module scoreboard_00000008_00000004
(
  clk_i,
  rst_ni,
  sb_full_o,
  flush_unissued_instr_i,
  flush_i,
  unresolved_branch_i,
  rd_clobber_gpr_o,
  rd_clobber_fpr_o,
  rs1_i,
  rs1_o,
  rs1_valid_o,
  rs2_i,
  rs2_o,
  rs2_valid_o,
  rs3_i,
  rs3_o,
  rs3_valid_o,
  commit_instr_o,
  commit_ack_i,
  decoded_instr_i,
  decoded_instr_valid_i,
  decoded_instr_ack_o,
  issue_instr_o,
  issue_instr_valid_o,
  issue_ack_i,
  resolved_branch_i,
  trans_id_i,
  wbdata_i,
  ex_i,
  wb_valid_i
);

  output [259:0] rd_clobber_gpr_o;
  output [259:0] rd_clobber_fpr_o;
  input [5:0] rs1_i;
  output [63:0] rs1_o;
  input [5:0] rs2_i;
  output [63:0] rs2_o;
  input [5:0] rs3_i;
  output [1:2] rs3_o;
  output [723:0] commit_instr_o;
  input [1:0] commit_ack_i;
  input [361:0] decoded_instr_i;
  output [361:0] issue_instr_o;
  input [133:0] resolved_branch_i;
  input [11:0] trans_id_i;
  input [255:0] wbdata_i;
  input [515:0] ex_i;
  input [3:0] wb_valid_i;
  input clk_i;
  input rst_ni;
  input flush_unissued_instr_i;
  input flush_i;
  input unresolved_branch_i;
  input decoded_instr_valid_i;
  input issue_ack_i;
  output sb_full_o;
  output rs1_valid_o;
  output rs2_valid_o;
  output rs3_valid_o;
  output decoded_instr_ack_o;
  output issue_instr_valid_o;
  wire [259:0] rd_clobber_gpr_o,rd_clobber_fpr_o;
  wire [63:0] rs1_o,rs2_o;
  wire [1:2] rs3_o;
  wire [723:0] commit_instr_o;
  wire sb_full_o,rs1_valid_o,rs2_valid_o,rs3_valid_o,decoded_instr_ack_o,
  issue_instr_valid_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,
  N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,
  N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,
  N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,
  N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,
  N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,
  N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,
  N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,
  N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,
  N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,
  N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,
  N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,
  N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,
  N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,
  N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,
  N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,
  N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,
  N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,
  N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,
  N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,
  N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,
  N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,
  N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,
  N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,
  N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,
  N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,
  N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,
  N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,
  N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,
  N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,
  N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,
  N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,
  N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,
  N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,
  N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,
  N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,
  N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,
  N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,
  N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,
  N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,
  N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,
  N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,
  N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,
  N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,
  N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,
  N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,
  N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,
  N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,
  N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,
  N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,
  N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
  N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,
  N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,
  N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,
  N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,
  N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,
  N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,
  N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,
  N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,
  N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,
  N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,
  N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,
  N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,
  N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,
  N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,
  N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,
  N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,
  N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,
  N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,
  N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,
  N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,
  N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,
  N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,
  N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,
  N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,
  N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,
  N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,
  N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,
  N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,
  N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,
  N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,
  N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,
  N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,
  N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,
  N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,
  N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,
  N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,
  N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,
  N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,
  N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,
  N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,
  N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,
  N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,
  N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,
  N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,
  N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,
  N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,
  N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,
  N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,
  N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,
  N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,
  N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,
  N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,
  N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,
  N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,
  N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,
  N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,
  N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,
  N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,
  N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,
  N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,
  N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,
  N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,
  N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,
  N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,
  N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,
  N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,
  N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,
  N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,
  N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,
  N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,
  N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,
  N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,
  N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,
  N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,
  N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,
  N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,
  N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,
  N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,
  N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,
  N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,
  N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,
  N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,
  N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,
  N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,
  N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,
  N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,
  N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,
  N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,
  N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,
  N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,
  N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,
  N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,
  N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,
  N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,
  N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,
  N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,
  N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,
  N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,
  N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,
  N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,
  N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,
  N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,
  N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,
  N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,
  N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,
  N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,
  N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,
  N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,
  N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,
  N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,
  N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,
  N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,
  N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,
  N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,
  N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,
  N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,
  N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,
  N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,
  N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,
  N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,
  N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,
  N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,
  N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,
  N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,
  N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,
  N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,
  N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,
  N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,
  N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,
  N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,
  N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,
  N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,
  N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,
  N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,
  N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,
  N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,
  N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,
  N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,
  N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,
  N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,
  N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,
  N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,
  N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,
  N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,
  N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,
  N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,
  N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,
  N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,
  N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,
  N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,
  N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,
  N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,
  N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,
  N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,
  N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,
  N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,
  N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,
  N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,
  N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,
  N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,
  N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,
  N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,
  N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,
  N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,
  N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,
  N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,
  N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,
  N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,
  N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,
  N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,
  N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,
  N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,N4143,
  N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,
  N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,
  N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,N4183,
  N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,
  N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,
  N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,N4223,
  N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,
  N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,
  N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,N4263,
  N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,
  N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,
  N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,N4303,
  N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,
  N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,
  N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,N4343,
  N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,
  N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,
  N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,N4383,
  N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,
  N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,
  N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,N4423,
  N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,
  N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,
  N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,N4463,
  N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,
  N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,
  N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,
  N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,
  N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,
  N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,
  N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,
  N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,
  N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,N4583,
  N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,
  N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,
  N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,
  N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,
  N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,
  N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,N4663,
  N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,
  N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,
  N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4703,
  N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,
  N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,
  N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,N4743,
  N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,
  N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,
  N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,
  N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,
  N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809,
  N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,N4821,N4822,N4823,
  N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,
  N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,N4849,
  N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,N4861,N4862,N4863,
  N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,
  N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,N4889,
  N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4903,
  N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,
  N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929,
  N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,N4941,N4942,N4943,
  N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,
  N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,N4969,
  N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,
  N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,
  N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,N5009,
  N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,N5021,N5022,N5023,
  N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,
  N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,N5049,
  N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,
  N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,
  N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,
  N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,
  N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,
  N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,
  N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,
  N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,
  N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,N5169,
  N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,
  N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,
  N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,
  N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,N5221,N5222,N5223,
  N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,
  N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,
  N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,N5263,
  N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,
  N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,N5289,
  N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5301,N5302,N5303,
  N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,
  N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,N5329,
  N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,N5341,N5342,N5343,
  N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,
  N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,N5369,
  N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,N5381,N5382,N5383,
  N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,
  N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,N5409,
  N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,N5421,N5422,N5423,
  N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,
  N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,N5449,
  N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,N5461,N5462,N5463,
  N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,
  N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,N5489,
  N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,N5501,N5502,N5503,
  N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,
  N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,N5529,
  N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,N5541,N5542,N5543,
  N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,
  N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,N5569,
  N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,N5581,N5582,N5583,
  N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,
  N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,N5609,
  N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5623,
  N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,
  N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,N5649,
  N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,N5661,N5662,N5663,
  N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,
  N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,N5689,
  N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,N5701,N5702,N5703,
  N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,
  N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,N5729,
  N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742,N5743,
  N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,
  N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,N5769,
  N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,N5781,N5782,N5783,
  N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,
  N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,N5809,
  N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,N5821,N5822,N5823,
  N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,
  N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,N5849,
  N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,N5861,N5862,N5863,
  N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,
  N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,N5889,
  N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,N5900,N5901,N5902,N5903,
  N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,
  N5917,N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,N5929,
  N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,N5940,N5941,N5942,N5943,
  N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,
  N5957,N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,N5969,
  N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5982,N5983,
  N5984,N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,
  N5997,N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,N6009,
  N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,N6019,N6020,N6021,N6022,N6023,
  N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,
  N6037,N6038,N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,N6048,N6049,
  N6050,N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060,N6061,N6062,N6063,
  N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,
  N6077,N6078,N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,N6088,N6089,
  N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,
  N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,
  N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,
  N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6141,N6142,N6143,
  N6144,N6145,N6146,N6147,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,
  N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,N6168,N6169,
  N6170,N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,N6179,N6180,N6181,N6182,N6183,
  N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,
  N6197,N6198,N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,N6208,N6209,
  N6210,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,N6219,N6220,N6221,N6222,N6223,
  N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6233,N6234,N6235,N6236,
  N6237,N6238,N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248,N6249,
  N6250,N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,N6263,
  N6264,N6265,N6266,N6267,N6268,N6269,N6270,N6271,N6272,N6273,N6274,N6275,N6276,
  N6277,N6278,N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,N6288,N6289,
  N6290,N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,N6299,N6300,N6301,N6302,N6303,
  N6304,N6305,N6306,N6307,N6308,N6309,N6310,N6311,N6312,N6313,N6314,N6315,N6316,
  N6317,N6318,N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,N6328,N6329,
  N6330,N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,N6339,N6340,N6341,N6342,N6343,
  N6344,N6345,N6346,N6347,N6348,N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356,
  N6357,N6358,N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,N6368,N6369,
  N6370,N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,N6379,N6380,N6381,N6382,N6383,
  N6384,N6385,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6393,N6394,N6395,N6396,
  N6397,N6398,N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,N6408,N6409,
  N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422,N6423,
  N6424,N6425,N6426,N6427,N6428,N6429,N6430,N6431,N6432,N6433,N6434,N6435,N6436,
  N6437,N6438,N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,N6448,N6449,
  N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,N6459,N6460,N6461,N6462,N6463,
  N6464,N6465,N6466,N6467,N6468,N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,
  N6477,N6478,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,N6488,N6489,
  N6490,N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,N6499,N6500,N6501,N6502,N6503,
  N6504,N6505,N6506,N6507,N6508,N6509,N6510,N6511,N6512,N6513,N6514,N6515,N6516,
  N6517,N6518,N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,N6528,N6529,
  N6530,N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,N6539,N6540,N6541,N6542,N6543,
  N6544,N6545,N6546,N6547,N6548,N6549,N6550,N6551,N6552,N6553,N6554,N6555,N6556,
  N6557,N6558,N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568,N6569,
  N6570,N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,N6579,N6580,N6581,N6582,N6583,
  N6584,N6585,N6586,N6587,N6588,N6589,N6590,N6591,N6592,N6593,N6594,N6595,N6596,
  N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,N6608,N6609,
  N6610,N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,N6619,N6620,N6621,N6622,N6623,
  N6624,N6625,N6626,N6627,N6628,N6629,N6630,N6631,N6632,N6633,N6634,N6635,N6636,
  N6637,N6638,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,
  N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6662,N6663,
  N6664,N6665,N6666,N6667,N6668,N6669,N6670,N6671,N6672,N6673,N6674,N6675,N6676,
  N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,
  N6690,N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,N6699,N6700,N6701,N6702,N6703,
  N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6716,
  N6717,N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,N6728,N6729,
  N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,N6739,N6740,N6741,N6742,N6743,
  N6744,N6745,N6746,N6747,N6748,N6749,N6750,N6751,N6752,N6753,N6754,N6755,N6756,
  N6757,N6758,N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,N6768,N6769,
  N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,N6783,
  N6784,N6785,N6786,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,
  N6797,N6798,N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,
  N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,N6819,N6820,N6821,N6822,N6823,
  N6824,N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6832,N6833,N6834,N6835,N6836,
  N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,N6848,N6849,
  N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,N6863,
  N6864,N6865,N6866,N6867,N6868,N6869,N6870,N6871,N6872,N6873,N6874,N6875,N6876,
  N6877,N6878,N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,N6888,N6889,
  N6890,N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,N6899,N6900,N6901,N6902,N6903,
  N6904,N6905,N6906,N6907,N6908,N6909,N6910,N6911,N6912,N6913,N6914,N6915,N6916,
  N6917,N6918,N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,N6928,N6929,
  N6930,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,N6939,N6940,N6941,N6942,N6943,
  N6944,N6945,N6946,N6947,N6948,N6949,N6950,N6951,N6952,N6953,N6954,N6955,N6956,
  N6957,N6958,N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,N6968,N6969,
  N6970,N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,N6979,N6980,N6981,N6982,N6983,
  N6984,N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992,N6993,N6994,N6995,N6996,
  N6997,N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,N7008,N7009,
  N7010,N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,N7019,N7020,N7021,N7022,N7023,
  N7024,N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032,N7033,N7034,N7035,N7036,
  N7037,N7038,N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,N7048,N7049,
  N7050,N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,N7059,N7060,N7061,N7062,N7063,
  N7064,N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072,N7073,N7074,N7075,N7076,
  N7077,N7078,N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088,N7089,
  N7090,N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,N7099,N7100,N7101,N7102,N7103,
  N7104,N7105,N7106,N7107,N7108,N7109,N7110,N7111,N7112,N7113,N7114,N7115,N7116,
  N7117,N7118,N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,N7128,N7129,
  N7130,N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,N7139,N7140,N7141,N7142,N7143,
  N7144,N7145,N7146,N7147,N7148,N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156,
  N7157,N7158,N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,N7168,N7169,
  N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,N7180,N7181,N7182,N7183,
  N7184,N7185,N7186,N7187,N7188,N7189,N7190,N7191,N7192,N7193,N7194,N7195,N7196,
  N7197,N7198,N7199,N7200,N7201,N7202,N7203,N7204,N7205,N7206,N7207,N7208,N7209,
  N7210,N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,N7219,N7220,N7221,N7222,N7223,
  N7224,N7225,N7226,N7227,N7228,N7229,N7230,N7231,N7232,N7233,N7234,N7235,N7236,
  N7237,N7238,N7239,N7240,N7241,N7242,N7243,N7244,N7245,N7246,N7247,N7248,N7249,
  N7250,N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,N7259,N7260,N7261,N7262,N7263,
  N7264,N7265,N7266,N7267,N7268,N7269,N7270,N7271,N7272,N7273,N7274,N7275,N7276,
  N7277,N7278,N7279,N7280,N7281,N7282,N7283,N7284,N7285,N7286,N7287,N7288,N7289,
  N7290,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,N7299,N7300,N7301,N7302,N7303,
  N7304,N7305,N7306,N7307,N7308,N7309,N7310,N7311,N7312,N7313,N7314,N7315,N7316,
  N7317,N7318,N7319,N7320,N7321,N7322,N7323,N7324,N7325,N7326,N7327,N7328,N7329,
  N7330,N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,N7339,N7340,N7341,N7342,N7343,
  N7344,N7345,N7346,N7347,N7348,N7349,N7350,N7351,N7352,N7353,N7354,N7355,N7356,
  N7357,N7358,N7359,N7360,N7361,N7362,N7363,N7364,N7365,N7366,N7367,N7368,N7369,
  N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,N7379,N7380,N7381,N7382,N7383,
  N7384,N7385,N7386,N7387,N7388,N7389,N7390,N7391,N7392,N7393,N7394,N7395,N7396,
  N7397,N7398,N7399,N7400,N7401,N7402,N7403,N7404,N7405,N7406,N7407,N7408,N7409,
  N7410,N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,N7419,N7420,N7421,N7422,N7423,
  N7424,N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7432,N7433,N7434,N7435,N7436,
  N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,N7449,
  N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,N7460,N7461,N7462,N7463,
  N7464,N7465,N7466,N7467,N7468,N7469,N7470,N7471,N7472,N7473,N7474,N7475,N7476,
  N7477,N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,N7487,N7488,N7489,
  N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,N7499,N7500,N7501,N7502,N7503,
  N7504,N7505,N7506,N7507,N7508,N7509,N7510,N7511,N7512,N7513,N7514,N7515,N7516,
  N7517,N7518,N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527,N7528,N7529,
  N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,N7539,N7540,N7541,N7542,N7543,
  N7544,N7545,N7546,N7547,N7548,N7549,N7550,N7551,N7552,N7553,N7554,N7555,N7556,
  N7557,N7558,N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567,N7568,N7569,
  N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,N7579,N7580,N7581,N7582,N7583,
  N7584,N7585,N7586,N7587,N7588,N7589,N7590,N7591,N7592,N7593,N7594,N7595,N7596,
  N7597,N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7608,N7609,
  N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,N7619,N7620,N7621,N7622,N7623,
  N7624,N7625,N7626,N7627,N7628,N7629,N7630,N7631,N7632,N7633,N7634,N7635,N7636,
  N7637,N7638,N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,N7647,N7648,N7649,
  N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,N7659,N7660,N7661,N7662,N7663,
  N7664,N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,
  N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,N7689,
  N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,N7699,N7700,N7701,N7702,N7703,
  N7704,N7705,N7706,N7707,N7708,N7709,N7710,N7711,N7712,N7713,N7714,N7715,N7716,
  N7717,N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,N7727,N7728,N7729,
  N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7743,
  N7744,N7745,N7746,N7747,N7748,N7749,N7750,N7751,N7752,N7753,N7754,N7755,N7756,
  N7757,N7758,N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,N7767,N7768,N7769,
  N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,N7779,N7780,N7781,N7782,N7783,
  N7784,N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792,N7793,N7794,N7795,N7796,
  N7797,N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,N7807,N7808,N7809,
  N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,N7819,N7820,N7821,N7822,N7823,
  N7824,N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832,N7833,N7834,N7835,N7836,
  N7837,N7838,N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,N7847,N7848,N7849,
  N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,N7859,N7860,N7861,N7862,N7863,
  N7864,N7865,N7866,N7867,N7868,N7869,N7870,N7871,N7872,N7873,N7874,N7875,N7876,
  N7877,N7878,N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,N7887,N7888,N7889,
  N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,N7899,N7900,N7901,N7902,N7903,
  N7904,N7905,N7906,N7907,N7908,N7909,N7910,N7911,N7912,N7913,N7914,N7915,N7916,
  N7917,N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,N7927,N7928,N7929,
  N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,N7939,N7940,N7941,N7942,N7943,
  N7944,N7945,N7946,N7947,N7948,N7949,N7950,N7951,N7952,N7953,N7954,N7955,N7956,
  N7957,N7958,N7959,N7960,N7961,N7962,N7963,N7964,N7965,N7966,N7967,N7968,N7969,
  N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,N7979,N7980,N7981,N7982,N7983,
  N7984,N7985,N7986,N7987,N7988,N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,
  N7997,N7998,N7999,N8000,N8001,N8002,N8003,N8004,N8005,N8006,N8007,N8008,N8009,
  N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,N8019,N8020,N8021,N8022,N8023,
  N8024,N8025,N8026,N8027,N8028,N8029,N8030,N8031,N8032,N8033,N8034,N8035,N8036,
  N8037,N8038,N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046,N8047,N8048,N8049,
  N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,N8059,N8060,N8061,N8062,N8063,
  N8064,N8065,N8066,N8067,N8068,N8069,N8070,N8071,N8072,N8073,N8074,N8075,N8076,
  N8077,N8078,N8079,N8080,N8081,N8082,N8083,N8084,N8085,N8086,N8087,N8088,N8089,
  N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,N8099,N8100,N8101,N8102,N8103,
  N8104,N8105,N8106,N8107,N8108,N8109,N8110,N8111,N8112,N8113,N8114,N8115,N8116,
  N8117,N8118,N8119,N8120,N8121,N8122,N8123,N8124,N8125,N8126,N8127,N8128,N8129,
  N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,N8139,N8140,N8141,N8142,N8143,
  N8144,N8145,N8146,N8147,N8148,N8149,N8150,N8151,N8152,N8153,N8154,N8155,N8156,
  N8157,N8158,N8159,N8160,N8161,N8162,N8163,N8164,N8165,N8166,N8167,N8168,N8169,
  N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,N8179,N8180,N8181,N8182,N8183,
  N8184,N8185,N8186,N8187,N8188,N8189,N8190,N8191,N8192,N8193,N8194,N8195,N8196,
  N8197,N8198,N8199,N8200,N8201,N8202,N8203,N8204,N8205,N8206,N8207,N8208,N8209,
  N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,N8219,N8220,N8221,N8222,N8223,
  N8224,N8225,N8226,N8227,N8228,N8229,N8230,N8231,N8232,N8233,N8234,N8235,N8236,
  N8237,N8238,N8239,N8240,N8241,N8242,N8243,N8244,N8245,N8246,N8247,N8248,N8249,
  N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,N8259,N8260,N8261,N8262,N8263,
  N8264,N8265,N8266,N8267,N8268,N8269,N8270,N8271,N8272,N8273,N8274,N8275,N8276,
  N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8286,N8287,N8288,N8289,
  N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,N8299,N8300,N8301,N8302,N8303,
  N8304,N8305,N8306,N8307,N8308,N8309,N8310,N8311,N8312,N8313,N8314,N8315,N8316,
  N8317,N8318,N8319,N8320,N8321,N8322,N8323,N8324,N8325,N8326,N8327,N8328,N8329,
  N8330,N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,N8339,N8340,N8341,N8342,N8343,
  N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,
  N8357,N8358,N8359,N8360,N8361,N8362,N8363,N8364,N8365,N8366,N8367,N8368,N8369,
  N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,
  N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,N8394,N8395,N8396,
  N8397,N8398,N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8406,N8407,N8408,N8409,
  N8410,N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,N8419,N8420,N8421,N8422,N8423,
  N8424,N8425,N8426,N8427,N8428,N8429,N8430,N8431,N8432,N8433,N8434,N8435,N8436,
  N8437,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8445,N8446,N8447,N8448,N8449,
  N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,N8459,N8460,N8461,N8462,N8463,
  N8464,N8465,N8466,N8467,N8468,N8469,N8470,N8471,N8472,N8473,N8474,N8475,N8476,
  N8477,N8478,N8479,N8480,N8481,N8482,N8483,N8484,N8485,N8486,N8487,N8488,N8489,
  N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,N8499,N8500,N8501,N8502,N8503,
  N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,N8513,N8514,N8515,N8516,
  N8517,N8518,N8519,N8520,N8521,N8522,N8523,N8524,N8525,N8526,N8527,N8528,N8529,
  N8530,N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,N8539,N8540,N8541,N8542,N8543,
  N8544,N8545,N8546,N8547,N8548,N8549,N8550,N8551,N8552,N8553,N8554,N8555,N8556,
  N8557,N8558,N8559,N8560,N8561,N8562,N8563,N8564,N8565,N8566,N8567,N8568,N8569,
  N8570,N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,N8579,N8580,N8581,N8582,N8583,
  N8584,N8585,N8586,N8587,N8588,N8589,N8590,N8591,N8592,N8593,N8594,N8595,N8596,
  N8597,N8598,N8599,N8600,N8601,N8602,N8603,N8604,N8605,N8606,N8607,N8608,N8609,
  N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,N8619,N8620,N8621,N8622,N8623,
  N8624,N8625,N8626,N8627,N8628,N8629,N8630,N8631,N8632,N8633,N8634,N8635,N8636,
  N8637,N8638,N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8646,N8647,N8648,N8649,
  N8650,N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,N8659,N8660,N8661,N8662,N8663,
  N8664,N8665,N8666,N8667,N8668,N8669,N8670,N8671,N8672,N8673,N8674,N8675,N8676,
  N8677,N8678,N8679,N8680,N8681,N8682,N8683,N8684,N8685,N8686,N8687,N8688,N8689,
  N8690,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,N8699,N8700,N8701,N8702,N8703,
  N8704,N8705,N8706,N8707,N8708,N8709,N8710,N8711,N8712,N8713,N8714,N8715,N8716,
  N8717,N8718,N8719,N8720,N8721,N8722,N8723,N8724,N8725,N8726,N8727,N8728,N8729,
  N8730,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,N8739,N8740,N8741,N8742,N8743,
  N8744,N8745,N8746,N8747,N8748,N8749,N8750,N8751,N8752,N8753,N8754,N8755,N8756,
  N8757,N8758,N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766,N8767,N8768,N8769,
  N8770,N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,N8779,N8780,N8781,N8782,N8783,
  N8784,N8785,N8786,N8787,N8788,N8789,N8790,N8791,N8792,N8793,N8794,N8795,N8796,
  N8797,N8798,N8799,N8800,N8801,N8802,N8803,N8804,N8805,N8806,N8807,N8808,N8809,
  N8810,N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,N8819,N8820,N8821,N8822,N8823,
  N8824,N8825,N8826,N8827,N8828,N8829,N8830,N8831,N8832,N8833,N8834,N8835,N8836,
  N8837,N8838,N8839,N8840,N8841,N8842,N8843,N8844,N8845,N8846,N8847,N8848,N8849,
  N8850,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,N8859,N8860,N8861,N8862,N8863,
  N8864,N8865,N8866,N8867,N8868,N8869,N8870,N8871,N8872,N8873,N8874,N8875,N8876,
  N8877,N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8889,
  N8890,N8891,N8892,N8893,N8894,N8895,N8896,N8897,N8898,N8899,N8900,N8901,N8902,N8903,
  N8904,N8905,N8906,N8907,N8908,N8909,N8910,N8911,N8912,N8913,N8914,N8915,N8916,
  N8917,N8918,N8919,N8920,N8921,N8922,N8923,N8924,N8925,N8926,N8927,N8928,N8929,
  N8930,N8931,N8932,N8933,N8934,N8935,N8936,N8937,N8938,N8939,N8940,N8941,N8942,N8943,
  N8944,N8945,N8946,N8947,N8948,N8949,N8950,N8951,N8952,N8953,N8954,N8955,N8956,
  N8957,N8958,N8959,N8960,N8961,N8962,N8963,N8964,N8965,N8966,N8967,N8968,N8969,
  N8970,N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978,N8979,N8980,N8981,N8982,N8983,
  N8984,N8985,N8986,N8987,N8988,N8989,N8990,N8991,N8992,N8993,N8994,N8995,N8996,
  N8997,N8998,N8999,N9000,N9001,N9002,N9003,N9004,N9005,N9006,N9007,N9008,N9009,
  N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017,N9018,N9019,N9020,N9021,N9022,N9023,
  N9024,N9025,N9026,N9027,N9028,N9029,N9030,N9031,N9032,N9033,N9034,N9035,N9036,
  N9037,N9038,N9039,N9040,N9041,N9042,N9043,N9044,N9045,N9046,N9047,N9048,N9049,
  N9050,N9051,N9052,N9053,N9054,N9055,N9056,N9057,N9058,N9059,N9060,N9061,N9062,N9063,
  N9064,N9065,N9066,N9067,N9068,N9069,N9070,N9071,N9072,N9073,N9074,N9075,N9076,
  N9077,N9078,N9079,N9080,N9081,N9082,N9083,N9084,N9085,N9086,N9087,N9088,N9089,
  N9090,N9091,N9092,N9093,N9094,N9095,N9096,N9097,N9098,N9099,N9100,N9101,N9102,N9103,
  N9104,N9105,N9106,N9107,N9108,N9109,N9110,N9111,N9112,N9113,N9114,N9115,N9116,
  N9117,N9118,N9119,N9120,N9121,N9122,N9123,N9124,N9125,N9126,N9127,N9128,N9129,
  N9130,N9131,N9132,N9133,N9134,N9135,N9136,N9137,N9138,N9139,N9140,N9141,N9142,N9143,
  N9144,N9145,N9146,N9147,N9148,N9149,N9150,N9151,N9152,N9153,N9154,N9155,N9156,
  N9157,N9158,N9159,N9160,N9161,N9162,N9163,N9164,N9165,N9166,N9167,N9168,N9169,
  N9170,N9171,N9172,N9173,N9174,N9175,N9176,N9177,N9178,N9179,N9180,N9181,N9182,N9183,
  N9184,N9185,N9186,N9187,N9188,N9189,N9190,N9191,N9192,N9193,N9194,N9195,N9196,
  N9197,N9198,N9199,N9200,N9201,N9202,N9203,N9204,N9205,N9206,N9207,N9208,N9209,
  N9210,N9211,N9212,N9213,N9214,N9215,N9216,N9217,N9218,N9219,N9220,N9221,N9222,N9223,
  N9224,N9225,N9226,N9227,N9228,N9229,N9230,N9231,N9232,N9233,N9234,N9235,N9236,
  N9237,N9238,N9239,N9240,N9241,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,
  N9250,N9251,N9252,N9253,N9254,N9255,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9263,
  N9264,N9265,N9266,N9267,N9268,N9269,N9270,N9271,N9272,N9273,N9274,N9275,N9276,
  N9277,N9278,N9279,N9280,N9281,N9282,N9283,N9284,N9285,N9286,N9287,N9288,N9289,
  N9290,N9291,N9292,N9293,N9294,N9295,N9296,N9297,N9298,N9299,N9300,N9301,N9302,N9303,
  N9304,N9305,N9306,N9307,N9308,N9309,N9310,N9311,N9312,N9313,N9314,N9315,N9316,
  N9317,N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9325,N9326,N9327,N9328,N9329,
  N9330,N9331,N9332,N9333,N9334,N9335,N9336,N9337,N9338,N9339,N9340,N9341,N9342,N9343,
  N9344,N9345,N9346,N9347,N9348,N9349,N9350,N9351,N9352,N9353,N9354,N9355,N9356,
  N9357,N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,
  N9370,N9371,N9372,N9373,N9374,N9375,N9376,N9377,N9378,N9379,N9380,N9381,N9382,N9383,
  N9384,N9385,N9386,N9387,N9388,N9389,N9390,N9391,N9392,N9393,N9394,N9395,N9396,
  N9397,N9398,N9399,N9400,N9401,N9402,N9403,N9404,N9405,N9406,N9407,N9408,N9409,
  N9410,N9411,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,N9420,N9421,N9422,N9423,
  N9424,N9425,N9426,N9427,N9428,N9429,N9430,N9431,N9432,N9433,N9434,N9435,N9436,
  N9437,N9438,N9439,N9440,N9441,N9442,N9443,N9444,N9445,N9446,N9447,N9448,N9449,
  N9450,N9451,N9452,N9453,N9454,N9455,N9456,N9457,N9458,N9459,N9460,N9461,N9462,N9463,
  N9464,N9465,N9466,N9467,N9468,N9469,N9470,N9471,N9472,N9473,N9474,N9475,N9476,
  N9477,N9478,N9479,N9480,N9481,N9482,N9483,N9484,N9485,N9486,N9487,N9488,N9489,
  N9490,N9491,N9492,N9493,N9494,N9495,N9496,N9497,N9498,N9499,N9500,N9501,N9502,N9503,
  N9504,N9505,N9506,N9507,N9508,N9509,N9510,N9511,N9512,N9513,N9514,N9515,N9516,
  N9517,N9518,N9519,N9520,N9521,N9522,N9523,N9524,N9525,N9526,N9527,N9528,N9529,
  N9530,N9531,N9532,N9533,N9534,N9535,N9536,N9537,N9538,N9539,N9540,N9541,N9542,N9543,
  N9544,N9545,N9546,N9547,N9548,N9549,N9550,N9551,N9552,N9553,N9554,N9555,N9556,
  N9557,N9558,N9559,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,N9569,
  N9570,N9571,N9572,N9573,N9574,N9575,N9576,N9577,N9578,N9579,N9580,N9581,N9582,N9583,
  N9584,N9585,N9586,N9587,N9588,N9589,N9590,N9591,N9592,N9593,N9594,N9595,N9596,
  N9597,N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9606,N9607,N9608,N9609,
  N9610,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,N9619,N9620,N9621,N9622,N9623,
  N9624,N9625,N9626,N9627,N9628,N9629,N9630,N9631,N9632,N9633,N9634,N9635,N9636,
  N9637,N9638,N9639,N9640,N9641,N9642,N9643,N9644,N9645,N9646,N9647,N9648,N9649,
  N9650,N9651,N9652,N9653,N9654,N9655,N9656,N9657,N9658,N9659,N9660,N9661,N9662,N9663,
  N9664,N9665,N9666,N9667,N9668,N9669,N9670,N9671,N9672,N9673,N9674,N9675,N9676,
  N9677,N9678,N9679,N9680,N9681,N9682,N9683,N9684,N9685,N9686,N9687,N9688,N9689,
  N9690,N9691,N9692,N9693,N9694,N9695,N9696,N9697,N9698,N9699,N9700,N9701,N9702,N9703,
  N9704,N9705,N9706,N9707,N9708,N9709,N9710,N9711,N9712,N9713,N9714,N9715,N9716,
  N9717,N9718,N9719,N9720,N9721,N9722,N9723,N9724,N9725,N9726,N9727,N9728,N9729,
  N9730,N9731,N9732,N9733,N9734,N9735,N9736,N9737,N9738,N9739,N9740,N9741,N9742,N9743,
  N9744,N9745,N9746,N9747,N9748,N9749,N9750,N9751,N9752,N9753,N9754,N9755,N9756,
  N9757,N9758,N9759,N9760,N9761,N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769,
  N9770,N9771,N9772,N9773,N9774,N9775,N9776,N9777,N9778,N9779,N9780,N9781,N9782,N9783,
  N9784,N9785,N9786,N9787,N9788,N9789,N9790,N9791,N9792,N9793,N9794,N9795,N9796,
  N9797,N9798,N9799,N9800,N9801,N9802,N9803,N9804,N9805,N9806,N9807,N9808,N9809,
  N9810,N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818,N9819,N9820,N9821,N9822,N9823,
  N9824,N9825,N9826,N9827,N9828,N9829,N9830,N9831,N9832,N9833,N9834,N9835,N9836,
  N9837,N9838,N9839,N9840,N9841,N9842,N9843,N9844,N9845,N9846,N9847,N9848,N9849,
  N9850,N9851,N9852,N9853,N9854,N9855,N9856,N9857,N9858,N9859,N9860,N9861,N9862,N9863,
  N9864,N9865,N9866,N9867,N9868,N9869,N9870,N9871,N9872,N9873,N9874,N9875,N9876,
  N9877,N9878,N9879,N9880,N9881,N9882,N9883,N9884,N9885,N9886,N9887,N9888,N9889,
  N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,N9902,N9903,
  N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9912,N9913,N9914,N9915,N9916,
  N9917,N9918,N9919,N9920,N9921,N9922,N9923,N9924,N9925,N9926,N9927,N9928,N9929,
  N9930,N9931,N9932,N9933,N9934,N9935,N9936,N9937,N9938,N9939,N9940,N9941,N9942,N9943,
  N9944,N9945,N9946,N9947,N9948,N9949,N9950,N9951,N9952,N9953,N9954,N9955,N9956,
  N9957,N9958,N9959,N9960,N9961,N9962,N9963,N9964,N9965,N9966,N9967,N9968,N9969,
  N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,N9979,N9980,N9981,N9982,N9983,
  N9984,N9985,N9986,N9987,N9988,N9989,N9990,N9991,N9992,N9993,N9994,N9995,N9996,
  N9997,N9998,N9999,N10000,N10001,N10002,N10003,N10004,N10005,N10006,N10007,N10008,
  N10009,N10010,N10011,N10012,N10013,N10014,N10015,N10016,N10017,N10018,N10019,
  N10020,N10021,N10022,N10023,N10024,N10025,N10026,N10027,N10028,N10029,N10030,N10031,
  N10032,N10033,N10034,N10035,N10036,N10037,N10038,N10039,N10040,N10041,N10042,
  N10043,N10044,N10045,N10046,N10047,N10048,N10049,N10050,N10051,N10052,N10053,
  N10054,N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10063,N10064,N10065,
  N10066,N10067,N10068,N10069,N10070,N10071,N10072,N10073,N10074,N10075,N10076,
  N10077,N10078,N10079,N10080,N10081,N10082,N10083,N10084,N10085,N10086,N10087,N10088,
  N10089,N10090,N10091,N10092,N10093,N10094,N10095,N10096,N10097,N10098,N10099,
  N10100,N10101,N10102,N10103,N10104,N10105,N10106,N10107,N10108,N10109,N10110,N10111,
  N10112,N10113,N10114,N10115,N10116,N10117,N10118,N10119,N10120,N10121,N10122,
  N10123,N10124,N10125,N10126,N10127,N10128,N10129,N10130,N10131,N10132,N10133,
  N10134,N10135,N10136,N10137,N10138,N10139,N10140,N10141,N10142,N10143,N10144,N10145,
  N10146,N10147,N10148,N10149,N10150,N10151,N10152,N10153,N10154,N10155,N10156,
  N10157,N10158,N10159,N10160,N10161,N10162,N10163,N10164,N10165,N10166,N10167,N10168,
  N10169,N10170,N10171,N10172,N10173,N10174,N10175,N10176,N10177,N10178,N10179,
  N10180,N10181,N10182,N10183,N10184,N10185,N10186,N10187,N10188,N10189,N10190,N10191,
  N10192,N10193,N10194,N10195,N10196,N10197,N10198,N10199,N10200,N10201,N10202,
  N10203,N10204,N10205,N10206,N10207,N10208,N10209,N10210,N10211,N10212,N10213,
  N10214,N10215,N10216,N10217,N10218,N10219,N10220,N10221,N10222,N10223,N10224,N10225,
  N10226,N10227,N10228,N10229,N10230,N10231,N10232,N10233,N10234,N10235,N10236,
  N10237,N10238,N10239,N10240,N10241,N10242,N10243,N10244,N10245,N10246,N10247,N10248,
  N10249,N10250,N10251,N10252,N10253,N10254,N10255,N10256,N10257,N10258,N10259,
  N10260,N10261,N10262,N10263,N10264,N10265,N10266,N10267,N10268,N10269,N10270,N10271,
  N10272,N10273,N10274,N10275,N10276,N10277,N10278,N10279,N10280,N10281,N10282,
  N10283,N10284,N10285,N10286,N10287,N10288,N10289,N10290,N10291,N10292,N10293,
  N10294,N10295,N10296,N10297,N10298,N10299,N10300,N10301,N10302,N10303,N10304,N10305,
  N10306,N10307,N10308,N10309,N10310,N10311,N10312,N10313,N10314,N10315,N10316,
  N10317,N10318,N10319,N10320,N10321,N10322,N10323,N10324,N10325,N10326,N10327,N10328,
  N10329,N10330,N10331,N10332,N10333,N10334,N10335,N10336,N10337,N10338,N10339,
  N10340,N10341,N10342,N10343,N10344,N10345,N10346,N10347,N10348,N10349,N10350,N10351,
  N10352,N10353,N10354,N10355,N10356,N10357,N10358,N10359,N10360,N10361,N10362,
  N10363,N10364,N10365,N10366,N10367,N10368,N10369,N10370,N10371,N10372,N10373,
  N10374,N10375,N10376,N10377,N10378,N10379,N10380,N10381,N10382,N10383,N10384,N10385,
  N10386,N10387,N10388,N10389,N10390,N10391,N10392,N10393,N10394,N10395,N10396,
  N10397,N10398,N10399,N10400,N10401,N10402,N10403,N10404,N10405,N10406,N10407,N10408,
  N10409,N10410,N10411,N10412,N10413,N10414,N10415,N10416,N10417,N10418,N10419,
  N10420,N10421,N10422,N10423,N10424,N10425,N10426,N10427,N10428,N10429,N10430,N10431,
  N10432,N10433,N10434,N10435,N10436,N10437,N10438,N10439,N10440,N10441,N10442,
  N10443,N10444,N10445,N10446,N10447,N10448,N10449,N10450,N10451,N10452,N10453,
  N10454,N10455,N10456,N10457,N10458,N10459,N10460,N10461,N10462,N10463,N10464,N10465,
  N10466,N10467,N10468,N10469,N10470,N10471,N10472,N10473,N10474,N10475,N10476,
  N10477,N10478,N10479,N10480,N10481,N10482,N10483,N10484,N10485,N10486,N10487,N10488,
  N10489,N10490,N10491,N10492,N10493,N10494,N10495,N10496,N10497,N10498,N10499,
  N10500,N10501,N10502,N10503,N10504,N10505,N10506,N10507,N10508,N10509,N10510,N10511,
  N10512,N10513,N10514,N10515,N10516,N10517,N10518,N10519,N10520,N10521,N10522,
  N10523,N10524,N10525,N10526,N10527,N10528,N10529,N10530,N10531,N10532,N10533,
  N10534,N10535,N10536,N10537,N10538,N10539,N10540,N10541,N10542,N10543,N10544,N10545,
  N10546,N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,
  N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,N10568,
  N10569,N10570,N10571,N10572,N10573,N10574,N10575,N10576,N10577,N10578,N10579,
  N10580,N10581,N10582,N10583,N10584,N10585,N10586,N10587,N10588,N10589,N10590,N10591,
  N10592,N10593,N10594,N10595,N10596,N10597,N10598,N10599,N10600,N10601,N10602,
  N10603,N10604,N10605,N10606,N10607,N10608,N10609,N10610,N10611,N10612,N10613,
  N10614,N10615,N10616,N10617,N10618,N10619,N10620,N10621,N10622,N10623,N10624,N10625,
  N10626,N10627,N10628,N10629,N10630,N10631,N10632,N10633,N10634,N10635,N10636,
  N10637,N10638,N10639,N10640,N10641,N10642,N10643,N10644,N10645,N10646,N10647,N10648,
  N10649,N10650,N10651,N10652,N10653,N10654,N10655,N10656,N10657,N10658,N10659,
  N10660,N10661,N10662,N10663,N10664,N10665,N10666,N10667,N10668,N10669,N10670,N10671,
  N10672,N10673,N10674,N10675,N10676,N10677,N10678,N10679,N10680,N10681,N10682,
  N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,N10692,N10693,
  N10694,N10695,N10696,N10697,N10698,N10699,N10700,N10701,N10702,N10703,N10704,N10705,
  N10706,N10707,N10708,N10709,N10710,N10711,N10712,N10713,N10714,N10715,N10716,
  N10717,N10718,N10719,N10720,N10721,N10722,N10723,N10724,N10725,N10726,N10727,N10728,
  N10729,N10730,N10731,N10732,N10733,N10734,N10735,N10736,N10737,N10738,N10739,
  N10740,N10741,N10742,N10743,N10744,N10745,N10746,N10747,N10748,N10749,N10750,N10751,
  N10752,N10753,N10754,N10755,N10756,N10757,N10758,N10759,N10760,N10761,N10762,
  N10763,N10764,N10765,N10766,N10767,N10768,N10769,N10770,N10771,N10772,N10773,
  N10774,N10775,N10776,N10777,N10778,N10779,N10780,N10781,N10782,N10783,N10784,N10785,
  N10786,N10787,N10788,N10789,N10790,N10791,N10792,N10793,N10794,N10795,N10796,
  N10797,N10798,N10799,N10800,N10801,N10802,N10803,N10804,N10805,N10806,N10807,N10808,
  N10809,N10810,N10811,N10812,N10813,N10814,N10815,N10816,N10817,N10818,N10819,
  N10820,N10821,N10822,N10823,N10824,N10825,N10826,N10827,N10828,N10829,N10830,N10831,
  N10832,N10833,N10834,N10835,N10836,N10837,N10838,N10839,N10840,N10841,N10842,
  N10843,N10844,N10845,N10846,N10847,N10848,N10849,N10850,N10851,N10852,N10853,
  N10854,N10855,N10856,N10857,N10858,N10859,N10860,N10861,N10862,N10863,N10864,N10865,
  N10866,N10867,N10868,N10869,N10870,N10871,N10872,N10873,N10874,N10875,N10876,
  N10877,N10878,N10879,N10880,N10881,N10882,N10883,N10884,N10885,N10886,N10887,N10888,
  N10889,N10890,N10891,N10892,N10893,N10894,N10895,N10896,N10897,N10898,N10899,
  N10900,N10901,N10902,N10903,N10904,N10905,N10906,N10907,N10908,N10909,N10910,N10911,
  N10912,N10913,N10914,N10915,N10916,N10917,N10918,N10919,N10920,N10921,N10922,
  N10923,N10924,N10925,N10926,N10927,N10928,N10929,N10930,N10931,N10932,N10933,
  N10934,N10935,N10936,N10937,N10938,N10939,N10940,N10941,N10942,N10943,N10944,N10945,
  N10946,N10947,N10948,N10949,N10950,N10951,N10952,N10953,N10954,N10955,N10956,
  N10957,N10958,N10959,N10960,N10961,N10962,N10963,N10964,N10965,N10966,N10967,N10968,
  N10969,N10970,N10971,N10972,N10973,N10974,N10975,N10976,N10977,N10978,N10979,
  N10980,N10981,N10982,N10983,N10984,N10985,N10986,N10987,N10988,N10989,N10990,N10991,
  N10992,N10993,N10994,N10995,N10996,N10997,N10998,N10999,N11000,N11001,N11002,
  N11003,N11004,N11005,N11006,N11007,N11008,N11009,N11010,N11011,N11012,N11013,
  N11014,N11015,N11016,N11017,N11018,N11019,N11020,N11021,N11022,N11023,N11024,N11025,
  N11026,N11027,N11028,N11029,N11030,N11031,N11032,N11033,N11034,N11035,N11036,
  N11037,N11038,N11039,N11040,N11041,N11042,N11043,N11044,N11045,N11046,N11047,N11048,
  N11049,N11050,N11051,N11052,N11053,N11054,N11055,N11056,N11057,N11058,N11059,
  N11060,N11061,N11062,N11063,N11064,N11065,N11066,N11067,N11068,N11069,N11070,N11071,
  N11072,N11073,N11074,N11075,N11076,N11077,N11078,N11079,N11080,N11081,N11082,
  N11083,N11084,N11085,N11086,N11087,N11088,N11089,N11090,N11091,N11092,N11093,
  N11094,N11095,N11096,N11097,N11098,N11099,N11100,N11101,N11102,N11103,N11104,N11105,
  N11106,N11107,N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,
  N11117,N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11125,N11126,N11127,N11128,
  N11129,N11130,N11131,N11132,N11133,N11134,N11135,N11136,N11137,N11138,N11139,
  N11140,N11141,N11142,N11143,N11144,N11145,N11146,N11147,N11148,N11149,N11150,N11151,
  N11152,N11153,N11154,N11155,N11156,N11157,N11158,N11159,N11160,N11161,N11162,
  N11163,N11164,N11165,N11166,N11167,N11168,N11169,N11170,N11171,N11172,N11173,
  N11174,N11175,N11176,N11177,N11178,N11179,N11180,N11181,N11182,N11183,N11184,N11185,
  N11186,N11187,N11188,N11189,N11190,N11191,N11192,N11193,N11194,N11195,N11196,
  N11197,N11198,N11199,N11200,N11201,N11202,N11203,N11204,N11205,N11206,N11207,N11208,
  N11209,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,
  N11220,N11221,N11222,N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11230,N11231,
  N11232,N11233,N11234,N11235,N11236,N11237,N11238,N11239,N11240,N11241,N11242,
  N11243,N11244,N11245,N11246,N11247,N11248,N11249,N11250,N11251,N11252,N11253,
  N11254,N11255,N11256,N11257,N11258,N11259,N11260,N11261,N11262,N11263,N11264,N11265,
  N11266,N11267,N11268,N11269,N11270,N11271,N11272,N11273,N11274,N11275,N11276,
  N11277,N11278,N11279,N11280,N11281,N11282,N11283,N11284,N11285,N11286,N11287,N11288,
  N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,N11298,N11299,
  N11300,N11301,N11302,N11303,N11304,N11305,N11306,N11307,N11308,N11309,N11310,N11311,
  N11312,N11313,N11314,N11315,N11316,N11317,N11318,N11319,N11320,N11321,N11322,
  N11323,N11324,N11325,N11326,N11327,N11328,N11329,N11330,N11331,N11332,N11333,
  N11334,N11335,N11336,N11337,N11338,N11339,N11340,N11341,N11342,N11343,N11344,N11345,
  N11346,N11347,N11348,N11349,N11350,N11351,N11352,N11353,N11354,N11355,N11356,
  N11357,N11358,N11359,N11360,N11361,N11362,N11363,N11364,N11365,N11366,N11367,N11368,
  N11369,N11370,N11371,N11372,N11373,N11374,N11375,N11376,N11377,N11378,N11379,
  N11380,N11381,N11382,N11383,N11384,N11385,N11386,N11387,N11388,N11389,N11390,N11391,
  N11392,N11393,N11394,N11395,N11396,N11397,N11398,N11399,N11400,N11401,N11402,
  N11403,N11404,N11405,N11406,N11407,N11408,N11409,N11410,N11411,N11412,N11413,
  N11414,N11415,N11416,N11417,N11418,N11419,N11420,N11421,N11422,N11423,N11424,N11425,
  N11426,N11427,N11428,N11429,N11430,N11431,N11432,N11433,N11434,N11435,N11436,
  N11437,N11438,N11439,N11440,N11441,N11442,N11443,N11444,N11445,N11446,N11447,N11448,
  N11449,N11450,N11451,N11452,N11453,N11454,N11455,N11456,N11457,N11458,N11459,
  N11460,N11461,N11462,N11463,N11464,N11465,N11466,N11467,N11468,N11469,N11470,N11471,
  N11472,N11473,N11474,N11475,N11476,N11477,N11478,N11479,N11480,N11481,N11482,
  N11483,N11484,N11485,N11486,N11487,N11488,N11489,N11490,N11491,N11492,N11493,
  N11494,N11495,N11496,N11497,N11498,N11499,N11500,N11501,N11502,N11503,N11504,N11505,
  N11506,N11507,N11508,N11509,N11510,N11511,N11512,N11513,N11514,N11515,N11516,
  N11517,N11518,N11519,N11520,N11521,N11522,N11523,N11524,N11525,N11526,N11527,N11528,
  N11529,N11530,N11531,N11532,N11533,N11534,N11535,N11536,N11537,N11538,N11539,
  N11540,N11541,N11542,N11543,N11544,N11545,N11546,N11547,N11548,N11549,N11550,N11551,
  N11552,N11553,N11554,N11555,N11556,N11557,N11558,N11559,N11560,N11561,N11562,
  N11563,N11564,N11565,N11566,N11567,N11568,N11569,N11570,N11571,N11572,N11573,
  N11574,N11575,N11576,N11577,N11578,N11579,N11580,N11581,N11582,N11583,N11584,N11585,
  N11586,N11587,N11588,N11589,N11590,N11591,N11592,N11593,N11594,N11595,N11596,
  N11597,N11598,N11599,N11600,N11601,N11602,N11603,N11604,N11605,N11606,N11607,N11608,
  N11609,N11610,N11611,N11612,N11613,N11614,N11615,N11616,N11617,N11618,N11619,
  N11620,N11621,N11622,N11623,N11624,N11625,N11626,N11627,N11628,N11629,N11630,N11631,
  N11632,N11633,N11634,N11635,N11636,N11637,N11638,N11639,N11640,N11641,N11642,
  N11643,N11644,N11645,N11646,N11647,N11648,N11649,N11650,N11651,N11652,N11653,
  N11654,N11655,N11656,N11657,N11658,N11659,N11660,N11661,N11662,N11663,N11664,N11665,
  N11666,N11667,N11668,N11669,N11670,N11671,N11672,N11673,N11674,N11675,N11676,
  N11677,N11678,N11679,N11680,N11681,N11682,N11683,N11684,N11685,N11686,N11687,N11688,
  N11689,N11690,N11691,N11692,N11693,N11694,N11695,N11696,N11697,N11698,N11699,
  N11700,N11701,N11702,N11703,N11704,N11705,N11706,N11707,N11708,N11709,N11710,N11711,
  N11712,N11713,N11714,N11715,N11716,N11717,N11718,N11719,N11720,N11721,N11722,
  N11723,N11724,N11725,N11726,N11727,N11728,N11729,N11730,N11731,N11732,N11733,
  N11734,N11735,N11736,N11737,N11738,N11739,N11740,N11741,N11742,N11743,N11744,N11745,
  N11746,N11747,N11748,N11749,N11750,N11751,N11752,N11753,N11754,N11755,N11756,
  N11757,N11758,N11759,N11760,N11761,N11762,N11763,N11764,N11765,N11766,N11767,N11768,
  N11769,N11770,N11771,N11772,N11773,N11774,N11775,N11776,N11777,N11778,N11779,
  N11780,N11781,N11782,N11783,N11784,N11785,N11786,N11787,N11788,N11789,N11790,N11791,
  N11792,N11793,N11794,N11795,N11796,N11797,N11798,N11799,N11800,N11801,N11802,
  N11803,N11804,N11805,N11806,N11807,N11808,N11809,N11810,N11811,N11812,N11813,
  N11814,N11815,N11816,N11817,N11818,N11819,N11820,N11821,N11822,N11823,N11824,N11825,
  N11826,N11827,N11828,N11829,N11830,N11831,N11832,N11833,N11834,N11835,N11836,
  N11837,N11838,N11839,N11840,N11841,N11842,N11843,N11844,N11845,N11846,N11847,N11848,
  N11849,N11850,N11851,N11852,N11853,N11854,N11855,N11856,N11857,N11858,N11859,
  N11860,N11861,N11862,N11863,N11864,N11865,N11866,N11867,N11868,N11869,N11870,N11871,
  N11872,N11873,N11874,N11875,N11876,N11877,N11878,N11879,N11880,N11881,N11882,
  N11883,N11884,N11885,N11886,N11887,N11888,N11889,N11890,N11891,N11892,N11893,
  N11894,N11895,N11896,N11897,N11898,N11899,N11900,N11901,N11902,N11903,N11904,N11905,
  N11906,N11907,N11908,N11909,N11910,N11911,N11912,N11913,N11914,N11915,N11916,
  N11917,N11918,N11919,N11920,N11921,N11922,N11923,N11924,N11925,N11926,N11927,N11928,
  N11929,N11930,N11931,N11932,N11933,N11934,N11935,N11936,N11937,N11938,N11939,
  N11940,N11941,N11942,N11943,N11944,N11945,N11946,N11947,N11948,N11949,N11950,N11951,
  N11952,N11953,N11954,N11955,N11956,N11957,N11958,N11959,N11960,N11961,N11962,
  N11963,N11964,N11965,N11966,N11967,N11968,N11969,N11970,N11971,N11972,N11973,
  N11974,N11975,N11976,N11977,N11978,N11979,N11980,N11981,N11982,N11983,N11984,N11985,
  N11986,N11987,N11988,N11989,N11990,N11991,N11992,N11993,N11994,N11995,N11996,
  N11997,N11998,N11999,N12000,N12001,N12002,N12003,N12004,N12005,N12006,N12007,N12008,
  N12009,N12010,N12011,N12012,N12013,N12014,N12015,N12016,N12017,N12018,N12019,
  N12020,N12021,N12022,N12023,N12024,N12025,N12026,N12027,N12028,N12029,N12030,N12031,
  N12032,N12033,N12034,N12035,N12036,N12037,N12038,N12039,N12040,N12041,N12042,
  N12043,N12044,N12045,N12046,N12047,N12048,N12049,N12050,N12051,N12052,N12053,
  N12054,N12055,N12056,N12057,N12058,N12059,N12060,N12061,N12062,N12063,N12064,N12065,
  N12066,N12067,N12068,N12069,N12070,N12071,N12072,N12073,N12074,N12075,N12076,
  N12077,N12078,N12079,N12080,N12081,N12082,N12083,N12084,N12085,N12086,N12087,N12088,
  N12089,N12090,N12091,N12092,N12093,N12094,N12095,N12096,N12097,N12098,N12099,
  N12100,N12101,N12102,N12103,N12104,N12105,N12106,N12107,N12108,N12109,N12110,N12111,
  N12112,N12113,N12114,N12115,N12116,N12117,N12118,N12119,N12120,N12121,N12122,
  N12123,N12124,N12125,N12126,N12127,N12128,N12129,N12130,N12131,N12132,N12133,
  N12134,N12135,N12136,N12137,N12138,N12139,N12140,N12141,N12142,N12143,N12144,N12145,
  N12146,N12147,N12148,N12149,N12150,N12151,N12152,N12153,N12154,N12155,N12156,
  N12157,N12158,N12159,N12160,N12161,N12162,N12163,N12164,N12165,N12166,N12167,N12168,
  N12169,N12170,N12171,N12172,N12173,N12174,N12175,N12176,N12177,N12178,N12179,
  N12180,N12181,N12182,N12183,N12184,N12185,N12186,N12187,N12188,N12189,N12190,N12191,
  N12192,N12193,N12194,N12195,N12196,N12197,N12198,N12199,N12200,N12201,N12202,
  N12203,N12204,N12205,N12206,N12207,N12208,N12209,N12210,N12211,N12212,N12213,
  N12214,N12215,N12216,N12217,N12218,N12219,N12220,N12221,N12222,N12223,N12224,N12225,
  N12226,N12227,N12228,N12229,N12230,N12231,N12232,N12233,N12234,N12235,N12236,
  N12237,N12238,N12239,N12240,N12241,N12242,N12243,N12244,N12245,N12246,N12247,N12248,
  N12249,N12250,N12251,N12252,N12253,N12254,N12255,N12256,N12257,N12258,N12259,
  N12260,N12261,N12262,N12263,N12264,N12265,N12266,N12267,N12268,N12269,N12270,N12271,
  N12272,N12273,N12274,N12275,N12276,N12277,N12278,N12279,N12280,N12281,N12282,
  N12283,N12284,N12285,N12286,N12287,N12288,N12289,N12290,N12291,N12292,N12293,
  N12294,N12295,N12296,N12297,N12298,N12299,N12300,N12301,N12302,N12303,N12304,N12305,
  N12306,N12307,N12308,N12309,N12310,N12311,N12312,N12313,N12314,N12315,N12316,
  N12317,N12318,N12319,N12320,N12321,N12322,N12323,N12324,N12325,N12326,N12327,N12328,
  N12329,N12330,N12331,N12332,N12333,N12334,N12335,N12336,N12337,N12338,N12339,
  N12340,N12341,N12342,N12343,N12344,N12345,N12346,N12347,N12348,N12349,N12350,N12351,
  N12352,N12353,N12354,N12355,N12356,N12357,N12358,N12359,N12360,N12361,N12362,
  N12363,N12364,N12365,N12366,N12367,N12368,N12369,N12370,N12371,N12372,N12373,
  N12374,N12375,N12376,N12377,N12378,N12379,N12380,N12381,N12382,N12383,N12384,N12385,
  N12386,N12387,N12388,N12389,N12390,N12391,N12392,N12393,N12394,N12395,N12396,
  N12397,N12398,N12399,N12400,N12401,N12402,N12403,N12404,N12405,N12406,N12407,N12408,
  N12409,N12410,N12411,N12412,N12413,N12414,N12415,N12416,N12417,N12418,N12419,
  N12420,N12421,N12422,N12423,N12424,N12425,N12426,N12427,N12428,N12429,N12430,N12431,
  N12432,N12433,N12434,N12435,N12436,N12437,N12438,N12439,N12440,N12441,N12442,
  N12443,N12444,N12445,N12446,N12447,N12448,N12449,N12450,N12451,N12452,N12453,
  N12454,N12455,N12456,N12457,N12458,N12459,N12460,N12461,N12462,N12463,N12464,N12465,
  N12466,N12467,N12468,N12469,N12470,N12471,N12472,N12473,N12474,N12475,N12476,
  N12477,N12478,N12479,N12480,N12481,N12482,N12483,N12484,N12485,N12486,N12487,N12488,
  N12489,N12490,N12491,N12492,N12493,N12494,N12495,N12496,N12497,N12498,N12499,
  N12500,N12501,N12502,N12503,N12504,N12505,N12506,N12507,N12508,N12509,N12510,N12511,
  N12512,N12513,N12514,N12515,N12516,N12517,N12518,N12519,N12520,N12521,N12522,
  N12523,N12524,N12525,N12526,N12527,N12528,N12529,N12530,N12531,N12532,N12533,
  N12534,N12535,N12536,N12537,N12538,N12539,N12540,N12541,N12542,N12543,N12544,N12545,
  N12546,N12547,N12548,N12549,N12550,N12551,N12552,N12553,N12554,N12555,N12556,
  N12557,N12558,N12559,N12560,N12561,N12562,N12563,N12564,N12565,N12566,N12567,N12568,
  N12569,N12570,N12571,N12572,N12573,N12574,N12575,N12576,N12577,N12578,N12579,
  N12580,N12581,N12582,N12583,N12584,N12585,N12586,N12587,N12588,N12589,N12590,N12591,
  N12592,N12593,N12594,N12595,N12596,N12597,N12598,N12599,N12600,N12601,N12602,
  N12603,N12604,N12605,N12606,N12607,N12608,N12609,N12610,N12611,N12612,N12613,
  N12614,N12615,N12616,N12617,N12618,N12619,N12620,N12621,N12622,N12623,N12624,N12625,
  N12626,N12627,N12628,N12629,N12630,N12631,N12632,N12633,N12634,N12635,N12636,
  N12637,N12638,N12639,N12640,N12641,N12642,N12643,N12644,N12645,N12646,N12647,N12648,
  N12649,N12650,N12651,N12652,N12653,N12654,N12655,N12656,N12657,N12658,N12659,
  N12660,N12661,N12662,N12663,N12664,N12665,N12666,N12667,N12668,N12669,N12670,N12671,
  N12672,N12673,N12674,N12675,N12676,N12677,N12678,N12679,N12680,N12681,N12682,
  N12683,N12684,N12685,N12686,N12687,N12688,N12689,N12690,N12691,N12692,N12693,
  N12694,N12695,N12696,N12697,N12698,N12699,N12700,N12701,N12702,N12703,N12704,N12705,
  N12706,N12707,N12708,N12709,N12710,N12711,N12712,N12713,N12714,N12715,N12716,
  N12717,N12718,N12719,N12720,N12721,N12722,N12723,N12724,N12725,N12726,N12727,N12728,
  N12729,N12730,N12731,N12732,N12733,N12734,N12735,N12736,N12737,N12738,N12739,
  N12740,N12741,N12742,N12743,N12744,N12745,N12746,N12747,N12748,N12749,N12750,N12751,
  N12752,N12753,N12754,N12755,N12756,N12757,N12758,N12759,N12760,N12761,N12762,
  N12763,N12764,N12765,N12766,N12767,N12768,N12769,N12770,N12771,N12772,N12773,
  N12774,N12775,N12776,N12777,N12778,N12779,N12780,N12781,N12782,N12783,N12784,N12785,
  N12786,N12787,N12788,N12789,N12790,N12791,N12792,N12793,N12794,N12795,N12796,
  N12797,N12798,N12799,N12800,N12801,N12802,N12803,N12804,N12805,N12806,N12807,N12808,
  N12809,N12810,N12811,N12812,N12813,N12814,N12815,N12816,N12817,N12818,N12819,
  N12820,N12821,N12822,N12823,N12824,N12825,N12826,N12827,N12828,N12829,N12830,N12831,
  N12832,N12833,N12834,N12835,N12836,N12837,N12838,N12839,N12840,N12841,N12842,
  N12843,N12844,N12845,N12846,N12847,N12848,N12849,N12850,N12851,N12852,N12853,
  N12854,N12855,N12856,N12857,N12858,N12859,N12860,N12861,N12862,N12863,N12864,N12865,
  N12866,N12867,N12868,N12869,N12870,N12871,N12872,N12873,N12874,N12875,N12876,
  N12877,N12878,N12879,N12880,N12881,N12882,N12883,N12884,N12885,N12886,N12887,N12888,
  N12889,N12890,N12891,N12892,N12893,N12894,N12895,N12896,N12897,N12898,N12899,
  N12900,N12901,N12902,N12903,N12904,N12905,N12906,N12907,N12908,N12909,N12910,N12911,
  N12912,N12913,N12914,N12915,N12916,N12917,N12918,N12919,N12920,N12921,N12922,
  N12923,N12924,N12925,N12926,N12927,N12928,N12929,N12930,N12931,N12932,N12933,
  N12934,N12935,N12936,N12937,N12938,N12939,N12940,N12941,N12942,N12943,N12944,N12945,
  N12946,N12947,N12948,N12949,N12950,N12951,N12952,N12953,N12954,N12955,N12956,
  N12957,N12958,N12959,N12960,N12961,N12962,N12963,N12964,N12965,N12966,N12967,N12968,
  N12969,N12970,N12971,N12972,N12973,N12974,N12975,N12976,N12977,N12978,N12979,
  N12980,N12981,N12982,N12983,N12984,N12985,N12986,N12987,N12988,N12989,N12990,N12991,
  N12992,N12993,N12994,N12995,N12996,N12997,N12998,N12999,N13000,N13001,N13002,
  N13003,N13004,N13005,N13006,N13007,N13008,N13009,N13010,N13011,N13012,N13013,
  N13014,N13015,N13016,N13017,N13018,N13019,N13020,N13021,N13022,N13023,N13024,N13025,
  N13026,N13027,N13028,N13029,N13030,N13031,N13032,N13033,N13034,N13035,N13036,
  N13037,N13038,N13039,N13040,N13041,N13042,N13043,N13044,N13045,N13046,N13047,N13048,
  N13049,N13050,N13051,N13052,N13053,N13054,N13055,N13056,N13057,N13058,N13059,
  N13060,N13061,N13062,N13063,N13064,N13065,N13066,N13067,N13068,N13069,N13070,N13071,
  N13072,N13073,N13074,N13075,N13076,N13077,N13078,N13079,N13080,N13081,N13082,
  N13083,N13084,N13085,N13086,N13087,N13088,N13089,N13090,N13091,N13092,N13093,
  N13094,N13095,N13096,N13097,N13098,N13099,N13100,N13101,N13102,N13103,N13104,N13105,
  N13106,N13107,N13108,N13109,N13110,N13111,N13112,N13113,N13114,N13115,N13116,
  N13117,N13118,N13119,N13120,N13121,N13122,N13123,N13124,N13125,N13126,N13127,N13128,
  N13129,N13130,N13131,N13132,N13133,N13134,N13135,N13136,N13137,N13138,N13139,
  N13140,N13141,N13142,N13143,N13144,N13145,N13146,N13147,N13148,N13149,N13150,N13151,
  N13152,N13153,N13154,N13155,N13156,N13157,N13158,N13159,N13160,N13161,N13162,
  N13163,N13164,N13165,N13166,N13167,N13168,N13169,N13170,N13171,N13172,N13173,
  N13174,N13175,N13176,N13177,N13178,N13179,N13180,N13181,N13182,N13183,N13184,N13185,
  N13186,N13187,N13188,N13189,N13190,N13191,N13192,N13193,N13194,N13195,N13196,
  N13197,N13198,N13199,N13200,N13201,N13202,N13203,N13204,N13205,N13206,N13207,N13208,
  N13209,N13210,N13211,N13212,N13213,N13214,N13215,N13216,N13217,N13218,N13219,
  N13220,N13221,N13222,N13223,N13224,N13225,N13226,N13227,N13228,N13229,N13230,N13231,
  N13232,N13233,N13234,N13235,N13236,N13237,N13238,N13239,N13240,N13241,N13242,
  N13243,N13244,N13245,N13246,N13247,N13248,N13249,N13250,N13251,N13252,N13253,
  N13254,N13255,N13256,N13257,N13258,N13259,N13260,N13261,N13262,N13263,N13264,N13265,
  N13266,N13267,N13268,N13269,N13270,N13271,N13272,N13273,N13274,N13275,N13276,
  N13277,N13278,N13279,N13280,N13281,N13282,N13283,N13284,N13285,N13286,N13287,N13288,
  N13289,N13290,N13291,N13292,N13293,N13294,N13295,N13296,N13297,N13298,N13299,
  N13300,N13301,N13302,N13303,N13304,N13305,N13306,N13307,N13308,N13309,N13310,N13311,
  N13312,N13313,N13314,N13315,N13316,N13317,N13318,N13319,N13320,N13321,N13322,
  N13323,N13324,N13325,N13326,N13327,N13328,N13329,N13330,N13331,N13332,N13333,
  N13334,N13335,N13336,N13337,N13338,N13339,N13340,N13341,N13342,N13343,N13344,N13345,
  N13346,N13347,N13348,N13349,N13350,N13351,N13352,N13353,N13354,N13355,N13356,
  N13357,N13358,N13359,N13360,N13361,N13362,N13363,N13364,N13365,N13366,N13367,N13368,
  N13369,N13370,N13371,N13372,N13373,N13374,N13375,N13376,N13377,N13378,N13379,
  N13380,N13381,N13382,N13383,N13384,N13385,N13386,N13387,N13388,N13389,N13390,N13391,
  N13392,N13393,N13394,N13395,N13396,N13397,N13398,N13399,N13400,N13401,N13402,
  N13403,N13404,N13405,N13406,N13407,N13408,N13409,N13410,N13411,N13412,N13413,
  N13414,N13415,N13416,N13417,N13418,N13419,N13420,N13421,N13422,N13423,N13424,N13425,
  N13426,N13427,N13428,N13429,N13430,N13431,N13432,N13433,N13434,N13435,N13436,
  N13437,N13438,N13439,N13440,N13441,N13442,N13443,N13444,N13445,N13446,N13447,N13448,
  N13449,N13450,N13451,N13452,N13453,N13454,N13455,N13456,N13457,N13458,N13459,
  N13460,N13461,N13462,N13463,N13464,N13465,N13466,N13467,N13468,N13469,N13470,N13471,
  N13472,N13473,N13474,N13475,N13476,N13477,N13478,N13479,N13480,N13481,N13482,
  N13483,N13484,N13485,N13486,N13487,N13488,N13489,N13490,N13491,N13492,N13493,
  N13494,N13495,N13496,N13497,N13498,N13499,N13500,N13501,N13502,N13503,N13504,N13505,
  N13506,N13507,N13508,N13509,N13510,N13511,N13512,N13513,N13514,N13515,N13516,
  N13517,N13518,N13519,N13520,N13521,N13522,N13523,N13524,N13525,N13526,N13527,N13528,
  N13529,N13530,N13531,N13532,N13533,N13534,N13535,N13536,N13537,N13538,N13539,
  N13540,N13541,N13542,N13543,N13544,N13545,N13546,N13547,N13548,N13549,N13550,N13551,
  N13552,N13553,N13554,N13555,N13556,N13557,N13558,N13559,N13560,N13561,N13562,
  N13563,N13564,N13565,N13566,N13567,N13568,N13569,N13570,N13571,N13572,N13573,
  N13574,N13575,N13576,N13577,N13578,N13579,N13580,N13581,N13582,N13583,N13584,N13585,
  N13586,N13587,N13588,N13589,N13590,N13591,N13592,N13593,N13594,N13595,N13596,
  N13597,N13598,N13599,N13600,N13601,N13602,N13603,N13604,N13605,N13606,N13607,N13608,
  N13609,N13610,N13611,N13612,N13613,N13614,N13615,N13616,N13617,N13618,N13619,
  N13620,N13621,N13622,N13623,N13624,N13625,N13626,N13627,N13628,N13629,N13630,N13631,
  N13632,N13633,N13634,N13635,N13636,N13637,N13638,N13639,N13640,N13641,N13642,
  N13643,N13644,N13645,N13646,N13647,N13648,N13649,N13650,N13651,N13652,N13653,
  N13654,N13655,N13656,N13657,N13658,N13659,N13660,N13661,N13662,N13663,N13664,N13665,
  N13666,N13667,N13668,N13669,N13670,N13671,N13672,N13673,N13674,N13675,N13676,
  N13677,N13678,N13679,N13680,N13681,N13682,N13683,N13684,N13685,N13686,N13687,N13688,
  N13689,N13690,N13691,N13692,N13693,N13694,N13695,N13696,N13697,N13698,N13699,
  N13700,N13701,N13702,N13703,N13704,N13705,N13706,N13707,N13708,N13709,N13710,N13711,
  N13712,N13713,N13714,N13715,N13716,N13717,N13718,N13719,N13720,N13721,N13722,
  N13723,N13724,N13725,N13726,N13727,N13728,N13729,N13730,N13731,N13732,N13733,
  N13734,N13735,N13736,N13737,N13738,N13739,N13740,N13741,N13742,N13743,N13744,N13745,
  N13746,N13747,N13748,N13749,N13750,N13751,N13752,N13753,N13754,N13755,N13756,
  N13757,N13758,N13759,N13760,N13761,N13762,N13763,N13764,N13765,N13766,N13767,N13768,
  N13769,N13770,N13771,N13772,N13773,N13774,N13775,N13776,N13777,N13778,N13779,
  N13780,N13781,N13782,N13783,N13784,N13785,N13786,N13787,N13788,N13789,N13790,N13791,
  N13792,N13793,N13794,N13795,N13796,N13797,N13798,N13799,N13800,N13801,N13802,
  N13803,N13804,N13805,N13806,N13807,N13808,N13809,N13810,N13811,N13812,N13813,
  N13814,N13815,N13816,N13817,N13818,N13819,N13820,N13821,N13822,N13823,N13824,N13825,
  N13826,N13827,N13828,N13829,N13830,N13831,N13832,N13833,N13834,N13835,N13836,
  N13837,N13838,N13839,N13840,N13841,N13842,N13843,N13844,N13845,N13846,N13847,N13848,
  N13849,N13850,N13851,N13852,N13853,N13854,N13855,N13856,N13857,N13858,N13859,
  N13860,N13861,N13862,N13863,N13864,N13865,N13866,N13867,N13868,N13869,N13870,N13871,
  N13872,N13873,N13874,N13875,N13876,N13877,N13878,N13879,N13880,N13881,N13882,
  N13883,N13884,N13885,N13886,N13887,N13888,N13889,N13890,N13891,N13892,N13893,
  N13894,N13895,N13896,N13897,N13898,N13899,N13900,N13901,N13902,N13903,N13904,N13905,
  N13906,N13907,N13908,N13909,N13910,N13911,N13912,N13913,N13914,N13915,N13916,
  N13917,N13918,N13919,N13920,N13921,N13922,N13923,N13924,N13925,N13926,N13927,N13928,
  N13929,N13930,N13931,N13932,N13933,N13934,N13935,N13936,N13937,N13938,N13939,
  N13940,N13941,N13942,N13943,N13944,N13945,N13946,N13947,N13948,N13949,N13950,N13951,
  N13952,N13953,N13954,N13955,N13956,N13957,N13958,N13959,N13960,N13961,N13962,
  N13963,N13964,N13965,N13966,N13967,N13968,N13969,N13970,N13971,N13972,N13973,
  N13974,N13975,N13976,N13977,N13978,N13979,N13980,N13981,N13982,N13983,N13984,N13985,
  N13986,N13987,N13988,N13989,N13990,N13991,N13992,N13993,N13994,N13995,N13996,
  N13997,N13998,N13999,N14000,N14001,N14002,N14003,N14004,N14005,N14006,N14007,N14008,
  N14009,N14010,N14011,N14012,N14013,N14014,N14015,N14016,N14017,N14018,N14019,
  N14020,N14021,N14022,N14023,N14024,N14025,N14026,N14027,N14028,N14029,N14030,N14031,
  N14032,N14033,N14034,N14035,N14036,N14037,N14038,N14039,N14040,N14041,N14042,
  N14043,N14044,N14045,N14046,N14047,N14048,N14049,N14050,N14051,N14052,N14053,
  N14054,N14055,N14056,N14057,N14058,N14059,N14060,N14061,N14062,N14063,N14064,N14065,
  N14066,N14067,N14068,N14069,N14070,N14071,N14072,N14073,N14074,N14075,N14076,
  N14077,N14078,N14079,N14080,N14081,N14082,N14083,N14084,N14085,N14086,N14087,N14088,
  N14089,N14090,N14091,N14092,N14093,N14094,N14095,N14096,N14097,N14098,N14099,
  N14100,N14101,N14102,N14103,N14104,N14105,N14106,N14107,N14108,N14109,N14110,N14111,
  N14112,N14113,N14114,N14115,N14116,N14117,N14118,N14119,N14120,N14121,N14122,
  N14123,N14124,N14125,N14126,N14127,N14128,N14129,N14130,N14131,N14132,N14133,
  N14134,N14135,N14136,N14137,N14138,N14139,N14140,N14141,N14142,N14143,N14144,N14145,
  N14146,N14147,N14148,N14149,N14150,N14151,N14152,N14153,N14154,N14155,N14156,
  N14157,N14158,N14159,N14160,N14161,N14162,N14163,N14164,N14165,N14166,N14167,N14168,
  N14169,N14170,N14171,N14172,N14173,N14174,N14175,N14176,N14177,N14178,N14179,
  N14180,N14181,N14182,N14183,N14184,N14185,N14186,N14187,N14188,N14189,N14190,N14191,
  N14192,N14193,N14194,N14195,N14196,N14197,N14198,N14199,N14200,N14201,N14202,
  N14203,N14204,N14205,N14206,N14207,N14208,N14209,N14210,N14211,N14212,N14213,
  N14214,N14215,N14216,N14217,N14218,N14219,N14220,N14221,N14222,N14223,N14224,N14225,
  N14226,N14227,N14228,N14229,N14230,N14231,N14232,N14233,N14234,N14235,N14236,
  N14237,N14238,N14239,N14240,N14241,N14242,N14243,N14244,N14245,N14246,N14247,N14248,
  N14249,N14250,N14251,N14252,N14253,N14254,N14255,N14256,N14257,N14258,N14259,
  N14260,N14261,N14262,N14263,N14264,N14265,N14266,N14267,N14268,N14269,N14270,N14271,
  N14272,N14273,N14274,N14275,N14276,N14277,N14278,N14279,N14280,N14281,N14282,
  N14283,N14284,N14285,N14286,N14287,N14288,N14289,N14290,N14291,N14292,N14293,
  N14294,N14295,N14296,N14297,N14298,N14299,N14300,N14301,N14302,N14303,N14304,N14305,
  N14306,N14307,N14308,N14309,N14310,N14311,N14312,N14313,N14314,N14315,N14316,
  N14317,N14318,N14319,N14320,N14321,N14322,N14323,N14324,N14325,N14326,N14327,N14328,
  N14329,N14330,N14331,N14332,N14333,N14334,N14335,N14336,N14337,N14338,N14339,
  N14340,N14341,N14342,N14343,N14344,N14345,N14346,N14347,N14348,N14349,N14350,N14351,
  N14352,N14353,N14354,N14355,N14356,N14357,N14358,N14359,N14360,N14361,N14362,
  N14363,N14364,N14365,N14366,N14367,N14368,N14369,N14370,N14371,N14372,N14373,
  N14374,N14375,N14376,N14377,N14378,N14379,N14380,N14381,N14382,N14383,N14384,N14385,
  N14386,N14387,N14388,N14389,N14390,N14391,N14392,N14393,N14394,N14395,N14396,
  N14397,N14398,N14399,N14400,N14401,N14402,N14403,N14404,N14405,N14406,N14407,N14408,
  N14409,N14410,N14411,N14412,N14413,N14414,N14415,N14416,N14417,N14418,N14419,
  N14420,N14421,N14422,N14423,N14424,N14425,N14426,N14427,N14428,N14429,N14430,N14431,
  N14432,N14433,N14434,N14435,N14436,N14437,N14438,N14439,N14440,N14441,N14442,
  N14443,N14444,N14445,N14446,N14447,N14448,N14449,N14450,N14451,N14452,N14453,
  N14454,N14455,N14456,N14457,N14458,N14459,N14460,N14461,N14462,N14463,N14464,N14465,
  N14466,N14467,N14468,N14469,N14470,N14471,N14472,N14473,N14474,N14475,N14476,
  N14477,N14478,N14479,N14480,N14481,N14482,N14483,N14484,N14485,N14486,N14487,N14488,
  N14489,N14490,N14491,N14492,N14493,N14494,N14495,N14496,N14497,N14498,N14499,
  N14500,N14501,N14502,N14503,N14504,N14505,N14506,N14507,N14508,N14509,N14510,N14511,
  N14512,N14513,N14514,N14515,N14516,N14517,N14518,N14519,N14520,N14521,N14522,
  N14523,N14524,N14525,N14526,N14527,N14528,N14529,N14530,N14531,N14532,N14533,
  N14534,N14535,N14536,N14537,N14538,N14539,N14540,N14541,N14542,N14543,N14544,N14545,
  N14546,N14547,N14548,N14549,N14550,N14551,N14552,N14553,N14554,N14555,N14556,
  N14557,N14558,N14559,N14560,N14561,N14562,N14563,N14564,N14565,N14566,N14567,N14568,
  N14569,N14570,N14571,N14572,N14573,N14574,N14575,N14576,N14577,N14578,N14579,
  N14580,N14581,N14582,N14583,N14584,N14585,N14586,N14587,N14588,N14589,N14590,N14591,
  N14592,N14593,N14594,N14595,N14596,N14597,N14598,N14599,N14600,N14601,N14602,
  N14603,N14604,N14605,N14606,N14607,N14608,N14609,N14610,N14611,N14612,N14613,
  N14614,N14615,N14616,N14617,N14618,N14619,N14620,N14621,N14622,N14623,N14624,N14625,
  N14626,N14627,N14628,N14629,N14630,N14631,N14632,N14633,N14634,N14635,N14636,
  N14637,N14638,N14639,N14640,N14641,N14642,N14643,N14644,N14645,N14646,N14647,N14648,
  N14649,N14650,N14651,N14652,N14653,N14654,N14655,N14656,N14657,N14658,N14659,
  N14660,N14661,N14662,N14663,N14664,N14665,N14666,N14667,N14668,N14669,N14670,N14671,
  N14672,N14673,N14674,N14675,N14676,N14677,N14678,N14679,N14680,N14681,N14682,
  N14683,N14684,N14685,N14686,N14687,N14688,N14689,N14690,N14691,N14692,N14693,
  N14694,N14695,N14696,N14697,N14698,N14699,N14700,N14701,N14702,N14703,N14704,N14705,
  N14706,N14707,N14708,N14709,N14710,N14711,N14712,N14713,N14714,N14715,N14716,
  N14717,N14718,N14719,N14720,N14721,N14722,N14723,N14724,N14725,N14726,N14727,N14728,
  N14729,N14730,N14731,N14732,N14733,N14734,N14735,N14736,N14737,N14738,N14739,
  N14740,N14741,N14742,N14743,N14744,N14745,N14746,N14747,N14748,N14749,N14750,N14751,
  N14752,N14753,N14754,N14755,N14756,N14757,N14758,N14759,N14760,N14761,N14762,
  N14763,N14764,N14765,N14766,N14767,N14768,N14769,N14770,N14771,N14772,N14773,
  N14774,N14775,N14776,N14777,N14778,N14779,N14780,N14781,N14782,N14783,N14784,N14785,
  N14786,N14787,N14788,N14789,N14790,N14791,N14792,N14793,N14794,N14795,N14796,
  N14797,N14798,N14799,N14800,N14801,N14802,N14803,N14804,N14805,N14806,N14807,N14808,
  N14809,N14810,N14811,N14812,N14813,N14814,N14815,N14816,N14817,N14818,N14819,
  N14820,N14821,N14822,N14823,N14824,N14825,N14826,N14827,N14828,N14829,N14830,N14831,
  N14832,N14833,N14834,N14835,N14836,N14837,N14838,N14839,N14840,N14841,N14842,
  N14843,N14844,N14845,N14846,N14847,N14848,N14849,N14850,N14851,N14852,N14853,
  N14854,N14855,N14856,N14857,N14858,N14859,N14860,N14861,N14862,N14863,N14864,N14865,
  N14866,N14867,N14868,N14869,N14870,N14871,N14872,N14873,N14874,N14875,N14876,
  N14877,N14878,N14879,N14880,N14881,N14882,N14883,N14884,N14885,N14886,N14887,N14888,
  N14889,N14890,N14891,N14892,N14893,N14894,N14895,N14896,N14897,N14898,N14899,
  N14900,N14901,N14902,N14903,N14904,N14905,N14906,N14907,N14908,N14909,N14910,N14911,
  N14912,N14913,N14914,N14915,N14916,N14917,N14918,N14919,N14920,N14921,N14922,
  N14923,N14924,N14925,N14926,N14927,N14928,N14929,N14930,N14931,N14932,N14933,
  N14934,N14935,N14936,N14937,N14938,N14939,N14940,N14941,N14942,N14943,N14944,N14945,
  N14946,N14947,N14948,N14949,N14950,N14951,N14952,N14953,N14954,N14955,N14956,
  N14957,N14958,N14959,N14960,N14961,N14962,N14963,N14964,N14965,N14966,N14967,N14968,
  N14969,N14970,N14971,N14972,N14973,N14974,N14975,N14976,N14977,N14978,N14979,
  N14980,N14981,N14982,N14983,N14984,N14985,N14986,N14987,N14988,N14989,N14990,N14991,
  N14992,N14993,N14994,N14995,N14996,N14997,N14998,N14999,N15000,N15001,N15002,
  N15003,N15004,N15005,N15006,N15007,N15008,N15009,N15010,N15011,N15012,N15013,
  N15014,N15015,N15016,N15017,N15018,N15019,N15020,N15021,N15022,N15023,N15024,N15025,
  N15026,N15027,N15028,N15029,N15030,N15031,N15032,N15033,N15034,N15035,N15036,
  N15037,N15038,N15039,N15040,N15041,N15042,N15043,N15044,N15045,N15046,N15047,N15048,
  N15049,N15050,N15051,N15052,N15053,N15054,N15055,N15056,N15057,N15058,N15059,
  N15060,N15061,N15062,N15063,N15064,N15065,N15066,N15067,N15068,N15069,N15070,N15071,
  N15072,N15073,N15074,N15075,N15076,N15077,N15078,N15079,N15080,N15081,N15082,
  N15083,N15084,N15085,N15086,N15087,N15088,N15089,N15090,N15091,N15092,N15093,
  N15094,N15095,N15096,N15097,N15098,N15099,N15100,N15101,N15102,N15103,N15104,N15105,
  N15106,N15107,N15108,N15109,N15110,N15111,N15112,N15113,N15114,N15115,N15116,
  N15117,N15118,N15119,N15120,N15121,N15122,N15123,N15124,N15125,N15126,N15127,N15128,
  N15129,N15130,N15131,N15132,N15133,N15134,N15135,N15136,N15137,N15138,N15139,
  N15140,N15141,N15142,N15143,N15144,N15145,N15146,N15147,N15148,N15149,N15150,N15151,
  N15152,N15153,N15154,N15155,N15156,N15157,N15158,N15159,N15160,N15161,N15162,
  N15163,N15164,N15165,N15166,N15167,N15168,N15169,N15170,N15171,N15172,N15173,
  N15174,N15175,N15176,N15177,N15178,N15179,N15180,N15181,N15182,N15183,N15184,N15185,
  N15186,N15187,N15188,N15189,N15190,N15191,N15192,N15193,N15194,N15195,N15196,
  N15197,N15198,N15199,N15200,N15201,N15202,N15203,N15204,N15205,N15206,N15207,N15208,
  N15209,N15210,N15211,N15212,N15213,N15214,N15215,N15216,N15217,N15218,N15219,
  N15220,N15221,N15222,N15223,N15224,N15225,N15226,N15227,N15228,N15229,N15230,N15231,
  N15232,N15233,N15234,N15235,N15236,N15237,N15238,N15239,N15240,N15241,N15242,
  N15243,N15244,N15245,N15246,N15247,N15248,N15249,N15250,N15251,N15252,N15253,
  N15254,N15255,N15256,N15257,N15258,N15259,N15260,N15261,N15262,N15263,N15264,N15265,
  N15266,N15267,N15268,N15269,N15270,N15271,N15272,N15273,N15274,N15275,N15276,
  N15277,N15278,N15279,N15280,N15281,N15282,N15283,N15284,N15285,N15286,N15287,N15288,
  N15289,N15290,N15291,N15292,N15293,N15294,N15295,N15296,N15297,N15298,N15299,
  N15300,N15301,N15302,N15303,N15304,N15305,N15306,N15307,N15308,N15309,N15310,N15311,
  N15312,N15313,N15314,N15315,N15316,N15317,N15318,N15319,N15320,N15321,N15322,
  N15323,N15324,N15325,N15326,N15327,N15328,N15329,N15330,N15331,N15332,N15333,
  N15334,N15335,N15336,N15337,N15338,N15339,N15340,N15341,N15342,N15343,N15344,N15345,
  N15346,N15347,N15348,N15349,N15350,N15351,N15352,N15353,N15354,N15355,N15356,
  N15357,N15358,N15359,N15360,N15361,N15362,N15363,N15364,N15365,N15366,N15367,N15368,
  N15369,N15370,N15371,N15372,N15373,N15374,N15375,N15376,N15377,N15378,N15379,
  N15380,N15381,N15382,N15383,N15384,N15385,N15386,N15387,N15388,N15389,N15390,N15391,
  N15392,N15393,N15394,N15395,N15396,N15397,N15398,N15399,N15400,N15401,N15402,
  N15403,N15404,N15405,N15406,N15407,N15408,N15409,N15410,N15411,N15412,N15413,
  N15414,N15415,N15416,N15417,N15418,N15419,N15420,N15421,N15422,N15423,N15424,N15425,
  N15426,N15427,N15428,N15429,N15430,N15431,N15432,N15433,N15434,N15435,N15436,
  N15437,N15438,N15439,N15440,N15441,N15442,N15443,N15444,N15445,N15446,N15447,N15448,
  N15449,N15450,N15451,N15452,N15453,N15454,N15455,N15456,N15457,N15458,N15459,
  N15460,N15461,N15462,N15463,N15464,N15465,N15466,N15467,N15468,N15469,N15470,N15471,
  N15472,N15473,N15474,N15475,N15476,N15477,N15478,N15479,N15480,N15481,N15482,
  N15483,N15484,N15485,N15486,N15487,N15488,N15489,N15490,N15491,N15492,N15493,
  N15494,N15495,N15496,N15497,N15498,N15499,N15500,N15501,N15502,N15503,N15504,N15505,
  N15506,N15507,N15508,N15509,N15510,N15511,N15512,N15513,N15514,N15515,N15516,
  N15517,N15518,N15519,N15520,N15521,N15522,N15523,N15524,N15525,N15526,N15527,N15528,
  N15529,N15530,N15531,N15532,N15533,N15534,N15535,N15536,N15537,N15538,N15539,
  N15540,N15541,N15542,N15543,N15544,N15545,N15546,N15547,N15548,N15549,N15550,N15551,
  N15552,N15553,N15554,N15555,N15556,N15557,N15558,N15559,N15560,N15561,N15562,
  N15563,N15564,N15565,N15566,N15567,N15568,N15569,N15570,N15571,N15572,N15573,
  N15574,N15575,N15576,N15577,N15578,N15579,N15580,N15581,N15582,N15583,N15584,N15585,
  N15586,N15587,N15588,N15589,N15590,N15591,N15592,N15593,N15594,N15595,N15596,
  N15597,N15598,N15599,N15600,N15601,N15602,N15603,N15604,N15605,N15606,N15607,N15608,
  N15609,N15610,N15611,N15612,N15613,N15614,N15615,N15616,N15617,N15618,N15619,
  N15620,N15621,N15622,N15623,N15624,N15625,N15626,N15627,N15628,N15629,N15630,N15631,
  N15632,N15633,N15634,N15635,N15636,N15637,N15638,N15639,N15640,N15641,N15642,
  N15643,N15644,N15645,N15646,N15647,N15648,N15649,N15650,N15651,N15652,N15653,
  N15654,N15655,N15656,N15657,N15658,N15659,N15660,N15661,N15662,N15663,N15664,N15665,
  N15666,N15667,N15668,N15669,N15670,N15671,N15672,N15673,N15674,N15675,N15676,
  N15677,N15678,N15679,N15680,N15681,N15682,N15683,N15684,N15685,N15686,N15687,N15688,
  N15689,N15690,N15691,N15692,N15693,N15694,N15695,N15696,N15697,N15698,N15699,
  N15700,N15701,N15702,N15703,N15704,N15705,N15706,N15707,N15708,N15709,N15710,N15711,
  N15712,N15713,N15714,N15715,N15716,N15717,N15718,N15719,N15720,N15721,N15722,
  N15723,N15724,N15725,N15726,N15727,N15728,N15729,N15730,N15731,N15732,N15733,
  N15734,N15735,N15736,N15737,N15738,N15739,N15740,N15741,N15742,N15743,N15744,N15745,
  N15746,N15747,N15748,N15749,N15750,N15751,N15752,N15753,N15754,N15755,N15756,
  N15757,N15758,N15759,N15760,N15761,N15762,N15763,N15764,N15765,N15766,N15767,N15768,
  N15769,N15770,N15771,N15772,N15773,N15774,N15775,N15776,N15777,N15778,N15779,
  N15780,N15781,N15782,N15783,N15784,N15785,N15786,N15787,N15788,N15789,N15790,N15791,
  N15792,N15793,N15794,N15795,N15796,N15797,N15798,N15799,N15800,N15801,N15802,
  N15803,N15804,N15805,N15806,N15807,N15808,N15809,N15810,N15811,N15812,N15813,
  N15814,N15815,N15816,N15817,N15818,N15819,N15820,N15821,N15822,N15823,N15824,N15825,
  N15826,N15827,N15828,N15829,N15830,N15831,N15832,N15833,N15834,N15835,N15836,
  N15837,N15838,N15839,N15840,N15841,N15842,N15843,N15844,N15845,N15846,N15847,N15848,
  N15849,N15850,N15851,N15852,N15853,N15854,N15855,N15856,N15857,N15858,N15859,
  N15860,N15861,N15862,N15863,N15864,N15865,N15866,N15867,N15868,N15869,N15870,N15871,
  N15872,N15873,N15874,N15875,N15876,N15877,N15878,N15879,N15880,N15881,N15882,
  N15883,N15884,N15885,N15886,N15887,N15888,N15889,N15890,N15891,N15892,N15893,
  N15894,N15895,N15896,N15897,N15898,N15899,N15900,N15901,N15902,N15903,N15904,N15905,
  N15906,N15907,N15908,N15909,N15910,N15911,N15912,N15913,N15914,N15915,N15916,
  N15917,N15918,N15919,N15920,N15921,N15922,N15923,N15924,N15925,N15926,N15927,N15928,
  N15929,N15930,N15931,N15932,N15933,N15934,N15935,N15936,N15937,N15938,N15939,
  N15940,N15941,N15942,N15943,N15944,N15945,N15946,N15947,N15948,N15949,N15950,N15951,
  N15952,N15953,N15954,N15955,N15956,N15957,N15958,N15959,N15960,N15961,N15962,
  N15963,N15964,N15965,N15966,N15967,N15968,N15969,N15970,N15971,N15972,N15973,
  N15974,N15975,N15976,N15977,N15978,N15979,N15980,N15981,N15982,N15983,N15984,N15985,
  N15986,N15987,N15988,N15989,N15990,N15991,N15992,N15993,N15994,N15995,N15996,
  N15997,N15998,N15999,N16000,N16001,N16002,N16003,N16004,N16005,N16006,N16007,N16008,
  N16009,N16010,N16011,N16012,N16013,N16014,N16015,N16016,N16017,N16018,N16019,
  N16020,N16021,N16022,N16023,N16024,N16025,N16026,N16027,N16028,N16029,N16030,N16031,
  N16032,N16033,N16034,N16035,N16036,N16037,N16038,N16039,N16040,N16041,N16042,
  N16043,N16044,N16045,N16046,N16047,N16048,N16049,N16050,N16051,N16052,N16053,
  N16054,N16055,N16056,N16057,N16058,N16059,N16060,N16061,N16062,N16063,N16064,N16065,
  N16066,N16067,N16068,N16069,N16070,N16071,N16072,N16073,N16074,N16075,N16076,
  N16077,N16078,N16079,N16080,N16081,N16082,N16083,N16084,N16085,N16086,N16087,N16088,
  N16089,N16090,N16091,N16092,N16093,N16094,N16095,N16096,N16097,N16098,N16099,
  N16100,N16101,N16102,N16103,N16104,N16105,N16106,N16107,N16108,N16109,N16110,N16111,
  N16112,N16113,N16114,N16115,N16116,N16117,N16118,N16119,N16120,N16121,N16122,
  N16123,N16124,N16125,N16126,N16127,N16128,N16129,N16130,N16131,N16132,N16133,
  N16134,N16135,N16136,N16137,N16138,N16139,N16140,N16141,N16142,N16143,N16144,N16145,
  N16146,N16147,N16148,N16149,N16150,N16151,N16152,N16153,N16154,N16155,N16156,
  N16157,N16158,N16159,N16160,N16161,N16162,N16163,N16164,N16165,N16166,N16167,N16168,
  N16169,N16170,N16171,N16172,N16173,N16174,N16175,N16176,N16177,N16178,N16179,
  N16180,N16181,N16182,N16183,N16184,N16185,N16186,N16187,N16188,N16189,N16190,N16191,
  N16192,N16193,N16194,N16195,N16196,N16197,N16198,N16199,N16200,N16201,N16202,
  N16203,N16204,N16205,N16206,N16207,N16208,N16209,N16210,N16211,N16212,N16213,
  N16214,N16215,N16216,N16217,N16218,N16219,N16220,N16221,N16222,N16223,N16224,N16225,
  N16226,N16227,N16228,N16229,N16230,N16231,N16232,N16233,N16234,N16235,N16236,
  N16237,N16238,N16239,N16240,N16241,N16242,N16243,N16244,N16245,N16246,N16247,N16248,
  N16249,N16250,N16251,N16252,N16253,N16254,N16255,N16256,N16257,N16258,N16259,
  N16260,N16261,N16262,N16263,N16264,N16265,N16266,N16267,N16268,N16269,N16270,N16271,
  N16272,N16273,N16274,N16275,N16276,N16277,N16278,N16279,N16280,N16281,N16282,
  N16283,N16284,N16285,N16286,N16287,N16288,N16289,N16290,N16291,N16292,N16293,
  N16294,N16295,N16296,N16297,N16298,N16299,N16300,N16301,N16302,N16303,N16304,N16305,
  N16306,N16307,N16308,N16309,N16310,N16311,N16312,N16313,N16314,N16315,N16316,
  N16317,N16318,N16319,N16320,N16321,N16322,N16323,N16324,N16325,N16326,N16327,N16328,
  N16329,N16330,N16331,N16332,N16333,N16334,N16335,N16336,N16337,N16338,N16339,
  N16340,N16341,N16342,N16343,N16344,N16345,N16346,N16347,N16348,N16349,N16350,N16351,
  N16352,N16353,N16354,N16355,N16356,N16357,N16358,N16359,N16360,N16361,N16362,
  N16363,N16364,N16365,N16366,N16367,N16368,N16369,N16370,N16371,N16372,N16373,
  N16374,N16375,N16376,N16377,N16378,N16379,N16380,N16381,N16382,N16383,N16384,N16385,
  N16386,N16387,N16388,N16389,N16390,N16391,N16392,N16393,N16394,N16395,N16396,
  N16397,N16398,N16399,N16400,N16401,N16402,N16403,N16404,N16405,N16406,N16407,N16408,
  N16409,N16410,N16411,N16412,N16413,N16414,N16415,N16416,N16417,N16418,N16419,
  N16420,N16421,N16422,N16423,N16424,N16425,N16426,N16427,N16428,N16429,N16430,N16431,
  N16432,N16433,N16434,N16435,N16436,N16437,N16438,N16439,N16440,N16441,N16442,
  N16443,N16444,N16445,N16446,N16447,N16448,N16449,N16450,N16451,N16452,N16453,
  N16454,N16455,N16456,N16457,N16458,N16459,N16460,N16461,N16462,N16463,N16464,N16465,
  N16466,N16467,N16468,N16469,N16470,N16471,N16472,N16473,N16474,N16475,N16476,
  N16477,N16478,N16479,N16480,N16481,N16482,N16483,N16484,N16485,N16486,N16487,N16488,
  N16489,N16490,N16491,N16492,N16493,N16494,N16495,N16496,N16497,N16498,N16499,
  N16500,N16501,N16502,N16503,N16504,N16505,N16506,N16507,N16508,N16509,N16510,N16511,
  N16512,N16513,N16514,N16515,N16516,N16517,N16518,N16519,N16520,N16521,N16522,
  N16523,N16524,N16525,N16526,N16527,N16528,N16529,N16530,N16531,N16532,N16533,
  N16534,N16535,N16536,N16537,N16538,N16539,N16540,N16541,N16542,N16543,N16544,N16545,
  N16546,N16547,N16548,N16549,N16550,N16551,N16552,N16553,N16554,N16555,N16556,
  N16557,N16558,N16559,N16560,N16561,N16562,N16563,N16564,N16565,N16566,N16567,N16568,
  N16569,N16570,N16571,N16572,N16573,N16574,N16575,N16576,N16577,N16578,N16579,
  N16580,N16581,N16582,N16583,N16584,N16585,N16586,N16587,N16588,N16589,N16590,N16591,
  N16592,N16593,N16594,N16595,N16596,N16597,N16598,N16599,N16600,N16601,N16602,
  N16603,N16604,N16605,N16606,N16607,N16608,N16609,N16610,N16611,N16612,N16613,
  N16614,N16615,N16616,N16617,N16618,N16619,N16620,N16621,N16622,N16623,N16624,N16625,
  N16626,N16627,N16628,N16629,N16630,N16631,N16632,N16633,N16634,N16635,N16636,
  N16637,N16638,N16639,N16640,N16641,N16642,N16643,N16644,N16645,N16646,N16647,N16648,
  N16649,N16650,N16651,N16652,N16653,N16654,N16655,N16656,N16657,N16658,N16659,
  N16660,N16661,N16662,N16663,N16664,N16665,N16666,N16667,N16668,N16669,N16670,N16671,
  N16672,N16673,N16674,N16675,N16676,N16677,N16678,N16679,N16680,N16681,N16682,
  N16683,N16684,N16685,N16686,N16687,N16688,N16689,N16690,N16691,N16692,N16693,
  N16694,N16695,N16696,N16697,N16698,N16699,N16700,N16701,N16702,N16703,N16704,N16705,
  N16706,N16707,N16708,N16709,N16710,N16711,N16712,N16713,N16714,N16715,N16716,
  N16717,N16718,N16719,N16720,N16721,N16722,N16723,N16724,N16725,N16726,N16727,N16728,
  N16729,N16730,N16731,N16732,N16733,N16734,N16735,N16736,N16737,N16738,N16739,
  N16740,N16741,N16742,N16743,N16744,N16745,N16746,N16747,N16748,N16749,N16750,N16751,
  N16752,N16753,N16754,N16755,N16756,N16757,N16758,N16759,N16760,N16761,N16762,
  N16763,N16764,N16765,N16766,N16767,N16768,N16769,N16770,N16771,N16772,N16773,
  N16774,N16775,N16776,N16777,N16778,N16779,N16780,N16781,N16782,N16783,N16784,N16785,
  N16786,N16787,N16788,N16789,N16790,N16791,N16792,N16793,N16794,N16795,N16796,
  N16797,N16798,N16799,N16800,N16801,N16802,N16803,N16804,N16805,N16806,N16807,N16808,
  N16809,N16810,N16811,N16812,N16813,N16814,N16815,N16816,N16817,N16818,N16819,
  N16820,N16821,N16822,N16823,N16824,N16825,N16826,N16827,N16828,N16829,N16830,N16831,
  N16832,N16833,N16834,N16835,N16836,N16837,N16838,N16839,N16840,N16841,N16842,
  N16843,N16844,N16845,N16846,N16847,N16848,N16849,N16850,N16851,N16852,N16853,
  N16854,N16855,N16856,N16857,N16858,N16859,N16860,N16861,N16862,N16863,N16864,N16865,
  N16866,N16867,N16868,N16869,N16870,N16871,N16872,N16873,N16874,N16875,N16876,
  N16877,N16878,N16879,N16880,N16881,N16882,N16883,N16884,N16885,N16886,N16887,N16888,
  N16889,N16890,N16891,N16892,N16893,N16894,N16895,N16896,N16897,N16898,N16899,
  N16900,N16901,N16902,N16903,N16904,N16905,N16906,N16907,N16908,N16909,N16910,N16911,
  N16912,N16913,N16914,N16915,N16916,N16917,N16918,N16919,N16920,N16921,N16922,
  N16923,N16924,N16925,N16926,N16927,N16928,N16929,N16930,N16931,N16932,N16933,
  N16934,N16935,N16936,N16937,N16938,N16939,N16940,N16941,N16942,N16943,N16944,N16945,
  N16946,N16947,N16948,N16949,N16950,N16951,N16952,N16953,N16954,N16955,N16956,
  N16957,N16958,N16959,N16960,N16961,N16962,N16963,N16964,N16965,N16966,N16967,N16968,
  N16969,N16970,N16971,N16972,N16973,N16974,N16975,N16976,N16977,N16978,N16979,
  N16980,N16981,N16982,N16983,N16984,N16985,N16986,N16987,N16988,N16989,N16990,N16991,
  N16992,N16993,N16994,N16995,N16996,N16997,N16998,N16999,N17000,N17001,N17002,
  N17003,N17004,N17005,N17006,N17007,N17008,N17009,N17010,N17011,N17012,N17013,
  N17014,N17015,N17016,N17017,N17018,N17019,N17020,N17021,N17022,N17023,N17024,N17025,
  N17026,N17027,N17028,N17029,N17030,N17031,N17032,N17033,N17034,N17035,N17036,
  N17037,N17038,N17039,N17040,N17041,N17042,N17043,N17044,N17045,N17046,N17047,N17048,
  N17049,N17050,N17051,N17052,N17053,N17054,N17055,N17056,N17057,N17058,N17059,
  N17060,N17061,N17062,N17063,N17064,N17065,N17066,N17067,N17068,N17069,N17070,N17071,
  N17072,N17073,N17074,N17075,N17076,N17077,N17078,N17079,N17080,N17081,N17082,
  N17083,N17084,N17085,N17086,N17087,N17088,N17089,N17090,N17091,N17092,N17093,
  N17094,N17095,N17096,N17097,N17098,N17099,N17100,N17101,N17102,N17103,N17104,N17105,
  N17106,N17107,N17108,N17109,N17110,N17111,N17112,N17113,N17114,N17115,N17116,
  N17117,N17118,N17119,N17120,N17121,N17122,N17123,N17124,N17125,N17126,N17127,N17128,
  N17129,N17130,N17131,N17132,N17133,N17134,N17135,N17136,N17137,N17138,N17139,
  N17140,N17141,N17142,N17143,N17144,N17145,N17146,N17147,N17148,N17149,N17150,N17151,
  N17152,N17153,N17154,N17155,N17156,N17157,N17158,N17159,N17160,N17161,N17162,
  N17163,N17164,N17165,N17166,N17167,N17168,N17169,N17170,N17171,N17172,N17173,
  N17174,N17175,N17176,N17177,N17178,N17179,N17180,N17181,N17182,N17183,N17184,N17185,
  N17186,N17187,N17188,N17189,N17190,N17191,N17192,N17193,N17194,N17195,N17196,
  N17197,N17198,N17199,N17200,N17201,N17202,N17203,N17204,N17205,N17206,N17207,N17208,
  N17209,N17210,N17211,N17212,N17213,N17214,N17215,N17216,N17217,N17218,N17219,
  N17220,N17221,N17222,N17223,N17224,N17225,N17226,N17227,N17228,N17229,N17230,N17231,
  N17232,N17233,N17234,N17235,N17236,N17237,N17238,N17239,N17240,N17241,N17242,
  N17243,N17244,N17245,N17246,N17247,N17248,N17249,N17250,N17251,N17252,N17253,
  N17254,N17255,N17256,N17257,N17258,N17259,N17260,N17261,N17262,N17263,N17264,N17265,
  N17266,N17267,N17268,N17269,N17270,N17271,N17272,N17273,N17274,N17275,N17276,
  N17277,N17278,N17279,N17280,N17281,N17282,N17283,N17284,N17285,N17286,N17287,N17288,
  N17289,N17290,N17291,N17292,N17293,N17294,N17295,N17296,N17297,N17298,N17299,
  N17300,N17301,N17302,N17303,N17304,N17305,N17306,N17307,N17308,N17309,N17310,N17311,
  N17312,N17313,N17314,N17315,N17316,N17317,N17318,N17319,N17320,N17321,N17322,
  N17323,N17324,N17325,N17326,N17327,N17328,N17329,N17330,N17331,N17332,N17333,
  N17334,N17335,N17336,N17337,N17338,N17339,N17340,N17341,N17342,N17343,N17344,N17345,
  N17346,N17347,N17348,N17349,N17350,N17351,N17352,N17353,N17354,N17355,N17356,
  N17357,N17358,N17359,N17360,N17361,N17362,N17363,N17364,N17365,N17366,N17367,N17368,
  N17369,N17370,N17371,N17372,N17373,N17374,N17375,N17376,N17377,N17378,N17379,
  N17380,N17381,N17382,N17383,N17384,N17385,N17386,N17387,N17388,N17389,N17390,N17391,
  N17392,N17393,N17394,N17395,N17396,N17397,N17398,N17399,N17400,N17401,N17402,
  N17403,N17404,N17405,N17406,N17407,N17408,N17409,N17410,N17411,N17412,N17413,
  N17414,N17415,N17416,N17417,N17418,N17419,N17420,N17421,N17422,N17423,N17424,N17425,
  N17426,N17427,N17428,N17429,N17430,N17431,N17432,N17433,N17434,N17435,N17436,
  N17437,N17438,N17439,N17440,N17441,N17442,N17443,N17444,N17445,N17446,N17447,N17448,
  N17449,N17450,N17451,N17452,N17453,N17454,N17455,N17456,N17457,N17458,N17459,
  N17460,N17461,N17462,N17463,N17464,N17465,N17466,N17467,N17468,N17469,N17470,N17471,
  N17472,N17473,N17474,N17475,N17476,N17477,N17478,N17479,N17480,N17481,N17482,
  N17483,N17484,N17485,N17486,N17487,N17488,N17489,N17490,N17491,N17492,N17493,
  N17494,N17495,N17496,N17497,N17498,N17499,N17500,N17501,N17502,N17503,N17504,N17505,
  N17506,N17507,N17508,N17509,N17510,N17511,N17512,N17513,N17514,N17515,N17516,
  N17517,N17518,N17519,N17520,N17521,N17522,N17523,N17524,N17525,N17526,N17527,N17528,
  N17529,N17530,N17531,N17532,N17533,N17534,N17535,N17536,N17537,N17538,N17539,
  N17540,N17541,N17542,N17543,N17544,N17545,N17546,N17547,N17548,N17549,N17550,N17551,
  N17552,N17553,N17554,N17555,N17556,N17557,N17558,N17559,N17560,N17561,N17562,
  N17563,N17564,N17565,N17566,N17567,N17568,N17569,N17570,N17571,N17572,N17573,
  N17574,N17575,N17576,N17577,N17578,N17579,N17580,N17581,N17582,N17583,N17584,N17585,
  N17586,N17587,N17588,N17589,N17590,N17591,N17592,N17593,N17594,N17595,N17596,
  N17597,N17598,N17599,N17600,N17601,N17602,N17603,N17604,N17605,N17606,N17607,N17608,
  N17609,N17610,N17611,N17612,N17613,N17614,N17615,N17616,N17617,N17618,N17619,
  N17620,N17621,N17622,N17623,N17624,N17625,N17626,N17627,N17628,N17629,N17630,N17631,
  N17632,N17633,N17634,N17635,N17636,N17637,N17638,N17639,N17640,N17641,N17642,
  N17643,N17644,N17645,N17646,N17647,N17648,N17649,N17650,N17651,N17652,N17653,
  N17654,N17655,N17656,N17657,N17658,N17659,N17660,N17661,N17662,N17663,N17664,N17665,
  N17666,N17667,N17668,N17669,N17670,N17671,N17672,N17673,N17674,N17675,N17676,
  N17677,N17678,N17679,N17680,N17681,N17682,N17683,N17684,N17685,N17686,N17687,N17688,
  N17689,N17690,N17691,N17692,N17693,N17694,N17695,N17696,N17697,N17698,N17699,
  N17700,N17701,N17702,N17703,N17704,N17705,N17706,N17707,N17708,N17709,N17710,N17711,
  N17712,N17713,N17714,N17715,N17716,N17717,N17718,N17719,N17720,N17721,N17722,
  N17723,N17724,N17725,N17726,N17727,N17728,N17729,N17730,N17731,N17732,N17733,
  N17734,N17735,N17736,N17737,N17738,N17739,N17740,N17741,N17742,N17743,N17744,N17745,
  N17746,N17747,N17748,N17749,N17750,N17751,N17752,N17753,N17754,N17755,N17756,
  N17757,N17758,N17759,N17760,N17761,N17762,N17763,N17764,N17765,N17766,N17767,N17768,
  N17769,N17770,N17771,N17772,N17773,N17774,N17775,N17776,N17777,N17778,N17779,
  N17780,N17781,N17782,N17783,N17784,N17785,N17786,N17787,N17788,N17789,N17790,N17791,
  N17792,N17793,N17794,N17795,N17796,N17797,N17798,N17799,N17800,N17801,N17802,
  N17803,N17804,N17805,N17806,N17807,N17808,N17809,N17810,N17811,N17812,N17813,
  N17814,N17815,N17816,N17817,N17818,N17819,N17820,N17821,N17822,N17823,N17824,N17825,
  N17826,N17827,N17828,N17829,N17830,N17831,N17832,N17833,N17834,N17835,N17836,
  N17837,N17838,N17839,N17840,N17841,N17842,N17843,N17844,N17845,N17846,N17847,N17848,
  N17849,N17850,N17851,N17852,N17853,N17854,N17855,N17856,N17857,N17858,N17859,
  N17860,N17861,N17862,N17863,N17864,N17865,N17866,N17867,N17868,N17869,N17870,N17871,
  N17872,N17873,N17874,N17875,N17876,N17877,N17878,N17879,N17880,N17881,N17882,
  N17883,N17884,N17885,N17886,N17887,N17888,N17889,N17890,N17891,N17892,N17893,
  N17894,N17895,N17896,N17897,N17898,N17899,N17900,N17901,N17902,N17903,N17904,N17905,
  N17906,N17907,N17908,N17909,N17910,N17911,N17912,N17913,N17914,N17915,N17916,
  N17917,N17918,N17919,N17920,N17921,N17922,N17923,N17924,N17925,N17926,N17927,N17928,
  N17929,N17930,N17931,N17932,N17933,N17934,N17935,N17936,N17937,N17938,N17939,
  N17940,N17941,N17942,N17943,N17944,N17945,N17946,N17947,N17948,N17949,N17950,N17951,
  N17952,N17953,N17954,N17955,N17956,N17957,N17958,N17959,N17960,N17961,N17962,
  N17963,N17964,N17965,N17966,N17967,N17968,N17969,N17970,N17971,N17972,N17973,
  N17974,N17975,N17976,N17977,N17978,N17979,N17980,N17981,N17982,N17983,N17984,N17985,
  N17986,N17987,N17988,N17989,N17990,N17991,N17992,N17993,N17994,N17995,N17996,
  N17997,N17998,N17999,N18000,N18001,N18002,N18003,N18004,N18005,N18006,N18007,N18008,
  N18009,N18010,N18011,N18012,N18013,N18014,N18015,N18016,N18017,N18018,N18019,
  N18020,N18021,N18022,N18023,N18024,N18025,N18026,N18027,N18028,N18029,N18030,N18031,
  N18032,N18033,N18034,N18035,N18036,N18037,N18038,N18039,N18040,N18041,N18042,
  N18043,N18044,N18045,N18046,N18047,N18048,N18049,N18050,N18051,N18052,N18053,
  N18054,N18055,N18056,N18057,N18058,N18059,N18060,N18061,N18062,N18063,N18064,N18065,
  N18066,N18067,N18068,N18069,N18070,N18071,N18072,N18073,N18074,N18075,N18076,
  N18077,N18078,N18079,N18080,N18081,N18082,N18083,N18084,N18085,N18086,N18087,N18088,
  N18089,N18090,N18091,N18092,N18093,N18094,N18095,N18096,N18097,N18098,N18099,
  N18100,N18101,N18102,N18103,N18104,N18105,N18106,N18107,N18108,N18109,N18110,N18111,
  N18112,N18113,N18114,N18115,N18116,N18117,N18118,N18119,N18120,N18121,N18122,
  N18123,N18124,N18125,N18126,N18127,N18128,N18129,N18130,N18131,N18132,N18133,
  N18134,N18135,N18136,N18137,N18138,N18139,N18140,N18141,N18142,N18143,N18144,N18145,
  N18146,N18147,N18148,N18149,N18150,N18151,N18152,N18153,N18154,N18155,N18156,
  N18157,N18158,N18159,N18160,N18161,N18162,N18163,N18164,N18165,N18166,N18167,N18168,
  N18169,N18170,N18171,N18172,N18173,N18174,N18175,N18176,N18177,N18178,N18179,
  N18180,N18181,N18182,N18183,N18184,N18185,N18186,N18187,N18188,N18189,N18190,N18191,
  N18192,N18193,N18194,N18195,N18196,N18197,N18198,N18199,N18200,N18201,N18202,
  N18203,N18204,N18205,N18206,N18207,N18208,N18209,N18210,N18211,N18212,N18213,
  N18214,N18215,N18216,N18217,N18218,N18219,N18220,N18221,N18222,N18223,N18224,N18225,
  N18226,N18227,N18228,N18229,N18230,N18231,N18232,N18233,N18234,N18235,N18236,
  N18237,N18238,N18239,N18240,N18241,N18242,N18243,N18244,N18245,N18246,N18247,N18248,
  N18249,N18250,N18251,N18252,N18253,N18254,N18255,N18256,N18257,N18258,N18259,
  N18260,N18261,N18262,N18263,N18264,N18265,N18266,N18267,N18268,N18269,N18270,N18271,
  N18272,N18273,N18274,N18275,N18276,N18277,N18278,N18279,N18280,N18281,N18282,
  N18283,N18284,N18285,N18286,N18287,N18288,N18289,N18290,N18291,N18292,N18293,
  N18294,N18295,N18296,N18297,N18298,N18299,N18300,N18301,N18302,N18303,N18304,N18305,
  N18306,N18307,N18308,N18309,N18310,N18311,N18312,N18313,N18314,N18315,N18316,
  N18317,N18318,N18319,N18320,N18321,N18322,N18323,N18324,N18325,N18326,N18327,N18328,
  N18329,N18330,N18331,N18332,N18333,N18334,N18335,N18336,N18337,N18338,N18339,
  N18340,N18341,N18342,N18343,N18344,N18345,N18346,N18347,N18348,N18349,N18350,N18351,
  N18352,N18353,N18354,N18355,N18356,N18357,N18358,N18359,N18360,N18361,N18362,
  N18363,N18364,N18365,N18366,N18367,N18368,N18369,N18370,N18371,N18372,N18373,
  N18374,N18375,N18376,N18377,N18378,N18379,N18380,N18381,N18382,N18383,N18384,N18385,
  N18386,N18387,N18388,N18389,N18390,N18391,N18392,N18393,N18394,N18395,N18396,
  N18397,N18398,N18399,N18400,N18401,N18402,N18403,N18404,N18405,N18406,N18407,N18408,
  N18409,N18410,N18411,N18412,N18413,N18414,N18415,N18416,N18417,N18418,N18419,
  N18420,N18421,N18422,N18423,N18424,N18425,N18426,N18427,N18428,N18429,N18430,N18431,
  N18432,N18433,N18434,N18435,N18436,N18437,N18438,N18439,N18440,N18441,N18442,
  N18443,N18444,N18445,N18446,N18447,N18448,N18449,N18450,N18451,N18452,N18453,
  N18454,N18455,N18456,N18457,N18458,N18459,N18460,N18461,N18462,N18463,N18464,N18465,
  N18466,N18467,N18468,N18469,N18470,N18471,N18472,N18473,N18474,N18475,N18476,
  N18477,N18478,N18479,N18480,N18481,N18482,N18483,N18484,N18485,N18486,N18487,N18488,
  N18489,N18490,N18491,N18492,N18493,N18494,N18495,N18496,N18497,N18498,N18499,
  N18500,N18501,N18502,N18503,N18504,N18505,N18506,N18507,N18508,N18509,N18510,N18511,
  N18512,N18513,N18514,N18515,N18516,N18517,N18518,N18519,N18520,N18521,N18522,
  N18523,N18524,N18525,N18526,N18527,N18528,N18529,N18530,N18531,N18532,N18533,
  N18534,N18535,N18536,N18537,N18538,N18539,N18540,N18541,N18542,N18543,N18544,N18545,
  N18546,N18547,N18548,N18549,N18550,N18551,N18552,N18553,N18554,N18555,N18556,
  N18557,N18558,N18559,N18560,N18561,N18562,N18563,N18564,N18565,N18566,N18567,N18568,
  N18569,N18570,N18571,N18572,N18573,N18574,N18575,N18576,N18577,N18578,N18579,
  N18580,N18581,N18582,N18583,N18584,N18585,N18586,N18587,N18588,N18589,N18590,N18591,
  N18592,N18593,N18594,N18595,N18596,N18597,N18598,N18599,N18600,N18601,N18602,
  N18603,N18604,N18605,N18606,N18607,N18608,N18609,N18610,N18611,N18612,N18613,
  N18614,N18615,N18616,N18617,N18618,N18619,N18620,N18621,N18622,N18623,N18624,N18625,
  N18626,N18627,N18628,N18629,N18630,N18631,N18632,N18633,N18634,N18635,N18636,
  N18637,N18638,N18639,N18640,N18641,N18642,N18643,N18644,N18645,N18646,N18647,N18648,
  N18649,N18650,N18651,N18652,N18653,N18654,N18655,N18656,N18657,N18658,N18659,
  N18660,N18661,N18662,N18663,N18664,N18665,N18666,N18667,N18668,N18669,N18670,N18671,
  N18672,N18673,N18674,N18675,N18676,N18677,N18678,N18679,N18680,N18681,N18682,
  N18683,N18684,N18685,N18686,N18687,N18688,N18689,N18690,N18691,N18692,N18693,
  N18694,N18695,N18696,N18697,N18698,N18699,N18700,N18701,N18702,N18703,N18704,N18705,
  N18706,N18707,N18708,N18709,N18710,N18711,N18712,N18713,N18714,N18715,N18716,
  N18717,N18718,N18719,N18720,N18721,N18722,N18723,N18724,N18725,N18726,N18727,N18728,
  N18729,N18730,N18731,N18732,N18733,N18734,N18735,N18736,N18737,N18738,N18739,
  N18740,N18741,N18742,N18743,N18744,N18745,N18746,N18747,N18748,N18749,N18750,N18751,
  N18752,N18753,N18754,N18755,N18756,N18757,N18758,N18759,N18760,N18761,N18762,
  N18763,N18764,N18765,N18766,N18767,N18768,N18769,N18770,N18771,N18772,N18773,
  N18774,N18775,N18776,N18777,N18778,N18779,N18780,N18781,N18782,N18783,N18784,N18785,
  N18786,N18787,N18788,N18789,N18790,N18791,N18792,N18793,N18794,N18795,N18796,
  N18797,N18798,N18799,N18800,N18801,N18802,N18803,N18804,N18805,N18806,N18807,N18808,
  N18809,N18810,N18811,N18812,N18813,N18814,N18815,N18816,N18817,N18818,N18819,
  N18820,N18821,N18822,N18823,N18824,N18825,N18826,N18827,N18828,N18829,N18830,N18831,
  N18832,N18833,N18834,N18835,N18836,N18837,N18838,N18839,N18840,N18841,N18842,
  N18843,N18844,N18845,N18846,N18847,N18848,N18849,N18850,N18851,N18852,N18853,
  N18854,N18855,N18856,N18857,N18858,N18859,N18860,N18861,N18862,N18863,N18864,N18865,
  N18866,N18867,N18868,N18869,N18870,N18871,N18872,N18873,N18874,N18875,N18876,
  N18877,N18878,N18879,N18880,N18881,N18882,N18883,N18884,N18885,N18886,N18887,N18888,
  N18889,N18890,N18891,N18892,N18893,N18894,N18895,N18896,N18897,N18898,N18899,
  N18900,N18901,N18902,N18903,N18904,N18905,N18906,N18907,N18908,N18909,N18910,N18911,
  N18912,N18913,N18914,N18915,N18916,N18917,N18918,N18919,N18920,N18921,N18922,
  N18923,N18924,N18925,N18926,N18927,N18928,N18929,N18930,N18931,N18932,N18933,
  N18934,N18935,N18936,N18937,N18938,N18939,N18940,N18941,N18942,N18943,N18944,N18945,
  N18946,N18947,N18948,N18949,N18950,N18951,N18952,N18953,N18954,N18955,N18956,
  N18957,N18958,N18959,N18960,N18961,N18962,N18963,N18964,N18965,N18966,N18967,N18968,
  N18969,N18970,N18971,N18972,N18973,N18974,N18975,N18976,N18977,N18978,N18979,
  N18980,N18981,N18982,N18983,N18984,N18985,N18986,N18987,N18988,N18989,N18990,N18991,
  N18992,N18993,N18994,N18995,N18996,N18997,N18998,N18999,N19000,N19001,N19002,
  N19003,N19004,N19005,N19006,N19007,N19008,N19009,N19010,N19011,N19012,N19013,
  N19014,N19015,N19016,N19017,N19018,N19019,N19020,N19021,N19022,N19023,N19024,N19025,
  N19026,N19027,N19028,N19029,N19030,N19031,N19032,N19033,N19034,N19035,N19036,
  N19037,N19038,N19039,N19040,N19041,N19042,N19043,N19044,N19045,N19046,N19047,N19048,
  N19049,N19050,N19051,N19052,N19053,N19054,N19055,N19056,N19057,N19058,N19059,
  N19060,N19061,N19062,N19063,N19064,N19065,N19066,N19067,N19068,N19069,N19070,N19071,
  N19072,N19073,N19074,N19075,N19076,N19077,N19078,N19079,N19080,N19081,N19082,
  N19083,N19084,N19085,N19086,N19087,N19088,N19089,N19090,N19091,N19092,N19093,
  N19094,N19095,N19096,N19097,N19098,N19099,N19100,N19101,N19102,N19103,N19104,N19105,
  N19106,N19107,N19108,N19109,N19110,N19111,N19112,N19113,N19114,N19115,N19116,
  N19117,N19118,N19119,N19120,N19121,N19122,N19123,N19124,N19125,N19126,N19127,N19128,
  N19129,N19130,N19131,N19132,N19133,N19134,N19135,N19136,N19137,N19138,N19139,
  N19140,N19141,N19142,N19143,N19144,N19145,N19146,N19147,N19148,N19149,N19150,N19151,
  N19152,N19153,N19154,N19155,N19156,N19157,N19158,N19159,N19160,N19161,N19162,
  N19163,N19164,N19165,N19166,N19167,N19168,N19169,N19170,N19171,N19172,N19173,
  N19174,N19175,N19176,N19177,N19178,N19179,N19180,N19181,N19182,N19183,N19184,N19185,
  N19186,N19187,N19188,N19189,N19190,N19191,N19192,N19193,N19194,N19195,N19196,
  N19197,N19198,N19199,N19200,N19201,N19202,N19203,N19204,N19205,N19206,N19207,N19208,
  N19209,N19210,N19211,N19212,N19213,N19214,N19215,N19216,N19217,N19218,N19219,
  N19220,N19221,N19222,N19223,N19224,N19225,N19226,N19227,N19228,N19229,N19230,N19231,
  N19232,N19233,N19234,N19235,N19236,N19237,N19238,N19239,N19240,N19241,N19242,
  N19243,N19244,N19245,N19246,N19247,N19248,N19249,N19250,N19251,N19252,N19253,
  N19254,N19255,N19256,N19257,N19258,N19259,N19260,N19261,N19262,N19263,N19264,N19265,
  N19266,N19267,N19268,N19269,N19270,N19271,N19272,N19273,N19274,N19275,N19276,
  N19277,N19278,N19279,N19280,N19281,N19282,N19283,N19284,N19285,N19286,N19287,N19288,
  N19289,N19290,N19291,N19292,N19293,N19294,N19295,N19296,N19297,N19298,N19299,
  N19300,N19301,N19302,N19303,N19304,N19305,N19306,N19307,N19308,N19309,N19310,N19311,
  N19312,N19313,N19314,N19315,N19316,N19317,N19318,N19319,N19320,N19321,N19322,
  N19323,N19324,N19325,N19326,N19327,N19328,N19329,N19330,N19331,N19332,N19333,
  N19334,N19335,N19336,N19337,N19338,N19339,N19340,N19341,N19342,N19343,N19344,N19345,
  N19346,N19347,N19348,N19349,N19350,N19351,N19352,N19353,N19354,N19355,N19356,
  N19357,N19358,N19359,N19360,N19361,N19362,N19363,N19364,N19365,N19366,N19367,N19368,
  N19369,N19370,N19371,N19372,N19373,N19374,N19375,N19376,N19377,N19378,N19379,
  N19380,N19381,N19382,N19383,N19384,N19385,N19386,N19387,N19388,N19389,N19390,N19391,
  N19392,N19393,N19394,N19395,N19396,N19397,N19398,N19399,N19400,N19401,N19402,
  N19403,N19404,N19405,N19406,N19407,N19408,N19409,N19410,N19411,N19412,N19413,
  N19414,N19415,N19416,N19417,N19418,N19419,N19420,N19421,N19422,N19423,N19424,N19425,
  N19426,N19427,N19428,N19429,N19430,N19431,N19432,N19433,N19434,N19435,N19436,
  N19437,N19438,N19439,N19440,N19441,N19442,N19443,N19444,N19445,N19446,N19447,N19448,
  N19449,N19450,N19451,N19452,N19453,N19454,N19455,N19456,N19457,N19458,N19459,
  N19460,N19461,N19462,N19463,N19464,N19465,N19466,N19467,N19468,N19469,N19470,N19471,
  N19472,N19473,N19474,N19475,N19476,N19477,N19478,N19479,N19480,N19481,N19482,
  N19483,N19484,N19485,N19486,N19487,N19488,N19489,N19490,N19491,N19492,N19493,
  N19494,N19495,N19496,N19497,N19498,N19499,N19500,N19501,N19502,N19503,N19504,N19505,
  N19506,N19507,N19508,N19509,N19510,N19511,N19512,N19513,N19514,N19515,N19516,
  N19517,N19518,N19519,N19520,N19521,N19522,N19523,N19524,N19525,N19526,N19527,N19528,
  N19529,N19530,N19531,N19532,N19533,N19534,N19535,N19536,N19537,N19538,N19539,
  N19540,N19541,N19542,N19543,N19544,N19545,N19546,N19547,N19548,N19549,N19550,N19551,
  N19552,N19553,N19554,N19555,N19556,N19557,N19558,N19559,N19560,N19561,N19562,
  N19563,N19564,N19565,N19566,N19567,N19568,N19569,N19570,N19571,N19572,N19573,
  N19574,N19575,N19576,N19577,N19578,N19579,N19580,N19581,N19582,N19583,N19584,N19585,
  N19586,N19587,N19588,N19589,N19590,N19591,N19592,N19593,N19594,N19595,N19596,
  N19597,N19598,N19599,N19600,N19601,N19602,N19603,N19604,N19605,N19606,N19607,N19608,
  N19609,N19610,N19611,N19612,N19613,N19614,N19615,N19616,N19617,N19618,N19619,
  N19620,N19621,N19622,N19623,N19624,N19625,N19626,N19627,N19628,N19629,N19630,N19631,
  N19632,N19633,N19634,N19635,N19636,N19637,N19638,N19639,N19640,N19641,N19642,
  N19643,N19644,N19645,N19646,N19647,N19648,N19649,N19650,N19651,N19652,N19653,
  N19654,N19655,N19656,N19657,N19658,N19659,N19660,N19661,N19662,N19663,N19664,N19665,
  N19666,N19667,N19668,N19669,N19670,N19671,N19672,N19673,N19674,N19675,N19676,
  N19677,N19678,N19679,N19680,N19681,N19682,N19683,N19684,N19685,N19686,N19687,N19688,
  N19689,N19690,N19691,N19692,N19693,N19694,N19695,N19696,N19697,N19698,N19699,
  N19700,N19701,N19702,N19703,N19704,N19705,N19706,N19707,N19708,N19709,N19710,N19711,
  N19712,N19713,N19714,N19715,N19716,N19717,N19718,N19719,N19720,N19721,N19722,
  N19723,N19724,N19725,N19726,N19727,N19728,N19729,N19730,N19731,N19732,N19733,
  N19734,N19735,N19736,N19737,N19738,N19739,N19740,N19741,N19742,N19743,N19744,N19745,
  N19746,N19747,N19748,N19749,N19750,N19751,N19752,N19753,N19754,N19755,N19756,
  N19757,N19758,N19759,N19760,N19761,N19762,N19763,N19764,N19765,N19766,N19767,N19768,
  N19769,N19770,N19771,N19772,N19773,N19774,N19775,N19776,N19777,N19778,N19779,
  N19780,N19781,N19782,N19783,N19784,N19785,N19786,N19787,N19788,N19789,N19790,N19791,
  N19792,N19793,N19794,N19795,N19796,N19797,N19798,N19799,N19800,N19801,N19802,
  N19803,N19804,N19805,N19806,N19807,N19808,N19809,N19810,N19811,N19812,N19813,
  N19814,N19815,N19816,N19817,N19818,N19819,N19820,N19821,N19822,N19823,N19824,N19825,
  N19826,N19827,N19828,N19829,N19830,N19831,N19832,N19833,N19834,N19835,N19836,
  N19837,N19838,N19839,N19840,N19841,N19842,N19843,N19844,N19845,N19846,N19847,N19848,
  N19849,N19850,N19851,N19852,N19853,N19854,N19855,N19856,N19857,N19858,N19859,
  N19860,N19861,N19862,N19863,N19864,N19865,N19866,N19867,N19868,N19869,N19870,N19871,
  N19872,N19873,N19874,N19875,N19876,N19877,N19878,N19879,N19880,N19881,N19882,
  N19883,N19884,N19885,N19886,N19887,N19888,N19889,N19890,N19891,N19892,N19893,
  N19894,N19895,N19896,N19897,N19898,N19899,N19900,N19901,N19902,N19903,N19904,N19905,
  N19906,N19907,N19908,N19909,N19910,N19911,N19912,N19913,N19914,N19915,N19916,
  N19917,N19918,N19919,N19920,N19921,N19922,N19923,N19924,N19925,N19926,N19927,N19928,
  N19929,N19930,N19931,N19932,N19933,N19934,N19935,N19936,N19937,N19938,N19939,
  N19940,N19941,N19942,N19943,N19944,N19945,N19946,N19947,N19948,N19949,N19950,N19951,
  N19952,N19953,N19954,N19955,N19956,N19957,N19958,N19959,N19960,N19961,N19962,
  N19963,N19964,N19965,N19966,N19967,N19968,N19969,N19970,N19971,N19972,N19973,
  N19974,N19975,N19976,N19977,N19978,N19979,N19980,N19981,N19982,N19983,N19984,N19985,
  N19986,N19987,N19988,N19989,N19990,N19991,N19992,N19993,N19994,N19995,N19996,
  N19997,N19998,N19999,N20000,N20001,N20002,N20003,N20004,N20005,N20006,N20007,N20008,
  N20009,N20010,N20011,N20012,N20013,N20014,N20015,N20016,N20017,N20018,N20019,
  N20020,N20021,N20022,N20023,N20024,N20025,N20026,N20027,N20028,N20029,N20030,N20031,
  N20032,N20033,N20034,N20035,N20036,N20037,N20038,N20039,N20040,N20041,N20042,
  N20043,N20044,N20045,N20046,N20047,N20048,N20049,N20050,N20051,N20052,N20053,
  N20054,N20055,N20056,N20057,N20058,N20059,N20060,N20061,N20062,N20063,N20064,N20065,
  N20066,N20067,N20068,N20069,N20070,N20071,N20072,N20073,N20074,N20075,N20076,
  N20077,N20078,N20079,N20080,N20081,N20082,N20083,N20084,N20085,N20086,N20087,N20088,
  N20089,N20090,N20091,N20092,N20093,N20094,N20095,N20096,N20097,N20098,N20099,
  N20100,N20101,N20102,N20103,N20104,N20105,N20106,N20107,N20108,N20109,N20110,N20111,
  N20112,N20113,N20114,N20115,N20116,N20117,N20118,N20119,N20120,N20121,N20122,
  N20123,N20124,N20125,N20126,N20127,N20128,N20129,N20130,N20131,N20132,N20133,
  N20134,N20135,N20136,N20137,N20138,N20139,N20140,N20141,N20142,N20143,N20144,N20145,
  N20146,N20147,N20148,N20149,N20150,N20151,N20152,N20153,N20154,N20155,N20156,
  N20157,N20158,N20159,N20160,N20161,N20162,N20163,N20164,N20165,N20166,N20167,N20168,
  N20169,N20170,N20171,N20172,N20173,N20174,N20175,N20176,N20177,N20178,N20179,
  N20180,N20181,N20182,N20183,N20184,N20185,N20186,N20187,N20188,N20189,N20190,N20191,
  N20192,N20193,N20194,N20195,N20196,N20197,N20198,N20199,N20200,N20201,N20202,
  N20203,N20204,N20205,N20206,N20207,N20208,N20209,N20210,N20211,N20212,N20213,
  N20214,N20215,N20216,N20217,N20218,N20219,N20220,N20221,N20222,N20223,N20224,N20225,
  N20226,N20227,N20228,N20229,N20230,N20231,N20232,N20233,N20234,N20235,N20236,
  N20237,N20238,N20239,N20240,N20241,N20242,N20243,N20244,N20245,N20246,N20247,N20248,
  N20249,N20250,N20251,N20252,N20253,N20254,N20255,N20256,N20257,N20258,N20259,
  N20260,N20261,N20262,N20263,N20264,N20265,N20266,N20267,N20268,N20269,N20270,N20271,
  N20272,N20273,N20274,N20275,N20276,N20277,N20278,N20279,N20280,N20281,N20282,
  N20283,N20284,N20285,N20286,N20287,N20288,N20289,N20290,N20291,N20292,N20293,
  N20294,N20295,N20296,N20297,N20298,N20299,N20300,N20301,N20302,N20303,N20304,N20305,
  N20306,N20307,N20308,N20309,N20310,N20311,N20312,N20313,N20314,N20315,N20316,
  N20317,N20318,N20319,N20320,N20321,N20322,N20323,N20324,N20325,N20326,N20327,N20328,
  N20329,N20330,N20331,N20332,N20333,N20334,N20335,N20336,N20337,N20338,N20339,
  N20340,N20341,N20342,N20343,N20344,N20345,N20346,N20347,N20348,N20349,N20350,N20351,
  N20352,N20353,N20354,N20355,N20356,N20357,N20358,N20359,N20360,N20361,N20362,
  N20363,N20364,N20365,N20366,N20367,N20368,N20369,N20370,N20371,N20372,N20373,
  N20374,N20375,N20376,N20377,N20378,N20379,N20380,N20381,N20382,N20383,N20384,N20385,
  N20386,N20387,N20388,N20389,N20390,N20391,N20392,N20393,N20394,N20395,N20396,
  N20397,N20398,N20399,N20400,N20401,N20402,N20403,N20404,N20405,N20406,N20407,N20408,
  N20409,N20410,N20411,N20412,N20413,N20414,N20415,N20416,N20417,N20418,N20419,
  N20420,N20421,N20422,N20423,N20424,N20425,N20426,N20427,N20428,N20429,N20430,N20431,
  N20432,N20433,N20434,N20435,N20436,N20437,N20438,N20439,N20440,N20441,N20442,
  N20443,N20444,N20445,N20446,N20447,N20448,N20449,N20450,N20451,N20452,N20453,
  N20454,N20455,N20456,N20457,N20458,N20459,N20460,N20461,N20462,N20463,N20464,N20465,
  N20466,N20467,N20468,N20469,N20470,N20471,N20472,N20473,N20474,N20475,N20476,
  N20477,N20478,N20479,N20480,N20481,N20482,N20483,N20484,N20485,N20486,N20487,N20488,
  N20489,N20490,N20491,N20492,N20493,N20494,N20495,N20496,N20497,N20498,N20499,
  N20500,N20501,N20502,N20503,N20504,N20505,N20506,N20507,N20508,N20509,N20510,N20511,
  N20512,N20513,N20514,N20515,N20516,N20517,N20518,N20519,N20520,N20521,N20522,
  N20523,N20524,N20525,N20526,N20527,N20528,N20529,N20530,N20531,N20532,N20533,
  N20534,N20535,N20536,N20537,N20538,N20539,N20540,N20541,N20542,N20543,N20544,N20545,
  N20546,N20547,N20548,N20549,N20550,N20551,N20552,N20553,N20554,N20555,N20556,
  N20557,N20558,N20559,N20560,N20561,N20562,N20563,N20564,N20565,N20566,N20567,N20568,
  N20569,N20570,N20571,N20572,N20573,N20574,N20575,N20576,N20577,N20578,N20579,
  N20580,N20581,N20582,N20583,N20584,N20585,N20586,N20587,N20588,N20589,N20590,N20591,
  N20592,N20593,N20594,N20595,N20596,N20597,N20598,N20599,N20600,N20601,N20602,
  N20603,N20604,N20605,N20606,N20607,N20608,N20609,N20610,N20611,N20612,N20613,
  N20614,N20615,N20616,N20617,N20618,N20619,N20620,N20621,N20622,N20623,N20624,N20625,
  N20626,N20627,N20628,N20629,N20630,N20631,N20632,N20633,N20634,N20635,N20636,
  N20637,N20638,N20639,N20640,N20641,N20642,N20643,N20644,N20645,N20646,N20647,N20648,
  N20649,N20650,N20651,N20652,N20653,N20654,N20655,N20656,N20657,N20658,N20659,
  N20660,N20661,N20662,N20663,N20664,N20665,N20666,N20667,N20668,N20669,N20670,N20671,
  N20672,N20673,N20674,N20675,N20676,N20677,N20678,N20679,N20680,N20681,N20682,
  N20683,N20684,N20685,N20686,N20687,N20688,N20689,N20690,N20691,N20692,N20693,
  N20694,N20695,N20696,N20697,N20698,N20699,N20700,N20701,N20702,N20703,N20704,N20705,
  N20706,N20707,N20708,N20709,N20710,N20711,N20712,N20713,N20714,N20715,N20716,
  N20717,N20718,N20719,N20720,N20721,N20722,N20723,N20724,N20725,N20726,N20727,N20728,
  N20729,N20730,N20731,N20732,N20733,N20734,N20735,N20736,N20737,N20738,N20739,
  N20740,N20741,N20742,N20743,N20744,N20745,N20746,N20747,N20748,N20749,N20750,N20751,
  N20752,N20753,N20754,N20755,N20756,N20757,N20758,N20759,N20760,N20761,N20762,
  N20763,N20764,N20765,N20766,N20767,N20768,N20769,N20770,N20771,N20772,N20773,
  N20774,N20775,N20776,N20777,N20778,N20779,N20780,N20781,N20782,N20783,N20784,N20785,
  N20786,N20787,N20788,N20789,N20790,N20791,N20792,N20793,N20794,N20795,N20796,
  N20797,N20798,N20799,N20800,N20801,N20802,N20803,N20804,N20805,N20806,N20807,N20808,
  N20809,N20810,N20811,N20812,N20813,N20814,N20815,N20816,N20817,N20818,N20819,
  N20820,N20821,N20822,N20823,N20824,N20825,N20826,N20827,N20828,N20829,N20830,N20831,
  N20832,N20833,N20834,N20835,N20836,N20837,N20838,N20839,N20840,N20841,N20842,
  N20843,N20844,N20845,N20846,N20847,N20848,N20849,N20850,N20851,N20852,N20853,
  N20854,N20855,N20856,N20857,N20858,N20859,N20860,N20861,N20862,N20863,N20864,N20865,
  N20866,N20867,N20868,N20869,N20870,N20871,N20872,N20873,N20874,N20875,N20876,
  N20877,N20878,N20879,N20880,N20881,N20882,N20883,N20884,N20885,N20886,N20887,N20888,
  N20889,N20890,N20891,N20892,N20893,N20894,N20895,N20896,N20897,N20898,N20899,
  N20900,N20901,N20902,N20903,N20904,N20905,N20906,N20907,N20908,N20909,N20910,N20911,
  N20912,N20913,N20914,N20915,N20916,N20917,N20918,N20919,N20920,N20921,N20922,
  N20923,N20924,N20925,N20926,N20927,N20928,N20929,N20930,N20931,N20932,N20933,
  N20934,N20935,N20936,N20937,N20938,N20939,N20940,N20941,N20942,N20943,N20944,N20945,
  N20946,N20947,N20948,N20949,N20950,N20951,N20952,N20953,N20954,N20955,N20956,
  N20957,N20958,N20959,N20960,N20961,N20962,N20963,N20964,N20965,N20966,N20967,N20968,
  N20969,N20970,N20971,N20972,N20973,N20974,N20975,N20976,N20977,N20978,N20979,
  N20980,N20981,N20982,N20983,N20984,N20985,N20986,N20987,N20988,N20989,N20990,N20991,
  N20992,N20993,N20994,N20995,N20996,N20997,N20998,N20999,N21000,N21001,N21002,
  N21003,N21004,N21005,N21006,N21007,N21008,N21009,N21010,N21011,N21012,N21013,
  N21014,N21015,N21016,N21017,N21018,N21019,N21020,N21021,N21022,N21023,N21024,N21025,
  N21026,N21027,N21028,N21029,N21030,N21031,N21032,N21033,N21034,N21035,N21036,
  N21037,N21038,N21039,N21040,N21041,N21042,N21043,N21044,N21045,N21046,N21047,N21048,
  N21049,N21050,N21051,N21052,N21053,N21054,N21055,N21056,N21057,N21058,N21059,
  N21060,N21061,N21062,N21063,N21064,N21065,N21066,N21067,N21068,N21069,N21070,N21071,
  N21072,N21073,N21074,N21075,N21076,N21077,N21078,N21079,N21080,N21081,N21082,
  N21083,N21084,N21085,N21086,N21087,N21088,N21089,N21090,N21091,N21092,N21093,
  N21094,N21095,N21096,N21097,N21098,N21099,N21100,N21101,N21102,N21103,N21104,N21105,
  N21106,N21107,N21108,N21109,N21110,N21111,N21112,N21113,N21114,N21115,N21116,
  N21117,N21118,N21119,N21120,N21121,N21122,N21123,N21124,N21125,N21126,N21127,N21128,
  N21129,N21130,N21131,N21132,N21133,N21134,N21135,N21136,N21137,N21138,N21139,
  N21140,N21141,N21142,N21143,N21144,N21145,N21146,N21147,N21148,N21149,N21150,N21151,
  N21152,N21153,N21154,N21155,N21156,N21157,N21158,N21159,N21160,N21161,N21162,
  N21163,N21164,N21165,N21166,N21167,N21168,N21169,N21170,N21171,N21172,N21173,
  N21174,N21175,N21176,N21177,N21178,N21179,N21180,N21181,N21182,N21183,N21184,N21185,
  N21186,N21187,N21188,N21189,N21190,N21191,N21192,N21193,N21194,N21195,N21196,
  N21197,N21198,N21199,N21200,N21201,N21202,N21203,N21204,N21205,N21206,N21207,N21208,
  N21209,N21210,N21211,N21212,N21213,N21214,N21215,N21216,N21217,N21218,N21219,
  N21220,N21221,N21222,N21223,N21224,N21225,N21226,N21227,N21228,N21229,N21230,N21231,
  N21232,N21233,N21234,N21235,N21236,N21237,N21238,N21239,N21240,N21241,N21242,
  N21243,N21244,N21245,N21246,N21247,N21248,N21249,N21250,N21251,N21252,N21253,
  N21254,N21255,N21256,N21257,N21258,N21259,N21260,N21261,N21262,N21263,N21264,N21265,
  N21266,N21267,N21268,N21269,N21270,N21271,N21272,N21273,N21274,N21275,N21276,
  N21277,N21278,N21279,N21280,N21281,N21282,N21283,N21284,N21285,N21286,N21287,N21288,
  N21289,N21290,N21291,N21292,N21293,N21294,N21295,N21296,N21297,N21298,N21299,
  N21300,N21301,N21302,N21303,N21304,N21305,N21306,N21307,N21308,N21309,N21310,N21311,
  N21312,N21313,N21314,N21315,N21316,N21317,N21318,N21319,N21320,N21321,N21322,
  N21323,N21324,N21325,N21326,N21327,N21328,N21329,N21330,N21331,N21332,N21333,
  N21334,N21335,N21336,N21337,N21338,N21339,N21340,N21341,N21342,N21343,N21344,N21345,
  N21346,N21347,N21348,N21349,N21350,N21351,N21352,N21353,N21354,N21355,N21356,
  N21357,N21358,N21359,N21360,N21361,N21362,N21363,N21364,N21365,N21366,N21367,N21368,
  N21369,N21370,N21371,N21372,N21373,N21374,N21375,N21376,N21377,N21378,N21379,
  N21380,N21381,N21382,N21383,N21384,N21385,N21386,N21387,N21388,N21389,N21390,N21391,
  N21392,N21393,N21394,N21395,N21396,N21397,N21398,N21399,N21400,N21401,N21402,
  N21403,N21404,N21405,N21406,N21407,N21408,N21409,N21410,N21411,N21412,N21413,
  N21414,N21415,N21416,N21417,N21418,N21419,N21420,N21421,N21422,N21423,N21424,N21425,
  N21426,N21427,N21428,N21429,N21430,N21431,N21432,N21433,N21434,N21435,N21436,
  N21437,N21438,N21439,N21440,N21441,N21442,N21443,N21444,N21445,N21446,N21447,N21448,
  N21449,N21450,N21451,N21452,N21453,N21454,N21455,N21456,N21457,N21458,N21459,
  N21460,N21461,N21462,N21463,N21464,N21465,N21466,N21467,N21468,N21469,N21470,N21471,
  N21472,N21473,N21474,N21475,N21476,N21477,N21478,N21479,N21480,N21481,N21482,
  N21483,N21484,N21485,N21486,N21487,N21488,N21489,N21490,N21491,N21492,N21493,
  N21494,N21495,N21496,N21497,N21498,N21499,N21500,N21501,N21502,N21503,N21504,N21505,
  N21506,N21507,N21508,N21509,N21510,N21511,N21512,N21513,N21514,N21515,N21516,
  N21517,N21518,N21519,N21520,N21521,N21522,N21523,N21524,N21525,N21526,N21527,N21528,
  N21529,N21530,N21531,N21532,N21533,N21534,N21535,N21536,N21537,N21538,N21539,
  N21540,N21541,N21542,N21543,N21544,N21545,N21546,N21547,N21548,N21549,N21550,N21551,
  N21552,N21553,N21554,N21555,N21556,N21557,N21558,N21559,N21560,N21561,N21562,
  N21563,N21564,N21565,N21566,N21567,N21568,N21569,N21570,N21571,N21572,N21573,
  N21574,N21575,N21576,N21577,N21578,N21579,N21580,N21581,N21582,N21583,N21584,N21585,
  N21586,N21587,N21588,N21589,N21590,N21591,N21592,N21593,N21594,N21595,N21596,
  N21597,N21598,N21599,N21600,N21601,N21602,N21603,N21604,N21605,N21606,N21607,N21608,
  N21609,N21610,N21611,N21612,N21613,N21614,N21615,N21616,N21617,N21618,N21619,
  N21620,N21621,N21622,N21623,N21624,N21625,N21626,N21627,N21628,N21629,N21630,N21631,
  N21632,N21633,N21634,N21635,N21636,N21637,N21638,N21639,N21640,N21641,N21642,
  N21643,N21644,N21645,N21646,N21647,N21648,N21649,N21650,N21651,N21652,N21653,
  N21654,N21655,N21656,N21657,N21658,N21659,N21660,N21661,N21662,N21663,N21664,N21665,
  N21666,N21667,N21668,N21669,N21670,N21671,N21672,N21673,N21674,N21675,N21676,
  N21677,N21678,N21679,N21680,N21681,N21682,N21683,N21684,N21685,N21686,N21687,N21688,
  N21689,N21690,N21691,N21692,N21693,N21694,N21695,N21696,N21697,N21698,N21699,
  N21700,N21701,N21702,N21703,N21704,N21705,N21706,N21707,N21708,N21709,N21710,N21711,
  N21712,N21713,N21714,N21715,N21716,N21717,N21718,N21719,N21720,N21721,N21722,
  N21723,N21724,N21725,N21726,N21727,N21728,N21729,N21730,N21731,N21732,N21733,
  N21734,N21735,N21736,N21737,N21738,N21739,N21740,N21741,N21742,N21743,N21744,N21745,
  N21746,N21747,N21748,N21749,N21750,N21751,N21752,N21753,N21754,N21755,N21756,
  N21757,N21758,N21759,N21760,N21761,N21762,N21763,N21764,N21765,N21766,N21767,N21768,
  N21769,N21770,N21771,N21772,N21773,N21774,N21775,N21776,N21777,N21778,N21779,
  N21780,N21781,N21782,N21783,N21784,N21785,N21786,N21787,N21788,N21789,N21790,N21791,
  N21792,N21793,N21794,N21795,N21796,N21797,N21798,N21799,N21800,N21801,N21802,
  N21803,N21804,N21805,N21806,N21807,N21808,N21809,N21810,N21811,N21812,N21813,
  N21814,N21815,N21816,N21817,N21818,N21819,N21820,N21821,N21822,N21823,N21824,N21825,
  N21826,N21827,N21828,N21829,N21830,N21831,N21832,N21833,N21834,N21835,N21836,
  N21837,N21838,N21839,N21840,N21841,N21842,N21843,N21844,N21845,N21846,N21847,N21848,
  N21849,N21850,N21851,N21852,N21853,N21854,N21855,N21856,N21857,N21858,N21859,
  N21860,N21861,N21862,N21863,N21864,N21865,N21866,N21867,N21868,N21869,N21870,N21871,
  N21872,N21873,N21874,N21875,N21876,N21877,N21878,N21879,N21880,N21881,N21882,
  N21883,N21884,N21885,N21886,N21887,N21888,N21889,N21890,N21891,N21892,N21893,
  N21894,N21895,N21896,N21897,N21898,N21899,N21900,N21901,N21902,N21903,N21904,N21905,
  N21906,N21907,N21908,N21909,N21910,N21911,N21912,N21913,N21914,N21915,N21916,
  N21917,N21918,N21919,N21920,N21921,N21922,N21923,N21924,N21925,N21926,N21927,N21928,
  N21929,N21930,N21931,N21932,N21933,N21934,N21935,N21936,N21937,N21938,N21939,
  N21940,N21941,N21942,N21943,N21944,N21945,N21946,N21947,N21948,N21949,N21950,N21951,
  N21952,N21953,N21954,N21955,N21956,N21957,N21958,N21959,N21960,N21961,N21962,
  N21963,N21964,N21965,N21966,N21967,N21968,N21969,N21970,N21971,N21972,N21973,
  N21974,N21975,N21976,N21977,N21978,N21979,N21980,N21981,N21982,N21983,N21984,N21985,
  N21986,N21987,N21988,N21989,N21990,N21991,N21992,N21993,N21994,N21995,N21996,
  N21997,N21998,N21999,N22000,N22001,N22002,N22003,N22004,N22005,N22006,N22007,N22008,
  N22009,N22010,N22011,N22012,N22013,N22014,N22015,N22016,N22017,N22018,N22019,
  N22020,N22021,N22022,N22023,N22024,N22025,N22026,N22027,N22028,N22029,N22030,N22031,
  N22032,N22033,N22034,N22035,N22036,N22037,N22038,N22039,N22040,N22041,N22042,
  N22043,N22044,N22045,N22046,N22047,N22048,N22049,N22050,N22051,N22052,N22053,
  N22054,N22055,N22056,N22057,N22058,N22059,N22060,N22061,N22062,N22063,N22064,N22065,
  N22066,N22067,N22068,N22069,N22070,N22071,N22072,N22073,N22074,N22075,N22076,
  N22077,N22078,N22079,N22080,N22081,N22082,N22083,N22084,N22085,N22086,N22087,N22088,
  N22089,N22090,N22091,N22092,N22093,N22094,N22095,N22096,N22097,N22098,N22099,
  N22100,N22101,N22102,N22103,N22104,N22105,N22106,N22107,N22108,N22109,N22110,N22111,
  N22112,N22113,N22114,N22115,N22116,N22117,N22118,N22119,N22120,N22121,N22122,
  N22123,N22124,N22125,N22126,N22127,N22128,N22129,N22130,N22131,N22132,N22133,
  N22134,N22135,N22136,N22137,N22138,N22139,N22140,N22141,N22142,N22143,N22144,N22145,
  N22146,N22147,N22148,N22149,N22150,N22151,N22152,N22153,N22154,N22155,N22156,
  N22157,N22158,N22159,N22160,N22161,N22162,N22163,N22164,N22165,N22166,N22167,N22168,
  N22169,N22170,N22171,N22172,N22173,N22174,N22175,N22176,N22177,N22178,N22179,
  N22180,N22181,N22182,N22183,N22184,N22185,N22186,N22187,N22188,N22189,N22190,N22191,
  N22192,N22193,N22194,N22195,N22196,N22197,N22198,N22199,N22200,N22201,N22202,
  N22203,N22204,N22205,N22206,N22207,N22208,N22209,N22210,N22211,N22212,N22213,
  N22214,N22215,N22216,N22217,N22218,N22219,N22220,N22221,N22222,N22223,N22224,N22225,
  N22226,N22227,N22228,N22229,N22230,N22231,N22232,N22233,N22234,N22235,N22236,
  N22237,N22238,N22239,N22240,N22241,N22242,N22243,N22244,N22245,N22246,N22247,N22248,
  N22249,N22250,N22251,N22252,N22253,N22254,N22255,N22256,N22257,N22258,N22259,
  N22260,N22261,N22262,N22263,N22264,N22265,N22266,N22267,N22268,N22269,N22270,N22271,
  N22272,N22273,N22274,N22275,N22276,N22277,N22278,N22279,N22280,N22281,N22282,
  N22283,N22284,N22285,N22286,N22287,N22288,N22289,N22290,N22291,N22292,N22293,
  N22294,N22295,N22296,N22297,N22298,N22299,N22300,N22301,N22302,N22303,N22304,N22305,
  N22306,N22307,N22308,N22309,N22310,N22311,N22312,N22313,N22314,N22315,N22316,
  N22317,N22318,N22319,N22320,N22321,N22322,N22323,N22324,N22325,N22326,N22327,N22328,
  N22329,N22330,N22331,N22332,N22333,N22334,N22335,N22336,N22337,N22338,N22339,
  N22340,N22341,N22342,N22343,N22344,N22345,N22346,N22347,N22348,N22349,N22350,N22351,
  N22352,N22353,N22354,N22355,N22356,N22357,N22358,N22359,N22360,N22361,N22362,
  N22363,N22364,N22365,N22366,N22367,N22368,N22369,N22370,N22371,N22372,N22373,
  N22374,N22375,N22376,N22377,N22378,N22379,N22380,N22381,N22382,N22383,N22384,N22385,
  N22386,N22387,N22388,N22389,N22390,N22391,N22392,N22393,N22394,N22395,N22396,
  N22397,N22398,N22399,N22400,N22401,N22402,N22403,N22404,N22405,N22406,N22407,N22408,
  N22409,N22410,N22411,N22412,N22413,N22414,N22415,N22416,N22417,N22418,N22419,
  N22420,N22421,N22422,N22423,N22424,N22425,N22426,N22427,N22428,N22429,N22430,N22431,
  N22432,N22433,N22434,N22435,N22436,N22437,N22438,N22439,N22440,N22441,N22442,
  N22443,N22444,N22445,N22446,N22447,N22448,N22449,N22450,N22451,N22452,N22453,
  N22454,N22455,N22456,N22457,N22458,N22459,N22460,N22461,N22462,N22463,N22464,N22465,
  N22466,N22467,N22468,N22469,N22470,N22471,N22472,N22473,N22474,N22475,N22476,
  N22477,N22478,N22479,N22480,N22481,N22482,N22483,N22484,N22485,N22486,N22487,N22488,
  N22489,N22490,N22491,N22492,N22493,N22494,N22495,N22496,N22497,N22498,N22499,
  N22500,N22501,N22502,N22503,N22504,N22505,N22506,N22507,N22508,N22509,N22510,N22511,
  N22512,N22513,N22514,N22515,N22516,N22517,N22518,N22519,N22520,N22521,N22522,
  N22523,N22524,N22525,N22526,N22527,N22528,N22529,N22530,N22531,N22532,N22533,
  N22534,N22535,N22536,N22537,N22538,N22539,N22540,N22541,N22542,N22543,N22544,N22545,
  N22546,N22547,N22548,N22549,N22550,N22551,N22552,N22553,N22554,N22555,N22556,
  N22557,N22558,N22559,N22560,N22561,N22562,N22563,N22564,N22565,N22566,N22567,N22568,
  N22569,N22570,N22571,N22572,N22573,N22574,N22575,N22576,N22577,N22578,N22579,
  N22580,N22581,N22582,N22583,N22584,N22585,N22586,N22587,N22588,N22589,N22590,N22591,
  N22592,N22593,N22594,N22595,N22596,N22597,N22598,N22599,N22600,N22601,N22602,
  N22603,N22604,N22605,N22606,N22607,N22608,N22609,N22610,N22611,N22612,N22613,
  N22614,N22615,N22616,N22617,N22618,N22619,N22620,N22621,N22622,N22623,N22624,N22625,
  N22626,N22627,N22628,N22629,N22630,N22631,N22632,N22633,N22634,N22635,N22636,
  N22637,N22638,N22639,N22640,N22641,N22642,N22643,N22644,N22645,N22646,N22647,N22648,
  N22649,N22650,N22651,N22652,N22653,N22654,N22655,N22656,N22657,N22658,N22659,
  N22660,N22661,N22662,N22663,N22664,N22665,N22666,N22667,N22668,N22669,N22670,N22671,
  N22672,N22673,N22674,N22675,N22676,N22677,N22678,N22679,N22680,N22681,N22682,
  N22683,N22684,N22685,N22686,N22687,N22688,N22689,N22690,N22691,N22692,N22693,
  N22694,N22695,N22696,N22697,N22698,N22699,N22700,N22701,N22702,N22703,N22704,N22705,
  N22706,N22707,N22708,N22709,N22710,N22711,N22712,N22713,N22714,N22715,N22716,
  N22717,N22718,N22719,N22720,N22721,N22722,N22723,N22724,N22725,N22726,N22727,N22728,
  N22729,N22730,N22731,N22732,N22733,N22734,N22735,N22736,N22737,N22738,N22739,
  N22740,N22741,N22742,N22743,N22744,N22745,N22746,N22747,N22748,N22749,N22750,N22751,
  N22752,N22753,N22754,N22755,N22756,N22757,N22758,N22759,N22760,N22761,N22762,
  N22763,N22764,N22765,N22766,N22767,N22768,N22769,N22770,N22771,N22772,N22773,
  N22774,N22775,N22776,N22777,N22778,N22779,N22780,N22781,N22782,N22783,N22784,N22785,
  N22786,N22787,N22788,N22789,N22790,N22791,N22792,N22793,N22794,N22795,N22796,
  N22797,N22798,N22799,N22800,N22801,N22802,N22803,N22804,N22805,N22806,N22807,N22808,
  N22809,N22810,N22811,N22812,N22813,N22814,N22815,N22816,N22817,N22818,N22819,
  N22820,N22821,N22822,N22823,N22824,N22825,N22826,N22827,N22828,N22829,N22830,N22831,
  N22832,N22833,N22834,N22835,N22836,N22837,N22838,N22839,N22840,N22841,N22842,
  N22843,N22844,N22845,N22846,N22847,N22848,N22849,N22850,N22851,N22852,N22853,
  N22854,N22855,N22856,N22857,N22858,N22859,N22860,N22861,N22862,N22863,N22864,N22865,
  N22866,N22867,N22868,N22869,N22870,N22871,N22872,N22873,N22874,N22875,N22876,
  N22877,N22878,N22879,N22880,N22881,N22882,N22883,N22884,N22885,N22886,N22887,N22888,
  N22889,N22890,N22891,N22892,N22893,N22894,N22895,N22896,N22897,N22898,N22899,
  N22900,N22901,N22902,N22903,N22904,N22905,N22906,N22907,N22908,N22909,N22910,N22911,
  N22912,N22913,N22914,N22915,N22916,N22917,N22918,N22919,N22920,N22921,N22922,
  N22923,N22924,N22925,N22926,N22927,N22928,N22929,N22930,N22931,N22932,N22933,
  N22934,N22935,N22936,N22937,N22938,N22939,N22940,N22941,N22942,N22943,N22944,N22945,
  N22946,N22947,N22948,N22949,N22950,N22951,N22952,N22953,N22954,N22955,N22956,
  N22957,N22958,N22959,N22960,N22961,N22962,N22963,N22964,N22965,N22966,N22967,N22968,
  N22969,N22970,N22971,N22972,N22973,N22974,N22975,N22976,N22977,N22978,N22979,
  N22980,N22981,N22982,N22983,N22984,N22985,N22986,N22987,N22988,N22989,N22990,N22991,
  N22992,N22993,N22994,N22995,N22996,N22997,N22998,N22999,N23000,N23001,N23002,
  N23003,N23004,N23005,N23006,N23007,N23008,N23009,N23010,N23011,N23012,N23013,
  N23014,N23015,N23016,N23017,N23018,N23019,N23020,N23021,N23022,N23023,N23024,N23025,
  N23026,N23027,N23028,N23029,N23030,N23031,N23032,N23033,N23034,N23035,N23036,
  N23037,N23038,N23039,N23040,N23041,N23042,N23043,N23044,N23045,N23046,N23047,N23048,
  N23049,N23050,N23051,N23052,N23053,N23054,N23055,N23056,N23057,N23058,N23059,
  N23060,N23061,N23062,N23063,N23064,N23065,N23066,N23067,N23068,N23069,N23070,N23071,
  N23072,N23073,N23074,N23075,N23076,N23077,N23078,N23079,N23080,N23081,N23082,
  N23083,N23084,N23085,N23086,N23087,N23088,N23089,N23090,N23091,N23092,N23093,
  N23094,N23095,N23096,N23097,N23098,N23099,N23100,N23101,N23102,N23103,N23104,N23105,
  N23106,N23107,N23108,N23109,N23110,N23111,N23112,N23113,N23114,N23115,N23116,
  N23117,N23118,N23119,N23120,N23121,N23122,N23123,N23124,N23125,N23126,N23127,N23128,
  N23129,N23130,N23131,N23132,N23133,N23134,N23135,N23136,N23137,N23138,N23139,
  N23140,N23141,N23142,N23143,N23144,N23145,N23146,N23147,N23148,N23149,N23150,N23151,
  N23152,N23153,N23154,N23155,N23156,N23157,N23158,N23159,N23160,N23161,N23162,
  N23163,N23164,N23165,N23166,N23167,N23168,N23169,N23170,N23171,N23172,N23173,
  N23174,N23175,N23176,N23177,N23178,N23179,N23180,N23181,N23182,N23183,N23184,N23185,
  N23186,N23187,N23188,N23189,N23190,N23191,N23192,N23193,N23194,N23195,N23196,
  N23197,N23198,N23199,N23200,N23201,N23202,N23203,N23204,N23205,N23206,N23207,N23208,
  N23209,N23210,N23211,N23212,N23213,N23214,N23215,N23216,N23217,N23218,N23219,
  N23220,N23221,N23222,N23223,N23224,N23225,N23226,N23227,N23228,N23229,N23230,N23231,
  N23232,N23233,N23234,N23235,N23236,N23237,N23238,N23239,N23240,N23241,N23242,
  N23243,N23244,N23245,N23246,N23247,N23248,N23249,N23250,N23251,N23252,N23253,
  N23254,N23255,N23256,N23257,N23258,N23259,N23260,N23261,N23262,N23263,N23264,N23265,
  N23266,N23267,N23268,N23269,N23270,N23271,N23272,N23273,N23274,N23275,N23276,
  N23277,N23278,N23279,N23280,N23281,N23282,N23283,N23284,N23285,N23286,N23287,N23288,
  N23289,N23290,N23291,N23292,N23293,N23294,N23295,N23296,N23297,N23298,N23299,
  N23300,N23301,N23302,N23303,N23304,N23305,N23306,N23307,N23308,N23309,N23310,N23311,
  N23312,N23313,N23314,N23315,N23316,N23317,N23318,N23319,N23320,N23321,N23322,
  N23323,N23324,N23325,N23326,N23327,N23328,N23329,N23330,N23331,N23332,N23333,
  N23334,N23335,N23336,N23337,N23338,N23339,N23340,N23341,N23342,N23343,N23344,N23345,
  N23346,N23347,N23348,N23349,N23350,N23351,N23352,N23353,N23354,N23355,N23356,
  N23357,N23358,N23359,N23360,N23361,N23362,N23363,N23364,N23365,N23366,N23367,N23368,
  N23369,N23370,N23371,N23372,N23373,N23374,N23375,N23376,N23377,N23378,N23379,
  N23380,N23381,N23382,N23383,N23384,N23385,N23386,N23387,N23388,N23389,N23390,N23391,
  N23392,N23393,N23394,N23395,N23396,N23397,N23398,N23399,N23400,N23401,N23402,
  N23403,N23404,N23405,N23406,N23407,N23408,N23409,N23410,N23411,N23412,N23413,
  N23414,N23415,N23416,N23417,N23418,N23419,N23420,N23421,N23422,N23423,N23424,N23425,
  N23426,N23427,N23428,N23429,N23430,N23431,N23432,N23433,N23434,N23435,N23436,
  N23437,N23438,N23439,N23440,N23441,N23442,N23443,N23444,N23445,N23446,N23447,N23448,
  N23449,N23450,N23451,N23452,N23453,N23454,N23455,N23456,N23457,N23458,N23459,
  N23460,N23461,N23462,N23463,N23464,N23465,N23466,N23467,N23468,N23469,N23470,N23471,
  N23472,N23473,N23474,N23475,N23476,N23477,N23478,N23479,N23480,N23481,N23482,
  N23483,N23484,N23485,N23486,N23487,N23488,N23489,N23490,N23491,N23492,N23493,
  N23494,N23495,N23496,N23497,N23498,N23499,N23500,N23501,N23502,N23503,N23504,N23505,
  N23506,N23507,N23508,N23509,N23510,N23511,N23512,N23513,N23514,N23515,N23516,
  N23517,N23518,N23519,N23520,N23521,N23522,N23523,N23524,N23525,N23526,N23527,N23528,
  N23529,N23530,N23531,N23532,N23533,N23534,N23535,N23536,N23537,N23538,N23539,
  N23540,N23541,N23542,N23543,N23544,N23545,N23546,N23547,N23548,N23549,N23550,N23551,
  N23552,N23553,N23554,N23555,N23556,N23557,N23558,N23559,N23560,N23561,N23562,
  N23563,N23564,N23565,N23566,N23567,N23568,N23569,N23570,N23571,N23572,N23573,
  N23574,N23575,N23576,N23577,N23578,N23579,N23580,N23581,N23582,N23583,N23584,N23585,
  N23586,N23587,N23588,N23589,N23590,N23591,N23592,N23593,N23594,N23595,N23596,
  N23597,N23598,N23599,N23600,N23601,N23602,N23603,N23604,N23605,N23606,N23607,N23608,
  N23609,N23610,N23611,N23612,N23613,N23614,N23615,N23616,N23617,N23618,N23619,
  N23620,N23621,N23622,N23623,N23624,N23625,N23626,N23627,N23628,N23629,N23630,N23631,
  N23632,N23633,N23634,N23635,N23636,N23637,N23638,N23639,N23640,N23641,N23642,
  N23643,N23644,N23645,N23646,N23647,N23648,N23649,N23650,N23651,N23652,N23653,
  N23654,N23655,N23656,N23657,N23658,N23659,N23660,N23661,N23662,N23663,N23664,N23665,
  N23666,N23667,N23668,N23669,N23670,N23671,N23672,N23673,N23674,N23675,N23676,
  N23677,N23678,N23679,N23680,N23681,N23682,N23683,N23684,N23685,N23686,N23687,N23688,
  N23689,N23690,N23691,N23692,N23693,N23694,N23695,N23696,N23697,N23698,N23699,
  N23700,N23701,N23702,N23703,N23704,N23705,N23706,N23707,N23708,N23709,N23710,N23711,
  N23712,N23713,N23714,N23715,N23716,N23717,N23718,N23719,N23720,N23721,N23722,
  N23723,N23724,N23725,N23726,N23727,N23728,N23729,N23730,N23731,N23732,N23733,
  N23734,N23735,N23736,N23737,N23738,N23739,N23740,N23741,N23742,N23743,N23744,N23745,
  N23746,N23747,N23748,N23749,N23750,N23751,N23752,N23753,N23754,N23755,N23756,
  N23757,N23758,N23759,N23760,N23761,N23762,N23763,N23764,N23765,N23766,N23767,N23768,
  N23769,N23770,N23771,N23772,N23773,N23774,N23775,N23776,N23777,N23778,N23779,
  N23780,N23781,N23782,N23783,N23784,N23785,N23786,N23787,N23788,N23789,N23790,N23791,
  N23792,N23793,N23794,N23795,N23796,N23797,N23798,N23799,N23800,N23801,N23802,
  N23803,N23804,N23805,N23806,N23807,N23808,N23809,N23810,N23811,N23812,N23813,
  N23814,N23815,N23816,N23817,N23818,N23819,N23820,N23821,N23822,N23823,N23824,N23825,
  N23826,N23827,N23828,N23829,N23830,N23831,N23832,N23833,N23834,N23835,N23836,
  N23837,N23838,N23839,N23840,N23841,N23842,N23843,N23844,N23845,N23846,N23847,N23848,
  N23849,N23850,N23851,N23852,N23853,N23854,N23855,N23856,N23857,N23858,N23859,
  N23860,N23861,N23862,N23863,N23864,N23865,N23866,N23867,N23868,N23869,N23870,N23871,
  N23872,N23873,N23874,N23875,N23876,N23877,N23878,N23879,N23880,N23881,N23882,
  N23883,N23884,N23885,N23886,N23887,N23888,N23889,N23890,N23891,N23892,N23893,
  N23894,N23895,N23896,N23897,N23898,N23899,N23900,N23901,N23902,N23903,N23904,N23905,
  N23906,N23907,N23908,N23909,N23910,N23911,N23912,N23913,N23914,N23915,N23916,
  N23917,N23918,N23919,N23920,N23921,N23922,N23923,N23924,N23925,N23926,N23927,N23928,
  N23929,N23930,N23931,N23932,N23933,N23934,N23935,N23936,N23937,N23938,N23939,
  N23940,N23941,N23942,N23943,N23944,N23945,N23946,N23947,N23948,N23949,N23950,N23951,
  N23952,N23953,N23954,N23955,N23956,N23957,N23958,N23959,N23960,N23961,N23962,
  N23963,N23964,N23965,N23966,N23967,N23968,N23969,N23970,N23971,N23972,N23973,
  N23974,N23975,N23976,N23977,N23978,N23979,N23980,N23981,N23982,N23983,N23984,N23985,
  N23986,N23987,N23988,N23989,N23990,N23991,N23992,N23993,N23994,N23995,N23996,
  N23997,N23998,N23999,N24000,N24001,N24002,N24003,N24004,N24005,N24006,N24007,N24008,
  N24009,N24010,N24011,N24012,N24013,N24014,N24015,N24016,N24017,N24018,N24019,
  N24020,N24021,N24022,N24023,N24024,N24025,N24026,N24027,N24028,N24029,N24030,N24031,
  N24032,N24033,N24034,N24035,N24036,N24037,N24038,N24039,N24040,N24041,N24042,
  N24043,N24044,N24045,N24046,N24047,N24048,N24049,N24050,N24051,N24052,N24053,
  N24054,N24055,N24056,N24057,N24058,N24059,N24060,N24061,N24062,N24063,N24064,N24065,
  N24066,N24067,N24068,N24069,N24070,N24071,N24072,N24073,N24074,N24075,N24076,
  N24077,N24078,N24079,N24080,N24081,N24082,N24083,N24084,N24085,N24086,N24087,N24088,
  N24089,N24090,N24091,N24092,N24093,N24094,N24095,N24096,N24097,N24098,N24099,
  N24100,N24101,N24102,N24103,N24104,N24105,N24106,N24107,N24108,N24109,N24110,N24111,
  N24112,N24113,N24114,N24115,N24116,N24117,N24118,N24119,N24120,N24121,N24122,
  N24123,N24124,N24125,N24126,N24127,N24128,N24129,N24130,N24131,N24132,N24133,
  N24134,N24135,N24136,N24137,N24138,N24139,N24140,N24141,N24142,N24143,N24144,N24145,
  N24146,N24147,N24148,N24149,N24150,N24151,N24152,N24153,N24154,N24155,N24156,
  N24157,N24158,N24159,N24160,N24161,N24162,N24163,N24164,N24165,N24166,N24167,N24168,
  N24169,N24170,N24171,N24172,N24173,N24174,N24175,N24176,N24177,N24178,N24179,
  N24180,N24181,N24182,N24183,N24184,N24185,N24186,N24187,N24188,N24189,N24190,N24191,
  N24192,N24193,N24194,N24195,N24196,N24197,N24198,N24199,N24200,N24201,N24202,
  N24203,N24204,N24205,N24206,N24207,N24208,N24209,N24210,N24211,N24212,N24213,
  N24214,N24215,N24216,N24217,N24218,N24219,N24220,N24221,N24222,N24223,N24224,N24225,
  N24226,N24227,N24228,N24229,N24230,N24231,N24232,N24233,N24234,N24235,N24236,
  N24237,N24238,N24239,N24240,N24241,N24242,N24243,N24244,N24245,N24246,N24247,N24248,
  N24249,N24250,N24251,N24252,N24253,N24254,N24255,N24256,N24257,N24258,N24259,
  N24260,N24261,N24262,N24263,N24264,N24265,N24266,N24267,N24268,N24269,N24270,N24271,
  N24272,N24273,N24274,N24275,N24276,N24277,N24278,N24279,N24280,N24281,N24282,
  N24283,N24284,N24285,N24286,N24287,N24288,N24289,N24290,N24291,N24292,N24293,
  N24294,N24295,N24296,N24297,N24298,N24299,N24300,N24301,N24302,N24303,N24304,N24305,
  N24306,N24307,N24308,N24309,N24310,N24311,N24312,N24313,N24314,N24315,N24316,
  N24317,N24318,N24319,N24320,N24321,N24322,N24323,N24324,N24325,N24326,N24327,N24328,
  N24329,N24330,N24331,N24332,N24333,N24334,N24335,N24336,N24337,N24338,N24339,
  N24340,N24341,N24342,N24343,N24344,N24345,N24346,N24347,N24348,N24349,N24350,N24351,
  N24352,N24353,N24354,N24355,N24356,N24357,N24358,N24359,N24360,N24361,N24362,
  N24363,N24364,N24365,N24366,N24367,N24368,N24369,N24370,N24371,N24372,N24373,
  N24374,N24375,N24376,N24377,N24378,N24379,N24380,N24381,N24382,N24383,N24384,N24385,
  N24386,N24387,N24388,N24389,N24390,N24391,N24392,N24393,N24394,N24395,N24396,
  N24397,N24398,N24399,N24400,N24401,N24402,N24403,N24404,N24405,N24406,N24407,N24408,
  N24409,N24410,N24411,N24412,N24413,N24414,N24415,N24416,N24417,N24418,N24419,
  N24420,N24421,N24422,N24423,N24424,N24425,N24426,N24427,N24428,N24429,N24430,N24431,
  N24432,N24433,N24434,N24435,N24436,N24437,N24438,N24439,N24440,N24441,N24442,
  N24443,N24444,N24445,N24446,N24447,N24448,N24449,N24450,N24451,N24452,N24453,
  N24454,N24455,N24456,N24457,N24458,N24459,N24460,N24461,N24462,N24463,N24464,N24465,
  N24466,N24467,N24468,N24469,N24470,N24471,N24472,N24473,N24474,N24475,N24476,
  N24477,N24478,N24479,N24480,N24481,N24482,N24483,N24484,N24485,N24486,N24487,N24488,
  N24489,N24490,N24491,N24492,N24493,N24494,N24495,N24496,N24497,N24498,N24499,
  N24500,N24501,N24502,N24503,N24504,N24505,N24506,N24507,N24508,N24509,N24510,N24511,
  N24512,N24513,N24514,N24515,N24516,N24517,N24518,N24519,N24520,N24521,N24522,
  N24523,N24524,N24525,N24526,N24527,N24528,N24529,N24530,N24531,N24532,N24533,
  N24534,N24535,N24536,N24537,N24538,N24539,N24540,N24541,N24542,N24543,N24544,N24545,
  N24546,N24547,N24548,N24549,N24550,N24551,N24552,N24553,N24554,N24555,N24556,
  N24557,N24558,N24559,N24560,N24561,N24562,N24563,N24564,N24565,N24566,N24567,N24568,
  N24569,N24570,N24571,N24572,N24573,N24574,N24575,N24576,N24577,N24578,N24579,
  N24580,N24581,N24582,N24583,N24584,N24585,N24586,N24587,N24588,N24589,N24590,N24591,
  N24592,N24593,N24594,N24595,N24596,N24597,N24598,N24599,N24600,N24601,N24602,
  N24603,N24604,N24605,N24606,N24607,N24608,N24609,N24610,N24611,N24612,N24613,
  N24614,N24615,N24616,N24617,N24618,N24619,N24620,N24621,N24622,N24623,N24624,N24625,
  N24626,N24627,N24628,N24629,N24630,N24631,N24632,N24633,N24634,N24635,N24636,
  N24637,N24638,N24639,N24640,N24641,N24642,N24643,N24644,N24645,N24646,N24647,N24648,
  N24649,N24650,N24651,N24652,N24653,N24654,N24655,N24656,N24657,N24658,N24659,
  N24660,N24661,N24662,N24663,N24664,N24665,N24666,N24667,N24668,N24669,N24670,N24671,
  N24672,N24673,N24674,N24675,N24676,N24677,N24678,N24679,N24680,N24681,N24682,
  N24683,N24684,N24685,N24686,N24687,N24688,N24689,N24690,N24691,N24692,N24693,
  N24694,N24695,N24696,N24697,N24698,N24699,N24700,N24701,N24702,N24703,N24704,N24705,
  N24706,N24707,N24708,N24709,N24710,N24711,N24712,N24713,N24714,N24715,N24716,
  N24717,N24718,N24719,N24720,N24721,N24722,N24723,N24724,N24725,N24726,N24727,N24728,
  N24729,N24730,N24731,N24732,N24733,N24734,N24735,N24736,N24737,N24738,N24739,
  N24740,N24741,N24742,N24743,N24744,N24745,N24746,N24747,N24748,N24749,N24750,N24751,
  N24752,N24753,N24754,N24755,N24756,N24757,N24758,N24759,N24760,N24761,N24762,
  N24763,N24764,N24765,N24766,N24767,N24768,N24769,N24770,N24771,N24772,N24773,
  N24774,N24775,N24776,N24777,N24778,N24779,N24780,N24781,N24782,N24783,N24784,N24785,
  N24786,N24787,N24788,N24789,N24790,N24791,N24792,N24793,N24794,N24795,N24796,
  N24797,N24798,N24799,N24800,N24801,N24802,N24803,N24804,N24805,N24806,N24807,N24808,
  N24809,N24810,N24811,N24812,N24813,N24814,N24815,N24816,N24817,N24818,N24819,
  N24820,N24821,N24822,N24823,N24824,N24825,N24826,N24827,N24828,N24829,N24830,N24831,
  N24832,N24833,N24834,N24835,N24836,N24837,N24838,N24839,N24840,N24841,N24842,
  N24843,N24844,N24845,N24846,N24847,N24848,N24849,N24850,N24851,N24852,N24853,
  N24854,N24855,N24856,N24857,N24858,N24859,N24860,N24861,N24862,N24863,N24864,N24865,
  N24866,N24867,N24868,N24869,N24870,N24871,N24872,N24873,N24874,N24875,N24876,
  N24877,N24878,N24879,N24880,N24881,N24882,N24883,N24884,N24885,N24886,N24887,N24888,
  N24889,N24890,N24891,N24892,N24893,N24894,N24895,N24896,N24897,N24898,N24899,
  N24900,N24901,N24902,N24903,N24904,N24905,N24906,N24907,N24908,N24909,N24910,N24911,
  N24912,N24913,N24914,N24915,N24916,N24917,N24918,N24919,N24920,N24921,N24922,
  N24923,N24924,N24925,N24926,N24927,N24928,N24929,N24930,N24931,N24932,N24933,
  N24934,N24935,N24936,N24937,N24938,N24939,N24940,N24941,N24942,N24943,N24944,N24945,
  N24946,N24947,N24948,N24949,N24950,N24951,N24952,N24953,N24954,N24955,N24956,
  N24957,N24958,N24959,N24960,N24961,N24962,N24963,N24964,N24965,N24966,N24967,N24968,
  N24969,N24970,N24971,N24972,N24973,N24974,N24975,N24976,N24977,N24978,N24979,
  N24980,N24981,N24982,N24983,N24984,N24985,N24986,N24987,N24988,N24989,N24990,N24991,
  N24992,N24993,N24994,N24995,N24996,N24997,N24998,N24999,N25000,N25001,N25002,
  N25003,N25004,N25005,N25006,N25007,N25008,N25009,N25010,N25011,N25012,N25013,
  N25014,N25015,N25016,N25017,N25018,N25019,N25020,N25021,N25022,N25023,N25024,N25025,
  N25026,N25027,N25028,N25029,N25030,N25031,N25032,N25033,N25034,N25035,N25036,
  N25037,N25038,N25039,N25040,N25041,N25042,N25043,N25044,N25045,N25046,N25047,N25048,
  N25049,N25050,N25051,N25052,N25053,N25054,N25055,N25056,N25057,N25058,N25059,
  N25060,N25061,N25062,N25063,N25064,N25065,N25066,N25067,N25068,N25069,N25070,N25071,
  N25072,N25073,N25074,N25075,N25076,N25077,N25078,N25079,N25080,N25081,N25082,
  N25083,N25084,N25085,N25086,N25087,N25088,N25089,N25090,N25091,N25092,N25093,
  N25094,N25095,N25096,N25097,N25098,N25099,N25100,N25101,N25102,N25103,N25104,N25105,
  N25106,N25107,N25108,N25109,N25110,N25111,N25112,N25113,N25114,N25115,N25116,
  N25117,N25118,N25119,N25120,N25121,N25122,N25123,N25124,N25125,N25126,N25127,N25128,
  N25129,N25130,N25131,N25132,N25133,N25134,N25135,N25136,N25137,N25138,N25139,
  N25140,N25141,N25142,N25143,N25144,N25145,N25146,N25147,N25148,N25149,N25150,N25151,
  N25152,N25153,N25154,N25155,N25156,N25157,N25158,N25159,N25160,N25161,N25162,
  N25163,N25164,N25165,N25166,N25167,N25168,N25169,N25170,N25171,N25172,N25173,
  N25174,N25175,N25176,N25177,N25178,N25179,N25180,N25181,N25182,N25183,N25184,N25185,
  N25186,N25187,N25188,N25189,N25190,N25191,N25192,N25193,N25194,N25195,N25196,
  N25197,N25198,N25199,N25200,N25201,N25202,N25203,N25204,N25205,N25206,N25207,N25208,
  N25209,N25210,N25211,N25212,N25213,N25214,N25215,N25216,N25217,N25218,N25219,
  N25220,N25221,N25222,N25223,N25224,N25225,N25226,N25227,N25228,N25229,N25230,N25231,
  N25232,N25233,N25234,N25235,N25236,N25237,N25238,N25239,N25240,N25241,N25242,
  N25243,N25244,N25245,N25246,N25247,N25248,N25249,N25250,N25251,N25252,N25253,
  N25254,N25255,N25256,N25257,N25258,N25259,N25260,N25261,N25262,N25263,N25264,N25265,
  N25266,N25267,N25268,N25269,N25270,N25271,N25272,N25273,N25274,N25275,N25276,
  N25277,N25278,N25279,N25280,N25281,N25282,N25283,N25284,N25285,N25286,N25287,N25288,
  N25289,N25290,N25291,N25292,N25293,N25294,N25295,N25296,N25297,N25298,N25299,
  N25300,N25301,N25302,N25303,N25304,N25305,N25306,N25307,N25308,N25309,N25310,N25311,
  N25312,N25313,N25314,N25315,N25316,N25317,N25318,N25319,N25320,N25321,N25322,
  N25323,N25324,N25325,N25326,N25327,N25328,N25329,N25330,N25331,N25332,N25333,
  N25334,N25335,N25336,N25337,N25338,N25339,N25340,N25341,N25342,N25343,N25344,N25345,
  N25346,N25347,N25348,N25349,N25350,N25351,N25352,N25353,N25354,N25355,N25356,
  N25357,N25358,N25359,N25360,N25361,N25362,N25363,N25364,N25365,N25366,N25367,N25368,
  N25369,N25370,N25371,N25372,N25373,N25374,N25375,N25376,N25377,N25378,N25379,
  N25380,N25381,N25382,N25383,N25384,N25385,N25386,N25387,N25388,N25389,N25390,N25391,
  N25392,N25393,N25394,N25395,N25396,N25397,N25398,N25399,N25400,N25401,N25402,
  N25403,N25404,N25405,N25406,N25407,N25408,N25409,N25410,N25411,N25412,N25413,
  N25414,N25415,N25416,N25417,N25418,N25419,N25420,N25421,N25422,N25423,N25424,N25425,
  N25426,N25427,N25428,N25429,N25430,N25431,N25432,N25433,N25434,N25435,N25436,
  N25437,N25438,N25439,N25440,N25441,N25442,N25443,N25444,N25445,N25446,N25447,N25448,
  N25449,N25450,N25451,N25452,N25453,N25454,N25455,N25456,N25457,N25458,N25459,
  N25460,N25461,N25462,N25463,N25464,N25465,N25466,N25467,N25468,N25469,N25470,N25471,
  N25472,N25473,N25474,N25475,N25476,N25477,N25478,N25479,N25480,N25481,N25482,
  N25483,N25484,N25485,N25486,N25487,N25488,N25489,N25490,N25491,N25492,N25493,
  N25494,N25495,N25496,N25497,N25498,N25499,N25500,N25501,N25502,N25503,N25504,N25505,
  N25506,N25507,N25508,N25509,N25510,N25511,N25512,N25513,N25514,N25515,N25516,
  N25517,N25518,N25519,N25520,N25521,N25522,N25523,N25524,N25525,N25526,N25527,N25528,
  N25529,N25530,N25531,N25532,N25533,N25534,N25535,N25536,N25537,N25538,N25539,
  N25540,N25541,N25542,N25543,N25544,N25545,N25546,N25547,N25548,N25549,N25550,N25551,
  N25552,N25553,N25554,N25555,N25556,N25557,N25558,N25559,N25560,N25561,N25562,
  N25563,N25564,N25565,N25566,N25567,N25568,N25569,N25570,N25571,N25572,N25573,
  N25574,N25575,N25576,N25577,N25578,N25579,N25580,N25581,N25582,N25583,N25584,N25585,
  N25586,N25587,N25588,N25589,N25590,N25591,N25592,N25593,N25594,N25595,N25596,
  N25597,N25598,N25599,N25600,N25601,N25602,N25603,N25604,N25605,N25606,N25607,N25608,
  N25609,N25610,N25611,N25612,N25613,N25614,N25615,N25616,N25617,N25618,N25619,
  N25620,N25621,N25622,N25623,N25624,N25625,N25626,N25627,N25628,N25629,N25630,N25631,
  N25632,N25633,N25634,N25635,N25636,N25637,N25638,N25639,N25640,N25641,N25642,
  N25643,N25644,N25645,N25646,N25647,N25648,N25649,N25650,N25651,N25652,N25653,
  N25654,N25655,N25656,N25657,N25658,N25659,N25660,N25661,N25662,N25663,N25664,N25665,
  N25666,N25667,N25668,N25669,N25670,N25671,N25672,N25673,N25674,N25675,N25676,
  N25677,N25678,N25679,N25680,N25681,N25682,N25683,N25684,N25685,N25686,N25687,N25688,
  N25689,N25690,N25691,N25692,N25693,N25694,N25695,N25696,N25697,N25698,N25699,
  N25700,N25701,N25702,N25703,N25704,N25705,N25706,N25707,N25708,N25709,N25710,N25711,
  N25712,N25713,N25714,N25715,N25716,N25717,N25718,N25719,N25720,N25721,N25722,
  N25723,N25724,N25725,N25726,N25727,N25728,N25729,N25730,N25731,N25732,N25733,
  N25734,N25735,N25736,N25737,N25738,N25739,N25740,N25741,N25742,N25743,N25744,N25745,
  N25746,N25747,N25748,N25749,N25750,N25751,N25752,N25753,N25754,N25755,N25756,
  N25757,N25758,N25759,N25760,N25761,N25762,N25763,N25764,N25765,N25766,N25767,N25768,
  N25769,N25770,N25771,N25772,N25773,N25774,N25775,N25776,N25777,N25778,N25779,
  N25780,N25781,N25782,N25783,N25784,N25785,N25786,N25787,N25788,N25789,N25790,N25791,
  N25792,N25793,N25794,N25795,N25796,N25797,N25798,N25799,N25800,N25801,N25802,
  N25803,N25804,N25805,N25806,N25807,N25808,N25809,N25810,N25811,N25812,N25813,
  N25814,N25815,N25816,N25817,N25818,N25819,N25820,N25821,N25822,N25823,N25824,N25825,
  N25826,N25827,N25828,N25829,N25830,N25831,N25832,N25833,N25834,N25835,N25836,
  N25837,N25838,N25839,N25840,N25841,N25842,N25843,N25844,N25845,N25846,N25847,N25848,
  N25849,N25850,N25851,N25852,N25853,N25854,N25855,N25856,N25857,N25858,N25859,
  N25860,N25861,N25862,N25863,N25864,N25865,N25866,N25867,N25868,N25869,N25870,N25871,
  N25872,N25873,N25874,N25875,N25876,N25877,N25878,N25879,N25880,N25881,N25882,
  N25883,N25884,N25885,N25886,N25887,N25888,N25889,N25890,N25891,N25892,N25893,
  N25894,N25895,N25896,N25897,N25898,N25899,N25900,N25901,N25902,N25903,N25904,N25905,
  N25906,N25907,N25908,N25909,N25910,N25911,N25912,N25913,N25914,N25915,N25916,
  N25917,N25918,N25919,N25920,N25921,N25922,N25923,N25924,N25925,N25926,N25927,N25928,
  N25929,N25930,N25931,N25932,N25933,N25934,N25935,N25936,N25937,N25938,N25939,
  N25940,N25941,N25942,N25943,N25944,N25945,N25946,N25947,N25948,N25949,N25950,N25951,
  N25952,N25953,N25954,N25955,N25956,N25957,N25958,N25959,N25960,N25961,N25962,
  N25963,N25964,N25965,N25966,N25967,N25968,N25969,N25970,N25971,N25972,N25973,
  N25974,N25975,N25976,N25977,N25978,N25979,N25980,N25981,N25982,N25983,N25984,N25985,
  N25986,N25987,N25988,N25989,N25990,N25991,N25992,N25993,N25994,N25995,N25996,
  N25997,N25998,N25999,N26000,N26001,N26002,N26003,N26004,N26005,N26006,N26007,N26008,
  N26009,N26010,N26011,N26012,N26013,N26014,N26015,N26016,N26017,N26018,N26019,
  N26020,N26021,N26022,N26023,N26024,N26025,N26026,N26027,N26028,N26029,N26030,N26031,
  N26032,N26033,N26034,N26035,N26036,N26037,N26038,N26039,N26040,N26041,N26042,
  N26043,N26044,N26045,N26046,N26047,N26048,N26049,N26050,N26051,N26052,N26053,
  N26054,N26055,N26056,N26057,N26058,N26059,N26060,N26061,N26062,N26063,N26064,N26065,
  N26066,N26067,N26068,N26069,N26070,N26071,N26072,N26073,N26074,N26075,N26076,
  N26077,N26078,N26079,N26080,N26081,N26082,N26083,N26084,N26085,N26086,N26087,N26088,
  N26089,N26090,N26091,N26092,N26093,N26094,N26095,N26096,N26097,N26098,N26099,
  N26100,N26101,N26102,N26103,N26104,N26105,N26106,N26107,N26108,N26109,N26110,N26111,
  N26112,N26113,N26114,N26115,N26116,N26117,N26118,N26119,N26120,N26121,N26122,
  N26123,N26124,N26125,N26126,N26127,N26128,N26129,N26130,N26131,N26132,N26133,
  N26134,N26135,N26136,N26137,N26138,N26139,N26140,N26141,N26142,N26143,N26144,N26145,
  N26146,N26147,N26148,N26149,N26150,N26151,N26152,N26153,N26154,N26155,N26156,
  N26157,N26158,N26159,N26160,N26161,N26162,N26163,N26164,N26165,N26166,N26167,N26168,
  N26169,N26170,N26171,N26172,N26173,N26174,N26175,N26176,N26177,N26178,N26179,
  N26180,N26181,N26182,N26183,N26184,N26185,N26186,N26187,N26188,N26189,N26190,N26191,
  N26192,N26193,N26194,N26195,N26196,N26197,N26198,N26199,N26200,N26201,N26202,
  N26203,N26204,N26205,N26206,N26207,N26208,N26209,N26210,N26211,N26212,N26213,
  N26214,N26215,N26216,N26217,N26218,N26219,N26220,N26221,N26222,N26223,N26224,N26225,
  N26226,N26227,N26228,N26229,N26230,N26231,N26232,N26233,N26234,N26235,N26236,
  N26237,N26238,N26239,N26240,N26241,N26242,N26243,N26244,N26245,N26246,N26247,N26248,
  N26249,N26250,N26251,N26252,N26253,N26254,N26255,N26256,N26257,N26258,N26259,
  N26260,N26261,N26262,N26263,N26264,N26265,N26266,N26267,N26268,N26269,N26270,N26271,
  N26272,N26273,N26274,N26275,N26276,N26277,N26278,N26279,N26280,N26281,N26282,
  N26283,N26284,N26285,N26286,N26287,N26288,N26289,N26290,N26291,N26292,N26293,
  N26294,N26295,N26296,N26297,N26298,N26299,N26300,N26301,N26302,N26303,N26304,N26305,
  N26306,N26307,N26308,N26309,N26310,N26311,N26312,N26313,N26314,N26315,N26316,
  N26317,N26318,N26319,N26320,N26321,N26322,N26323,N26324,N26325,N26326,N26327,N26328,
  N26329,N26330,N26331,N26332,N26333,N26334,N26335,N26336,N26337,N26338,N26339,
  N26340,N26341,N26342,N26343,N26344,N26345,N26346,N26347,N26348,N26349,N26350,N26351,
  N26352,N26353,N26354,N26355,N26356,N26357,N26358,N26359,N26360,N26361,N26362,
  N26363,N26364,N26365,N26366,N26367,N26368,N26369,N26370,N26371,N26372,N26373,
  N26374,N26375,N26376,N26377,N26378,N26379,N26380,N26381,N26382,N26383,N26384,N26385,
  N26386,N26387,N26388,N26389,N26390,N26391,N26392,N26393,N26394,N26395,N26396,
  N26397,N26398,N26399,N26400,N26401,N26402,N26403,N26404,N26405,N26406,N26407,N26408,
  N26409,N26410,N26411,N26412,N26413,N26414,N26415,N26416,N26417,N26418,N26419,
  N26420,N26421,N26422,N26423,N26424,N26425,N26426,N26427,N26428,N26429,N26430,N26431,
  N26432,N26433,N26434,N26435,N26436,N26437,N26438,N26439,N26440,N26441,N26442,
  N26443,N26444,N26445,N26446,N26447,N26448,N26449,N26450,N26451,N26452,N26453,
  N26454,N26455,N26456,N26457,N26458,N26459,N26460,N26461,N26462,N26463,N26464,N26465,
  N26466,N26467,N26468,N26469,N26470,N26471,N26472,N26473,N26474,N26475,N26476,
  N26477,N26478,N26479,N26480,N26481,N26482,N26483,N26484,N26485,N26486,N26487,N26488,
  N26489,N26490,N26491,N26492,N26493,N26494,N26495,N26496,N26497,N26498,N26499,
  N26500,N26501,N26502,N26503,N26504,N26505,N26506,N26507,N26508,N26509,N26510,N26511,
  N26512,N26513,N26514,N26515,N26516,N26517,N26518,N26519,N26520,N26521,N26522,
  N26523,N26524,N26525,N26526,N26527,N26528,N26529,N26530,N26531,N26532,N26533,
  N26534,N26535,N26536,N26537,N26538,N26539,N26540,N26541,N26542,N26543,N26544,N26545,
  N26546,N26547,N26548,N26549,N26550,N26551,N26552,N26553,N26554,N26555,N26556,
  N26557,N26558,N26559,N26560,N26561,N26562,N26563,N26564,N26565,N26566,N26567,N26568,
  N26569,N26570,N26571,N26572,N26573,N26574,N26575,N26576,N26577,N26578,N26579,
  N26580,N26581,N26582,N26583,N26584,N26585,N26586,N26587,N26588,N26589,N26590,N26591,
  N26592,N26593,N26594,N26595,N26596,N26597,N26598,N26599,N26600,N26601,N26602,
  N26603,N26604,N26605,N26606,N26607,N26608,N26609,N26610,N26611,N26612,N26613,
  N26614,N26615,N26616,N26617,N26618,N26619,N26620,N26621,N26622,N26623,N26624,N26625,
  N26626,N26627,N26628,N26629,N26630,N26631,N26632,N26633,N26634,N26635,N26636,
  N26637,N26638,N26639,N26640,N26641,N26642,N26643,N26644,N26645,N26646,N26647,N26648,
  N26649,N26650,N26651,N26652,N26653,N26654,N26655,N26656,N26657,N26658,N26659,
  N26660,N26661,N26662,N26663,N26664,N26665,N26666,N26667,N26668,N26669,N26670,N26671,
  N26672,N26673,N26674,N26675,N26676,N26677,N26678,N26679,N26680,N26681,N26682,
  N26683,N26684,N26685,N26686,N26687,N26688,N26689,N26690,N26691,N26692,N26693,
  N26694,N26695,N26696,N26697,N26698,N26699,N26700,N26701,N26702,N26703,N26704,N26705,
  N26706,N26707,N26708,N26709,N26710,N26711,N26712,N26713,N26714,N26715,N26716,
  N26717,N26718,N26719,N26720,N26721,N26722,N26723,N26724,N26725,N26726,N26727,N26728,
  N26729,N26730,N26731,N26732,N26733,N26734,N26735,N26736,N26737,N26738,N26739,
  N26740,N26741,N26742,N26743,N26744,N26745,N26746,N26747,N26748,N26749,N26750,N26751,
  N26752,N26753,N26754,N26755,N26756,N26757,N26758,N26759,N26760,N26761,N26762,
  N26763,N26764,N26765,N26766,N26767,N26768,N26769,N26770,N26771,N26772,N26773,
  N26774,N26775,N26776,N26777,N26778,N26779,N26780,N26781,N26782,N26783,N26784,N26785,
  N26786,N26787,N26788,N26789,N26790,N26791,N26792,N26793,N26794,N26795,N26796,
  N26797,N26798,N26799,N26800,N26801,N26802,N26803,N26804,N26805,N26806,N26807,N26808,
  N26809,N26810,N26811,N26812,N26813,N26814,N26815,N26816,N26817,N26818,N26819,
  N26820,N26821,N26822,N26823,N26824,N26825,N26826,N26827,N26828,N26829,N26830,N26831,
  N26832,N26833,N26834,N26835,N26836,N26837,N26838,N26839,N26840,N26841,N26842,
  N26843,N26844,N26845,N26846,N26847,N26848,N26849,N26850,N26851,N26852,N26853,
  N26854,N26855,N26856,N26857,N26858,N26859,N26860,N26861,N26862,N26863,N26864,N26865,
  N26866,N26867,N26868,N26869,N26870,N26871,N26872,N26873,N26874,N26875,N26876,
  N26877,N26878,N26879,N26880,N26881,N26882,N26883,N26884,N26885,N26886,N26887,N26888,
  N26889,N26890,N26891,N26892,N26893,N26894,N26895,N26896,N26897,N26898,N26899,
  N26900,N26901,N26902,N26903,N26904,N26905,N26906,N26907,N26908,N26909,N26910,N26911,
  N26912,N26913,N26914,N26915,N26916,N26917,N26918,N26919,N26920,N26921,N26922,
  N26923,N26924,N26925,N26926,N26927,N26928,N26929,N26930,N26931,N26932,N26933,
  N26934,N26935,N26936,N26937,N26938,N26939,N26940,N26941,N26942,N26943,N26944,N26945,
  N26946,N26947,N26948,N26949,N26950,N26951,N26952,N26953,N26954,N26955,N26956,
  N26957,N26958,N26959,N26960,N26961,N26962,N26963,N26964,N26965,N26966,N26967,N26968,
  N26969,N26970,N26971,N26972,N26973,N26974,N26975,N26976,N26977,N26978,N26979,
  N26980,N26981,N26982,N26983,N26984,N26985,N26986,N26987,N26988,N26989,N26990,N26991,
  N26992,N26993,N26994,N26995,N26996,N26997,N26998,N26999,N27000,N27001,N27002,
  N27003,N27004,N27005,N27006,N27007,N27008,N27009,N27010,N27011,N27012,N27013,
  N27014,N27015,N27016,N27017,N27018,N27019,N27020,N27021,N27022,N27023,N27024,N27025,
  N27026,N27027,N27028,N27029,N27030,N27031,N27032,N27033,N27034,N27035,N27036,
  N27037,N27038,N27039,N27040,N27041,N27042,N27043,N27044,N27045,N27046,N27047,N27048,
  N27049,N27050,N27051,N27052,N27053,N27054,N27055,N27056,N27057,N27058,N27059,
  N27060,N27061,N27062,N27063,N27064,N27065,N27066,N27067,N27068,N27069,N27070,N27071,
  N27072,N27073,N27074,N27075,N27076,N27077,N27078,N27079,N27080,N27081,N27082,
  N27083,N27084,N27085,N27086,N27087,N27088,N27089,N27090,N27091,N27092,N27093,
  N27094,N27095,N27096,N27097,N27098,N27099,N27100,N27101,N27102,N27103,N27104,N27105,
  N27106,N27107,N27108,N27109,N27110,N27111,N27112,N27113,N27114,N27115,N27116,
  N27117,N27118,N27119,N27120,N27121,N27122,N27123,N27124,N27125,N27126,N27127,N27128,
  N27129,N27130,N27131,N27132,N27133,N27134,N27135,N27136,N27137,N27138,N27139,
  N27140,N27141,N27142,N27143,N27144,N27145,N27146,N27147,N27148,N27149,N27150,N27151,
  N27152,N27153,N27154,N27155,N27156,N27157,N27158,N27159,N27160,N27161,N27162,
  N27163,N27164,N27165,N27166,N27167,N27168,N27169,N27170,N27171,N27172,N27173,
  N27174,N27175,N27176,N27177,N27178,N27179,N27180,N27181,N27182,N27183,N27184,N27185,
  N27186,N27187,N27188,N27189,N27190,N27191,N27192,N27193,N27194,N27195,N27196,
  N27197,N27198,N27199,N27200,N27201,N27202,N27203,N27204,N27205,N27206,N27207,N27208,
  N27209,N27210,N27211,N27212,N27213,N27214,N27215,N27216,N27217,N27218,N27219,
  N27220,N27221,N27222,N27223,N27224,N27225,N27226,N27227,N27228,N27229,N27230,N27231,
  N27232,N27233,N27234,N27235,N27236,N27237,N27238,N27239,N27240,N27241,N27242,
  N27243,N27244,N27245,N27246,N27247,N27248,N27249,N27250,N27251,N27252,N27253,
  N27254,N27255,N27256,N27257,N27258,N27259,N27260,N27261,N27262,N27263,N27264,N27265,
  N27266,N27267,N27268,N27269,N27270,N27271,N27272,N27273,N27274,N27275,N27276,
  N27277,N27278,N27279,N27280,N27281,N27282,N27283,N27284,N27285,N27286,N27287,N27288,
  N27289,N27290,N27291,N27292,N27293,N27294,N27295,N27296,N27297,N27298,N27299,
  N27300,N27301,N27302,N27303,N27304,N27305,N27306,N27307,N27308,N27309,N27310,N27311,
  N27312,N27313,N27314,N27315,N27316,N27317,N27318,N27319,N27320,N27321,N27322,
  N27323,N27324,N27325,N27326,N27327,N27328,N27329,N27330,N27331,N27332,N27333,
  N27334,N27335,N27336,N27337,N27338,N27339,N27340,N27341,N27342,N27343,N27344,N27345,
  N27346,N27347,N27348,N27349,N27350,N27351,N27352,N27353,N27354,N27355,N27356,
  N27357,N27358,N27359,N27360,N27361,N27362,N27363,N27364,N27365,N27366,N27367,N27368,
  N27369,N27370,N27371,N27372,N27373,N27374,N27375,N27376,N27377,N27378,N27379,
  N27380,N27381,N27382,N27383,N27384,N27385,N27386,N27387,N27388,N27389,N27390,N27391,
  N27392,N27393,N27394,N27395,N27396,N27397,N27398,N27399,N27400,N27401,N27402,
  N27403,N27404,N27405,N27406,N27407,N27408,N27409,N27410,N27411,N27412,N27413,
  N27414,N27415,N27416,N27417,N27418,N27419,N27420,N27421,N27422,N27423,N27424,N27425,
  N27426,N27427,N27428,N27429,N27430,N27431,N27432,N27433,N27434,N27435,N27436,
  N27437,N27438,N27439,N27440,N27441,N27442,N27443,N27444,N27445,N27446,N27447,N27448,
  N27449,N27450,N27451,N27452,N27453,N27454,N27455,N27456,N27457,N27458,N27459,
  N27460,N27461,N27462,N27463,N27464,N27465,N27466,N27467,N27468,N27469,N27470,N27471,
  N27472,N27473,N27474,N27475,N27476,N27477,N27478,N27479,N27480,N27481,N27482,
  N27483,N27484,N27485,N27486,N27487,N27488,N27489,N27490,N27491,N27492,N27493,
  N27494,N27495,N27496,N27497,N27498,N27499,N27500,N27501,N27502,N27503,N27504,N27505,
  N27506,N27507,N27508,N27509,N27510,N27511,N27512,N27513,N27514,N27515,N27516,
  N27517,N27518,N27519,N27520,N27521,N27522,N27523,N27524,N27525,N27526,N27527,N27528,
  N27529,N27530,N27531,N27532,N27533,N27534,N27535,N27536,N27537,N27538,N27539,
  N27540,N27541,N27542,N27543,N27544,N27545,N27546,N27547,N27548,N27549,N27550,N27551,
  N27552,N27553,N27554,N27555,N27556,N27557,N27558,N27559,N27560,N27561,N27562,
  N27563,N27564,N27565,N27566,N27567,N27568,N27569,N27570,N27571,N27572,N27573,
  N27574,N27575,N27576,N27577,N27578,N27579,N27580,N27581,N27582,N27583,N27584,N27585,
  N27586,N27587,N27588,N27589,N27590,N27591,N27592,N27593,N27594,N27595,N27596,
  N27597,N27598,N27599,N27600,N27601,N27602,N27603,N27604,N27605,N27606,N27607,N27608,
  N27609,N27610,N27611,N27612,N27613,N27614,N27615,N27616,N27617,N27618,N27619,
  N27620,N27621,N27622,N27623,N27624,N27625,N27626,N27627,N27628,N27629,N27630,N27631,
  N27632,N27633,N27634,N27635,N27636,N27637,N27638,N27639,N27640,N27641,N27642,
  N27643,N27644,N27645,N27646,N27647,N27648,N27649,N27650,N27651,N27652,N27653,
  N27654,N27655,N27656,N27657,N27658,N27659,N27660,N27661,N27662,N27663,N27664,N27665,
  N27666,N27667,N27668,N27669,N27670,N27671,N27672,N27673,N27674,N27675,N27676,
  N27677,N27678,N27679,N27680,N27681,N27682,N27683,N27684,N27685,N27686,N27687,N27688,
  N27689,N27690,N27691,N27692,N27693,N27694,N27695,N27696,N27697,N27698,N27699,
  N27700,N27701,N27702,N27703,N27704,N27705,N27706,N27707,N27708,N27709,N27710,N27711,
  N27712,N27713,N27714,N27715,N27716,N27717,N27718,N27719,N27720,N27721,N27722,
  N27723,N27724,N27725,N27726,N27727,N27728,N27729,N27730,N27731,N27732,N27733,
  N27734,N27735,N27736,N27737,N27738,N27739,N27740,N27741,N27742,N27743,N27744,N27745,
  N27746,N27747,N27748,N27749,N27750,N27751,N27752,N27753,N27754,N27755,N27756,
  N27757,N27758,N27759,N27760,N27761,N27762,N27763,N27764,N27765,N27766,N27767,N27768,
  N27769,N27770,N27771,N27772,N27773,N27774,N27775,N27776,N27777,N27778,N27779,
  N27780,N27781,N27782,N27783,N27784,N27785,N27786,N27787,N27788,N27789,N27790,N27791,
  N27792,N27793,N27794,N27795,N27796,N27797,N27798,N27799,N27800,N27801,N27802,
  N27803,N27804,N27805,N27806,N27807,N27808,N27809,N27810,N27811,N27812,N27813,
  N27814,N27815,N27816,N27817,N27818,N27819,N27820,N27821,N27822,N27823,N27824,N27825,
  N27826,N27827,N27828,N27829,N27830,N27831,N27832,N27833,N27834,N27835,N27836,
  N27837,N27838,N27839,N27840,N27841,N27842,N27843,N27844,N27845,N27846,N27847,N27848,
  N27849,N27850,N27851,N27852,N27853,N27854,N27855,N27856,N27857,N27858,N27859,
  N27860,N27861,N27862,N27863,N27864,N27865,N27866,N27867,N27868,N27869,N27870,N27871,
  N27872,N27873,N27874,N27875,N27876,N27877,N27878,N27879,N27880,N27881,N27882,
  N27883,N27884,N27885,N27886,N27887,N27888,N27889,N27890,N27891,N27892,N27893,
  N27894,N27895,N27896,N27897,N27898,N27899,N27900,N27901,N27902,N27903,N27904,N27905,
  N27906,N27907,N27908,N27909,N27910,N27911,N27912,N27913,N27914,N27915,N27916,
  N27917,N27918,N27919,N27920,N27921,N27922,N27923,N27924,N27925,N27926,N27927,N27928,
  N27929,N27930,N27931,N27932,N27933,N27934,N27935,N27936,N27937,N27938,N27939,
  N27940,N27941,N27942,N27943,N27944,N27945,N27946,N27947,N27948,N27949,N27950,N27951,
  N27952,N27953,N27954,N27955,N27956,N27957,N27958,N27959,N27960,N27961,N27962,
  N27963,N27964,N27965,N27966,N27967,N27968,N27969,N27970,N27971,N27972,N27973,
  N27974,N27975,N27976,N27977,N27978,N27979,N27980,N27981,N27982,N27983,N27984,N27985,
  N27986,N27987,N27988,N27989,N27990,N27991,N27992,N27993,N27994,N27995,N27996,
  N27997,N27998,N27999,N28000,N28001,N28002,N28003,N28004,N28005,N28006,N28007,N28008,
  N28009,N28010,N28011,N28012,N28013,N28014,N28015,N28016,N28017,N28018,N28019,
  N28020,N28021,N28022,N28023,N28024,N28025,N28026,N28027,N28028,N28029,N28030,N28031,
  N28032,N28033,N28034,N28035,N28036,N28037,N28038,N28039,N28040,N28041,N28042,
  N28043,N28044,N28045,N28046,N28047,N28048,N28049,N28050,N28051,N28052,N28053,
  N28054,N28055,N28056,N28057,N28058,N28059,N28060,N28061,N28062,N28063,N28064,N28065,
  N28066,N28067,N28068,N28069,N28070,N28071,N28072,N28073,N28074,N28075,N28076,
  N28077,N28078,N28079,N28080,N28081,N28082,N28083,N28084,N28085,N28086,N28087,N28088,
  N28089,N28090,N28091,N28092,N28093,N28094,N28095,N28096,N28097,N28098,N28099,
  N28100,N28101,N28102,N28103,N28104,N28105,N28106,N28107,N28108,N28109,N28110,N28111,
  N28112,N28113,N28114,N28115,N28116,N28117,N28118,N28119,N28120,N28121,N28122,
  N28123,N28124,N28125,N28126,N28127,N28128,N28129,N28130,N28131,N28132,N28133,
  N28134,N28135,N28136,N28137,N28138,N28139,N28140,N28141,N28142,N28143,N28144,N28145,
  N28146,N28147,N28148,N28149,N28150,N28151,N28152,N28153,N28154,N28155,N28156,
  N28157,N28158,N28159,N28160,N28161,N28162,N28163,N28164,N28165,N28166,N28167,N28168,
  N28169,N28170,N28171,N28172,N28173,N28174,N28175,N28176,N28177,N28178,N28179,
  N28180,N28181,N28182,N28183,N28184,N28185,N28186,N28187,N28188,N28189,N28190,N28191,
  N28192,N28193,N28194,N28195,N28196,N28197,N28198,N28199,N28200,N28201,N28202,
  N28203,N28204,N28205,N28206,N28207,N28208,N28209,N28210,N28211,N28212,N28213,
  N28214,N28215,N28216,N28217,N28218,N28219,N28220,N28221,N28222,N28223,N28224,N28225,
  N28226,N28227,N28228,N28229,N28230,N28231,N28232,N28233,N28234,N28235,N28236,
  N28237,N28238,N28239,N28240,N28241,N28242,N28243,N28244,N28245,N28246,N28247,N28248,
  N28249,N28250,N28251,N28252,N28253,N28254,N28255,N28256,N28257,N28258,N28259,
  N28260,N28261,N28262,N28263,N28264,N28265,N28266,N28267,N28268,N28269,N28270,N28271,
  N28272,N28273,N28274,N28275,N28276,N28277,N28278,N28279,N28280,N28281,N28282,
  N28283,N28284,N28285,N28286,N28287,N28288,N28289,N28290,N28291,N28292,N28293,
  N28294,N28295,N28296,N28297,N28298,N28299,N28300,N28301,N28302,N28303,N28304,N28305,
  N28306,N28307,N28308,N28309,N28310,N28311,N28312,N28313,N28314,N28315,N28316,
  N28317,N28318,N28319,N28320,N28321,N28322,N28323,N28324,N28325,N28326,N28327,N28328,
  N28329,N28330,N28331,N28332,N28333,N28334,N28335,N28336,N28337,N28338,N28339,
  N28340,N28341,N28342,N28343,N28344,N28345,N28346,N28347,N28348,N28349,N28350,N28351,
  N28352,N28353,N28354,N28355,N28356,N28357,N28358,N28359,N28360,N28361,N28362,
  N28363,N28364,N28365,N28366,N28367,N28368,N28369,N28370,N28371,N28372,N28373,
  N28374,N28375,N28376,N28377,N28378,N28379,N28380,N28381,N28382,N28383,N28384,N28385,
  N28386,N28387,N28388,N28389,N28390,N28391,N28392,N28393,N28394,N28395,N28396,
  N28397,N28398,N28399,N28400,N28401,N28402,N28403,N28404,N28405,N28406,N28407,N28408,
  N28409,N28410,N28411,N28412,N28413,N28414,N28415,N28416,N28417,N28418,N28419,
  N28420,N28421,N28422,N28423,N28424,N28425,N28426,N28427,N28428,N28429,N28430,N28431,
  N28432,N28433,N28434,N28435,N28436,N28437,N28438,N28439,N28440,N28441,N28442,
  N28443,N28444,N28445,N28446,N28447,N28448,N28449,N28450,N28451,N28452,N28453,
  N28454,N28455,N28456,N28457,N28458,N28459,N28460,N28461,N28462,N28463,N28464,N28465,
  N28466,N28467,N28468,N28469,N28470,N28471,N28472,N28473,N28474,N28475,N28476,
  N28477,N28478,N28479,N28480,N28481,N28482,N28483,N28484,N28485,N28486,N28487,N28488,
  N28489,N28490,N28491,N28492,N28493,N28494,N28495,N28496,N28497,N28498,N28499,
  N28500,N28501,N28502,N28503,N28504,N28505,N28506,N28507,N28508,N28509,N28510,N28511,
  N28512,N28513,N28514,N28515,N28516,N28517,N28518,N28519,N28520,N28521,N28522,
  N28523,N28524,N28525,N28526,N28527,N28528,N28529,N28530,N28531,N28532,N28533,
  N28534,N28535,N28536,N28537,N28538,N28539,N28540,N28541,N28542,N28543,N28544,N28545,
  N28546,N28547,N28548,N28549,N28550,N28551,N28552,N28553,N28554,N28555,N28556,
  N28557,N28558,N28559,N28560,N28561,N28562,N28563,N28564,N28565,N28566,N28567,N28568,
  N28569,N28570,N28571,N28572,N28573,N28574,N28575,N28576,N28577,N28578,N28579,
  N28580,N28581,N28582,N28583,N28584,N28585,N28586,N28587,N28588,N28589,N28590,N28591,
  N28592,N28593,N28594,N28595,N28596,N28597,N28598,N28599,N28600,N28601,N28602,
  N28603,N28604,N28605,N28606,N28607,N28608,N28609,N28610,N28611,N28612,N28613,
  N28614,N28615,N28616,N28617,N28618,N28619,N28620,N28621,N28622,N28623,N28624,N28625,
  N28626,N28627,N28628,N28629,N28630,N28631,N28632,N28633,N28634,N28635,N28636,
  N28637,N28638,N28639,N28640,N28641,N28642,N28643,N28644,N28645,N28646,N28647,N28648,
  N28649,N28650,N28651,N28652,N28653,N28654,N28655,N28656,N28657,N28658,N28659,
  N28660,N28661,N28662,N28663,N28664,N28665,N28666,N28667,N28668,N28669,N28670,N28671,
  N28672,N28673,N28674,N28675,N28676,N28677,N28678,N28679,N28680,N28681,N28682,
  N28683,N28684,N28685,N28686,N28687,N28688,N28689,N28690,N28691,N28692,N28693,
  N28694,N28695,N28696,N28697,N28698,N28699,N28700,N28701,N28702,N28703,N28704,N28705,
  N28706,N28707,N28708,N28709,N28710,N28711,N28712,N28713,N28714,N28715,N28716,
  N28717,N28718,N28719,N28720,N28721,N28722,N28723,N28724,N28725,N28726,N28727,N28728,
  N28729,N28730,N28731,N28732,N28733,N28734,N28735,N28736,N28737,N28738,N28739,
  N28740,N28741,N28742,N28743,N28744,N28745,N28746,N28747,N28748,N28749,N28750,N28751,
  N28752,N28753,N28754,N28755,N28756,N28757,N28758,N28759,N28760,N28761,N28762,
  N28763,N28764,N28765,N28766,N28767,N28768,N28769,N28770,N28771,N28772,N28773,
  N28774,N28775,N28776,N28777,N28778,N28779,N28780,N28781,N28782,N28783,N28784,N28785,
  N28786,N28787,N28788,N28789,N28790,N28791,N28792,N28793,N28794,N28795,N28796,
  N28797,N28798,N28799,N28800,N28801,N28802,N28803,N28804,N28805,N28806,N28807,N28808,
  N28809,N28810,N28811,N28812,N28813,N28814,N28815,N28816,N28817,N28818,N28819,
  N28820,N28821,N28822,N28823,N28824,N28825,N28826,N28827,N28828,N28829,N28830,N28831,
  N28832,N28833,N28834,N28835,N28836,N28837,N28838,N28839,N28840,N28841,N28842,
  N28843,N28844,N28845,N28846,N28847,N28848,N28849,N28850,N28851,N28852,N28853,
  N28854,N28855,N28856,N28857,N28858,N28859,N28860,N28861,N28862,N28863,N28864,N28865,
  N28866,N28867,N28868,N28869,N28870,N28871,N28872,N28873,N28874,N28875,N28876,
  N28877,N28878,N28879,N28880,N28881,N28882,N28883,N28884,N28885,N28886,N28887,N28888,
  N28889,N28890,N28891,N28892,N28893,N28894,N28895,N28896,N28897,N28898,N28899,
  N28900,N28901,N28902,N28903,N28904,N28905,N28906,N28907,N28908,N28909,N28910,N28911,
  N28912,N28913,N28914,N28915,N28916,N28917,N28918,N28919,N28920,N28921,N28922,
  N28923,N28924,N28925,N28926,N28927,N28928,N28929,N28930,N28931,N28932,N28933,
  N28934,N28935,N28936,N28937,N28938,N28939,N28940,N28941,N28942,N28943,N28944,N28945,
  N28946,N28947,N28948,N28949,N28950,N28951,N28952,N28953,N28954,N28955,N28956,
  N28957,N28958,N28959,N28960,N28961,N28962,N28963,N28964,N28965,N28966,N28967,N28968,
  N28969,N28970,N28971,N28972,N28973,N28974,N28975,N28976,N28977,N28978,N28979,
  N28980,N28981,N28982,N28983,N28984,N28985,N28986,N28987,N28988,N28989,N28990,N28991,
  N28992,N28993,N28994,N28995,N28996,N28997,N28998,N28999,N29000,N29001,N29002,
  N29003,N29004,N29005,N29006,N29007,N29008,N29009,N29010,N29011,N29012,N29013,
  N29014,N29015,N29016,N29017,N29018,N29019,N29020,N29021,N29022,N29023,N29024,N29025,
  N29026,N29027,N29028,N29029,N29030,N29031,N29032,N29033,N29034,N29035,N29036,
  N29037,N29038,N29039,N29040,N29041,N29042,N29043,N29044,N29045,N29046,N29047,N29048,
  N29049,N29050,N29051,N29052,N29053,N29054,N29055,N29056,N29057,N29058,N29059,
  N29060,N29061,N29062,N29063,N29064,N29065,N29066,N29067,N29068,N29069,N29070,N29071,
  N29072,N29073,N29074,N29075,N29076,N29077,N29078,N29079,N29080,N29081,N29082,
  N29083,N29084,N29085,N29086,N29087,N29088,N29089,N29090,N29091,N29092,N29093,
  N29094,N29095,N29096,N29097,N29098,N29099,N29100,N29101,N29102,N29103,N29104,N29105,
  N29106,N29107,N29108,N29109,N29110,N29111,N29112,N29113,N29114,N29115,N29116,
  N29117,N29118,N29119,N29120,N29121,N29122,N29123,N29124,N29125,N29126,N29127,N29128,
  N29129,N29130,N29131,N29132,N29133,N29134,N29135,N29136,N29137,N29138,N29139,
  N29140,N29141,N29142,N29143,N29144,N29145,N29146,N29147,N29148,N29149,N29150,N29151,
  N29152,N29153,N29154,N29155,N29156,N29157,N29158,N29159,N29160,N29161,N29162,
  N29163,N29164,N29165,N29166,N29167,N29168,N29169,N29170,N29171,N29172,N29173,
  N29174,N29175,N29176,N29177,N29178,N29179,N29180,N29181,N29182,N29183,N29184,N29185,
  N29186,N29187,N29188,N29189,N29190,N29191,N29192,N29193,N29194,N29195,N29196,
  N29197,N29198,N29199,N29200,N29201,N29202,N29203,N29204,N29205,N29206,N29207,N29208,
  N29209,N29210,N29211,N29212,N29213,N29214,N29215,N29216,N29217,N29218,N29219,
  N29220,N29221,N29222,N29223,N29224,N29225,N29226,N29227,N29228,N29229,N29230,N29231,
  N29232,N29233,N29234,N29235,N29236,N29237,N29238,N29239,N29240,N29241,N29242,
  N29243,N29244,N29245,N29246,N29247,N29248,N29249,N29250,N29251,N29252,N29253,
  N29254,N29255,N29256,N29257,N29258,N29259,N29260,N29261,N29262,N29263,N29264,N29265,
  N29266,N29267,N29268,N29269,N29270,N29271,N29272,N29273,N29274,N29275,N29276,
  N29277,N29278,N29279,N29280,N29281,N29282,N29283,N29284,N29285,N29286,N29287,N29288,
  N29289,N29290,N29291,N29292,N29293,N29294,N29295,N29296,N29297,N29298,N29299,
  N29300,N29301,N29302,N29303,N29304,N29305,N29306,N29307,N29308,N29309,N29310,N29311,
  N29312,N29313,N29314,N29315,N29316,N29317,N29318,N29319,N29320,N29321,N29322,
  N29323,N29324,N29325,N29326,N29327,N29328,N29329,N29330,N29331,N29332,N29333,
  N29334,N29335,N29336,N29337,N29338,N29339,N29340,N29341,N29342,N29343,N29344,N29345,
  N29346,N29347,N29348,N29349,N29350,N29351,N29352,N29353,N29354,N29355,N29356,
  N29357,N29358,N29359,N29360,N29361,N29362,N29363,N29364,N29365,N29366,N29367,N29368,
  N29369,N29370,N29371,N29372,N29373,N29374,N29375,N29376,N29377,N29378,N29379,
  N29380,N29381,N29382,N29383,N29384,N29385,N29386,N29387,N29388,N29389,N29390,N29391,
  N29392,N29393,N29394,N29395,N29396,N29397,N29398,N29399,N29400,N29401,N29402,
  N29403,N29404,N29405,N29406,N29407,N29408,N29409,N29410,N29411,N29412,N29413,
  N29414,N29415,N29416,N29417,N29418,N29419,N29420,N29421,N29422,N29423,N29424,N29425,
  N29426,N29427,N29428,N29429,N29430,N29431,N29432,N29433,N29434,N29435,N29436,
  N29437,N29438,N29439,N29440,N29441,N29442,N29443,N29444,N29445,N29446,N29447,N29448,
  N29449,N29450,N29451,N29452,N29453,N29454,N29455,N29456,N29457,N29458,N29459,
  N29460,N29461,N29462,N29463,N29464,N29465,N29466,N29467,N29468,N29469,N29470,N29471,
  N29472,N29473,N29474,N29475,N29476,N29477,N29478,N29479,N29480,N29481,N29482,
  N29483,N29484,N29485,N29486,N29487,N29488,N29489,N29490,N29491,N29492,N29493,
  N29494,N29495,N29496,N29497,N29498,N29499,N29500,N29501,N29502,N29503,N29504,N29505,
  N29506,N29507,N29508,N29509,N29510,N29511,N29512,N29513,N29514,N29515,N29516,
  N29517,N29518,N29519,N29520,N29521,N29522,N29523,N29524,N29525,N29526,N29527,N29528,
  N29529,N29530,N29531,N29532,N29533,N29534,N29535,N29536,N29537,N29538,N29539,
  N29540,N29541,N29542,N29543,N29544,N29545,N29546,N29547,N29548,N29549,N29550,N29551,
  N29552,N29553,N29554,N29555,N29556,N29557,N29558,N29559,N29560,N29561,N29562,
  N29563,N29564,N29565,N29566,N29567,N29568,N29569,N29570,N29571,N29572,N29573,
  N29574,N29575,N29576,N29577,N29578,N29579,N29580,N29581,N29582,N29583,N29584,N29585,
  N29586,N29587,N29588,N29589,N29590,N29591,N29592,N29593,N29594,N29595,N29596,
  N29597,N29598,N29599,N29600,N29601,N29602,N29603,N29604,N29605,N29606,N29607,N29608,
  N29609,N29610,N29611,N29612,N29613,N29614,N29615,N29616,N29617,N29618,N29619,
  N29620,N29621,N29622,N29623,N29624,N29625,N29626,N29627,N29628,N29629,N29630,N29631,
  N29632,N29633,N29634,N29635,N29636,N29637,N29638,N29639,N29640,N29641,N29642,
  N29643,N29644,N29645,N29646,N29647,N29648,N29649,N29650,N29651,N29652,N29653,
  N29654,N29655,N29656,N29657,N29658,N29659,N29660,N29661,N29662,N29663,N29664,N29665,
  N29666,N29667,N29668,N29669,N29670,N29671,N29672,N29673,N29674,N29675,N29676,
  N29677,N29678,N29679,N29680,N29681,N29682,N29683,N29684,N29685,N29686,N29687,N29688,
  N29689,N29690,N29691,N29692,N29693,N29694,N29695,N29696,N29697,N29698,N29699,
  N29700,N29701,N29702,N29703,N29704,N29705,N29706,N29707,N29708,N29709,N29710,N29711,
  N29712,N29713,N29714,N29715,N29716,N29717,N29718,N29719,N29720,N29721,N29722,
  N29723,N29724,N29725,N29726,N29727,N29728,N29729,N29730,N29731,N29732,N29733,
  N29734,N29735,N29736,N29737,N29738,N29739,N29740,N29741,N29742,N29743,N29744,N29745,
  N29746,N29747,N29748,N29749,N29750,N29751,N29752,N29753,N29754,N29755,N29756,
  N29757,N29758,N29759,N29760,N29761,N29762,N29763,N29764,N29765,N29766,N29767,N29768,
  N29769,N29770,N29771,N29772,N29773,N29774,N29775,N29776,N29777,N29778,N29779,
  N29780,N29781,N29782,N29783,N29784,N29785,N29786,N29787,N29788,N29789,N29790,N29791,
  N29792,N29793,N29794,N29795,N29796,N29797,N29798,N29799,N29800,N29801,N29802,
  N29803,N29804,N29805,N29806,N29807,N29808,N29809,N29810,N29811,N29812,N29813,
  N29814,N29815,N29816,N29817,N29818,N29819,N29820,N29821,N29822,N29823,N29824,N29825,
  N29826,N29827,N29828,N29829,N29830,N29831,N29832,N29833,N29834,N29835,N29836,
  N29837,N29838,N29839,N29840,N29841,N29842,N29843,N29844,N29845,N29846,N29847,N29848,
  N29849,N29850,N29851,N29852,N29853,N29854,N29855,N29856,N29857,N29858,N29859,
  N29860,N29861,N29862,N29863,N29864,N29865,N29866,N29867,N29868,N29869,N29870,N29871,
  N29872,N29873,N29874,N29875,N29876,N29877,N29878,N29879,N29880,N29881,N29882,
  N29883,N29884,N29885,N29886,N29887,N29888,N29889,N29890,N29891,N29892,N29893,
  N29894,N29895,N29896,N29897,N29898,N29899,N29900,N29901,N29902,N29903,N29904,N29905,
  N29906,N29907,N29908,N29909,N29910,N29911,N29912,N29913,N29914,N29915,N29916,
  N29917,N29918,N29919,N29920,N29921,N29922,N29923,N29924,N29925,N29926,N29927,N29928,
  N29929,N29930,N29931,N29932,N29933,N29934,N29935,N29936,N29937,N29938,N29939,
  N29940,N29941,N29942,N29943,N29944,N29945,N29946,N29947,N29948,N29949,N29950,N29951,
  N29952,N29953,N29954,N29955,N29956,N29957,N29958,N29959,N29960,N29961,N29962,
  N29963,N29964,N29965,N29966,N29967,N29968,N29969,N29970,N29971,N29972,N29973,
  N29974,N29975,N29976,N29977,N29978,N29979,N29980,N29981,N29982,N29983,N29984,N29985,
  N29986,N29987,N29988,N29989,N29990,N29991,N29992,N29993,N29994,N29995,N29996,
  N29997,N29998,N29999,N30000,N30001,N30002,N30003,N30004,N30005,N30006,N30007,N30008,
  N30009,N30010,N30011,N30012,N30013,N30014,N30015,N30016,N30017,N30018,N30019,
  N30020,N30021,N30022,N30023,N30024,N30025,N30026,N30027,N30028,N30029,N30030,N30031,
  N30032,N30033,N30034,N30035,N30036,N30037,N30038,N30039,N30040,N30041,N30042,
  N30043,N30044,N30045,N30046,N30047,N30048,N30049,N30050,N30051,N30052,N30053,
  N30054,N30055,N30056,N30057,N30058,N30059,N30060,N30061,N30062,N30063,N30064,N30065,
  N30066,N30067,N30068,N30069,N30070,N30071,N30072,N30073,N30074,N30075,N30076,
  N30077,N30078,N30079,N30080,N30081,N30082,N30083,N30084,N30085,N30086,N30087,N30088,
  N30089,N30090,N30091,N30092,N30093,N30094,N30095,N30096,N30097,N30098,N30099,
  N30100,N30101,N30102,N30103,N30104,N30105,N30106,N30107,N30108,N30109,N30110,N30111,
  N30112,N30113,N30114,N30115,N30116,N30117,N30118,N30119,N30120,N30121,N30122,
  N30123,N30124,N30125,N30126,N30127,N30128,N30129,N30130,N30131,N30132,N30133,
  N30134,N30135,N30136,N30137,N30138,N30139,N30140,N30141,N30142,N30143,N30144,N30145,
  N30146,N30147,N30148,N30149,N30150,N30151,N30152,N30153,N30154,N30155,N30156,
  N30157,N30158,N30159,N30160,N30161,N30162,N30163,N30164,N30165,N30166,N30167,N30168,
  N30169,N30170,N30171,N30172,N30173,N30174,N30175,N30176,N30177,N30178,N30179,
  N30180,N30181,N30182,N30183,N30184,N30185,N30186,N30187,N30188,N30189,N30190,N30191,
  N30192,N30193,N30194,N30195,N30196,N30197,N30198,N30199,N30200,N30201,N30202,
  N30203,N30204,N30205,N30206,N30207,N30208,N30209,N30210,N30211,N30212,N30213,
  N30214,N30215,N30216,N30217,N30218,N30219,N30220,N30221,N30222,N30223,N30224,N30225,
  N30226,N30227,N30228,N30229,N30230,N30231,N30232,N30233,N30234,N30235,N30236,
  N30237,N30238,N30239,N30240,N30241,N30242,N30243,N30244,N30245,N30246,N30247,N30248,
  N30249,N30250,N30251,N30252,N30253,N30254,N30255,N30256,N30257,N30258,N30259,
  N30260,N30261,N30262,N30263,N30264,N30265,N30266,N30267,N30268,N30269,N30270,N30271,
  N30272,N30273,N30274,N30275,N30276,N30277,N30278,N30279,N30280,N30281,N30282,
  N30283,N30284,N30285,N30286,N30287,N30288,N30289,N30290,N30291,N30292,N30293,
  N30294,N30295,N30296,N30297,N30298,N30299,N30300,N30301,N30302,N30303,N30304,N30305,
  N30306,N30307,N30308,N30309,N30310,N30311,N30312,N30313,N30314,N30315,N30316,
  N30317,N30318,N30319,N30320,N30321,N30322,N30323,N30324,N30325,N30326,N30327,N30328,
  N30329,N30330,N30331,N30332,N30333,N30334,N30335,N30336,N30337,N30338,N30339,
  N30340,N30341,N30342,N30343,N30344,N30345,N30346,N30347,N30348,N30349,N30350,N30351,
  N30352,N30353,N30354,N30355,N30356,N30357,N30358,N30359,N30360,N30361,N30362,
  N30363,N30364,N30365,N30366,N30367,N30368,N30369,N30370,N30371,N30372,N30373,
  N30374,N30375,N30376,N30377,N30378,N30379,N30380,N30381,N30382,N30383,N30384,N30385,
  N30386,N30387,N30388,N30389,N30390,N30391,N30392,N30393,N30394,N30395,N30396,
  N30397,N30398,N30399,N30400,N30401,N30402,N30403,N30404,N30405,N30406,N30407,N30408,
  N30409,N30410,N30411,N30412,N30413,N30414,N30415,N30416,N30417,N30418,N30419,
  N30420,N30421,N30422,N30423,N30424,N30425,N30426,N30427,N30428,N30429,N30430,N30431,
  N30432,N30433,N30434,N30435,N30436,N30437,N30438,N30439,N30440,N30441,N30442,
  N30443,N30444,N30445,N30446,N30447,N30448,N30449,N30450,N30451,N30452,N30453,
  N30454,N30455,N30456,N30457,N30458,N30459,N30460,N30461,N30462,N30463,N30464,N30465,
  N30466,N30467,N30468,N30469,N30470,N30471,N30472,N30473,N30474,N30475,N30476,
  N30477,N30478,N30479,N30480,N30481,N30482,N30483,N30484,N30485,N30486,N30487,N30488,
  N30489,N30490,N30491,N30492,N30493,N30494,N30495,N30496,N30497,N30498,N30499,
  N30500,N30501,N30502,N30503,N30504,N30505,N30506,N30507,N30508,N30509,N30510,N30511,
  N30512,N30513,N30514,N30515,N30516,N30517,N30518,N30519,N30520,N30521,N30522,
  N30523,N30524,N30525,N30526,N30527,N30528,N30529,N30530,N30531,N30532,N30533,
  N30534,N30535,N30536,N30537,N30538,N30539,N30540,N30541,N30542,N30543,N30544,N30545,
  N30546,N30547,N30548,N30549,N30550,N30551,N30552,N30553,N30554,N30555,N30556,
  N30557,N30558,N30559,N30560,N30561,N30562,N30563,N30564,N30565,N30566,N30567,N30568,
  N30569,N30570,N30571,N30572,N30573,N30574,N30575,N30576,N30577,N30578,N30579,
  N30580,N30581,N30582,N30583,N30584,N30585,N30586,N30587,N30588,N30589,N30590,N30591,
  N30592,N30593,N30594,N30595,N30596,N30597,N30598,N30599,N30600,N30601,N30602,
  N30603,N30604,N30605,N30606,N30607,N30608,N30609,N30610,N30611,N30612,N30613,
  N30614,N30615,N30616,N30617,N30618,N30619,N30620,N30621,N30622,N30623,N30624,N30625,
  N30626,N30627,N30628,N30629,N30630,N30631,N30632,N30633,N30634,N30635,N30636,
  N30637,N30638,N30639,N30640,N30641,N30642,N30643,N30644,N30645,N30646,N30647,N30648,
  N30649,N30650,N30651,N30652,N30653,N30654,N30655,N30656,N30657,N30658,N30659,
  N30660,N30661,N30662,N30663,N30664,N30665,N30666,N30667,N30668,N30669,N30670,N30671,
  N30672,N30673,N30674,N30675,N30676,N30677,N30678,N30679,N30680,N30681,N30682,
  N30683,N30684,N30685,N30686,N30687,N30688,N30689,N30690,N30691,N30692,N30693,
  N30694,N30695,N30696,N30697,N30698,N30699,N30700,N30701,N30702,N30703,N30704,N30705,
  N30706,N30707,N30708,N30709,N30710,N30711,N30712,N30713,N30714,N30715,N30716,
  N30717,N30718,N30719,N30720,N30721,N30722,N30723,N30724,N30725,N30726,N30727,N30728,
  N30729,N30730,N30731,N30732,N30733,N30734,N30735,N30736,N30737,N30738,N30739,
  N30740,N30741,N30742,N30743,N30744,N30745,N30746,N30747,N30748,N30749,N30750,N30751,
  N30752,N30753,N30754,N30755,N30756,N30757,N30758,N30759,N30760,N30761,N30762,
  N30763,N30764,N30765,N30766,N30767,N30768,N30769,N30770,N30771,N30772,N30773,
  N30774,N30775,N30776,N30777,N30778,N30779,N30780,N30781,N30782,N30783,N30784,N30785,
  N30786,N30787,N30788,N30789,N30790,N30791,N30792,N30793,N30794,N30795,N30796,
  N30797,N30798,N30799,N30800,N30801,N30802,N30803,N30804,N30805,N30806,N30807,N30808,
  N30809,N30810,N30811,N30812,N30813,N30814,N30815,N30816,N30817,N30818,N30819,
  N30820,N30821,N30822,N30823,N30824,N30825,N30826,N30827,N30828,N30829,N30830,N30831,
  N30832,N30833,N30834,N30835,N30836,N30837,N30838,N30839,N30840,N30841,N30842,
  N30843,N30844,N30845,N30846,N30847,N30848,N30849,N30850,N30851,N30852,N30853,
  N30854,N30855,N30856,N30857,N30858,N30859,N30860,N30861,N30862,N30863,N30864,N30865,
  N30866,N30867,N30868,N30869,N30870,N30871,N30872,N30873,N30874,N30875,N30876,
  N30877,N30878,N30879,N30880,N30881,N30882,N30883,N30884,N30885,N30886,N30887,N30888,
  N30889,N30890,N30891,N30892,N30893,N30894,N30895,N30896,N30897,N30898,N30899,
  N30900,N30901,N30902,N30903,N30904,N30905,N30906,N30907,N30908,N30909,N30910,N30911,
  N30912,N30913,N30914,N30915,N30916,N30917,N30918,N30919,N30920,N30921,N30922,
  N30923,N30924,N30925,N30926,N30927,N30928,N30929,N30930,N30931,N30932,N30933,
  N30934,N30935,N30936,N30937,N30938,N30939,N30940,N30941,N30942,N30943,N30944,N30945,
  N30946,N30947,N30948,N30949,N30950,N30951,N30952,N30953,N30954,N30955,N30956,
  N30957,N30958,N30959,N30960,N30961,N30962,N30963,N30964,N30965,N30966,N30967,N30968,
  N30969,N30970,N30971,N30972,N30973,N30974,N30975,N30976,N30977,N30978,N30979,
  N30980,N30981,N30982,N30983,N30984,N30985,N30986,N30987,N30988,N30989,N30990,N30991,
  N30992,N30993,N30994,N30995,N30996,N30997,N30998,N30999,N31000,N31001,N31002,
  N31003,N31004,N31005,N31006,N31007,N31008,N31009,N31010,N31011,N31012,N31013,
  N31014,N31015,N31016,N31017,N31018,N31019,N31020,N31021,N31022,N31023,N31024,N31025,
  N31026,N31027,N31028,N31029,N31030,N31031,N31032,N31033,N31034,N31035,N31036,
  N31037,N31038,N31039,N31040,N31041,N31042,N31043,N31044,N31045,N31046,N31047,N31048,
  N31049,N31050,N31051,N31052,N31053,N31054,N31055,N31056,N31057,N31058,N31059,
  N31060,N31061,N31062,N31063,N31064,N31065,N31066,N31067,N31068,N31069,N31070,N31071,
  N31072,N31073,N31074,N31075,N31076,N31077,N31078,N31079,N31080,N31081,N31082,
  N31083,N31084,N31085,N31086,N31087,N31088,N31089,N31090,N31091,N31092,N31093,
  N31094,N31095,N31096,N31097,N31098,N31099,N31100,N31101,N31102,N31103,N31104,N31105,
  N31106,N31107,N31108,N31109,N31110,N31111,N31112,N31113,N31114,N31115,N31116,
  N31117,N31118,N31119,N31120,N31121,N31122,N31123,N31124,N31125,N31126,N31127,N31128,
  N31129,N31130,N31131,N31132,N31133,N31134,N31135,N31136,N31137,N31138,N31139,
  N31140,N31141,N31142,N31143,N31144,N31145,N31146,N31147,N31148,N31149,N31150,N31151,
  N31152,N31153,N31154,N31155,N31156,N31157,N31158,N31159,N31160,N31161,N31162,
  N31163,N31164,N31165,N31166,N31167,N31168,N31169,N31170,N31171,N31172,N31173,
  N31174,N31175,N31176,N31177,N31178,N31179,N31180,N31181,N31182,N31183,N31184,N31185,
  N31186,N31187,N31188,N31189,N31190,N31191,N31192,N31193,N31194,N31195,N31196,
  N31197,N31198,N31199,N31200,N31201,N31202,N31203,N31204,N31205,N31206,N31207,N31208,
  N31209,N31210,N31211,N31212,N31213,N31214,N31215,N31216,N31217,N31218,N31219,
  N31220,N31221,N31222,N31223,N31224,N31225,N31226,N31227,N31228,N31229,N31230,N31231,
  N31232,N31233,N31234,N31235,N31236,N31237,N31238,N31239,N31240,N31241,N31242,
  N31243,N31244,N31245,N31246,N31247,N31248,N31249,N31250,N31251,N31252,N31253,
  N31254,N31255,N31256,N31257,N31258,N31259,N31260,N31261,N31262,N31263,N31264,N31265,
  N31266,N31267,N31268,N31269,N31270,N31271,N31272,N31273,N31274,N31275,N31276,
  N31277,N31278,N31279,N31280,N31281,N31282,N31283,N31284,N31285,N31286,N31287,N31288,
  N31289,N31290,N31291,N31292,N31293,N31294,N31295,N31296,N31297,N31298,N31299,
  N31300,N31301,N31302,N31303,N31304,N31305,N31306,N31307,N31308,N31309,N31310,N31311,
  N31312,N31313,N31314,N31315,N31316,N31317,N31318,N31319,N31320,N31321,N31322,
  N31323,N31324,N31325,N31326,N31327,N31328,N31329,N31330,N31331,N31332,N31333,
  N31334,N31335,N31336,N31337,N31338,N31339,N31340,N31341,N31342,N31343,N31344,N31345,
  N31346,N31347,N31348,N31349,N31350,N31351,N31352,N31353,N31354,N31355,N31356,
  N31357,N31358,N31359,N31360,N31361,N31362,N31363,N31364,N31365,N31366,N31367,N31368,
  N31369,N31370,N31371,N31372,N31373,N31374,N31375,N31376,N31377,N31378,N31379,
  N31380,N31381,N31382,N31383,N31384,N31385,N31386,N31387,N31388,N31389,N31390,N31391,
  N31392,N31393,N31394,N31395,N31396,N31397,N31398,N31399,N31400,N31401,N31402,
  N31403,N31404,N31405,N31406,N31407,N31408,N31409,N31410,N31411,N31412,N31413,
  N31414,N31415,N31416,N31417,N31418,N31419,N31420,N31421,N31422,N31423,N31424,N31425,
  N31426,N31427,N31428,N31429,N31430,N31431,N31432,N31433,N31434,N31435,N31436,
  N31437,N31438,N31439,N31440,N31441,N31442,N31443,N31444,N31445,N31446,N31447,N31448,
  N31449,N31450,N31451,N31452,N31453,N31454,N31455,N31456,N31457,N31458,N31459,
  N31460,N31461,N31462,N31463,N31464,N31465,N31466,N31467,N31468,N31469,N31470,N31471,
  N31472,N31473,N31474,N31475,N31476,N31477,N31478,N31479,N31480,N31481,N31482,
  N31483,N31484,N31485,N31486,N31487,N31488,N31489,N31490,N31491,N31492,N31493,
  N31494,N31495,N31496,N31497,N31498,N31499,N31500,N31501,N31502,N31503,N31504,N31505,
  N31506,N31507,N31508,N31509,N31510,N31511,N31512,N31513,N31514,N31515,N31516,
  N31517,N31518,N31519,N31520,N31521,N31522,N31523,N31524,N31525,N31526,N31527,N31528,
  N31529,N31530,N31531,N31532,N31533,N31534,N31535,N31536,N31537,N31538,N31539,
  N31540,N31541,N31542,N31543,N31544,N31545,N31546,N31547,N31548,N31549,N31550,N31551,
  N31552,N31553,N31554,N31555,N31556,N31557,N31558,N31559,N31560,N31561,N31562,
  N31563,N31564,N31565,N31566,N31567,N31568,N31569,N31570,N31571,N31572,N31573,
  N31574,N31575,N31576,N31577,N31578,N31579,N31580,N31581,N31582,N31583,N31584,N31585,
  N31586,N31587,N31588,N31589,N31590,N31591,N31592,N31593,N31594,N31595,N31596,
  N31597,N31598,N31599,N31600,N31601,N31602,N31603,N31604,N31605,N31606,N31607,N31608,
  N31609,N31610,N31611,N31612,N31613,N31614,N31615,N31616,N31617,N31618,N31619,
  N31620,N31621,N31622,N31623,N31624,N31625,N31626,N31627,N31628,N31629,N31630,N31631,
  N31632,N31633,N31634,N31635,N31636,N31637,N31638,N31639,N31640,N31641,N31642,
  N31643,N31644,N31645,N31646,N31647,N31648,N31649,N31650,N31651,N31652,N31653,
  N31654,N31655,N31656,N31657,N31658,N31659,N31660,N31661,N31662,N31663,N31664,N31665,
  N31666,N31667,N31668,N31669,N31670,N31671,N31672,N31673,N31674,N31675,N31676,
  N31677,N31678,N31679,N31680,N31681,N31682,N31683,N31684,N31685,N31686,N31687,N31688,
  N31689,N31690,N31691,N31692,N31693,N31694,N31695,N31696,N31697,N31698,N31699,
  N31700,N31701,N31702,N31703,N31704,N31705,N31706,N31707,N31708,N31709,N31710,N31711,
  N31712,N31713,N31714,N31715,N31716,N31717,N31718,N31719,N31720,N31721,N31722,
  N31723,N31724,N31725,N31726,N31727,N31728,N31729,N31730,N31731,N31732,N31733,
  N31734,N31735,N31736,N31737,N31738,N31739,N31740,N31741,N31742,N31743,N31744,N31745,
  N31746,N31747,N31748,N31749,N31750,N31751,N31752,N31753,N31754,N31755,N31756,
  N31757,N31758,N31759,N31760,N31761,N31762,N31763,N31764,N31765,N31766,N31767,N31768,
  N31769,N31770,N31771,N31772,N31773,N31774,N31775,N31776,N31777,N31778,N31779,
  N31780,N31781,N31782,N31783,N31784,N31785,N31786,N31787,N31788,N31789,N31790,N31791,
  N31792,N31793,N31794,N31795,N31796,N31797,N31798,N31799,N31800,N31801,N31802,
  N31803,N31804,N31805,N31806,N31807,N31808,N31809,N31810,N31811,N31812,N31813,
  N31814,N31815,N31816,N31817,N31818,N31819,N31820,N31821,N31822,N31823,N31824,N31825,
  N31826,N31827,N31828,N31829,N31830,N31831,N31832,N31833,N31834,N31835,N31836,
  N31837,N31838,N31839,N31840,N31841,N31842,N31843,N31844,N31845,N31846,N31847,N31848,
  N31849,N31850,N31851,N31852,N31853,N31854,N31855,N31856,N31857,N31858,N31859,
  N31860,N31861,N31862,N31863,N31864,N31865,N31866,N31867,N31868,N31869,N31870,N31871,
  N31872,N31873,N31874,N31875,N31876,N31877,N31878,N31879,N31880,N31881,N31882,
  N31883,N31884,N31885,N31886,N31887,N31888,N31889,N31890,N31891,N31892,N31893,
  N31894,N31895,N31896,N31897,N31898,N31899,N31900,N31901,N31902,N31903,N31904,N31905,
  N31906,N31907,N31908,N31909,N31910,N31911,N31912,N31913,N31914,N31915,N31916,
  N31917,N31918,N31919,N31920,N31921,N31922,N31923,N31924,N31925,N31926,N31927,N31928,
  N31929,N31930,N31931,N31932,N31933,N31934,N31935,N31936,N31937,N31938,N31939,
  N31940,N31941,N31942,N31943,N31944,N31945,N31946,N31947,N31948,N31949,N31950,N31951,
  N31952,N31953,N31954,N31955,N31956,N31957,N31958,N31959,N31960,N31961,N31962,
  N31963,N31964,N31965,N31966,N31967,N31968,N31969,N31970,N31971,N31972,N31973,
  N31974,N31975,N31976,N31977,N31978,N31979,N31980,N31981,N31982,N31983,N31984,N31985,
  N31986,N31987,N31988,N31989,N31990,N31991,N31992,N31993,N31994,N31995,N31996,
  N31997,N31998,N31999,N32000,N32001,N32002,N32003,N32004,N32005,N32006,N32007,N32008,
  N32009,N32010,N32011,N32012,N32013,N32014,N32015,N32016,N32017,N32018,N32019,
  N32020,N32021,N32022,N32023,N32024,N32025,N32026,N32027,N32028,N32029,N32030,N32031,
  N32032,N32033,N32034,N32035,N32036,N32037,N32038,N32039,N32040,N32041,N32042,
  N32043,N32044,N32045,N32046,N32047,N32048,N32049,N32050,N32051,N32052,N32053,
  N32054,N32055,N32056,N32057,N32058,N32059,N32060,N32061,N32062,N32063,N32064,N32065,
  N32066,N32067,N32068,N32069,N32070,N32071,N32072,N32073,N32074,N32075,N32076,
  N32077,N32078,N32079,N32080,N32081,N32082,N32083,N32084,N32085,N32086,N32087,N32088,
  N32089,N32090,N32091,N32092,N32093,N32094,N32095,N32096,N32097,N32098,N32099,
  N32100,N32101,N32102,N32103,N32104,N32105,N32106,N32107,N32108,N32109,N32110,N32111,
  N32112,N32113,N32114,N32115,N32116,N32117,N32118,N32119,N32120,N32121,N32122,
  N32123,N32124,N32125,N32126,N32127,N32128,N32129,N32130,N32131,N32132,N32133,
  N32134,N32135,N32136,N32137,N32138,N32139,N32140,N32141,N32142,N32143,N32144,N32145,
  N32146,N32147,N32148,N32149,N32150,N32151,N32152,N32153,N32154,N32155,N32156,
  N32157,N32158,N32159,N32160,N32161,N32162,N32163,N32164,N32165,N32166,N32167,N32168,
  N32169,N32170,N32171,N32172,N32173,N32174,N32175,N32176,N32177,N32178,N32179,
  N32180,N32181,N32182,N32183,N32184,N32185,N32186,N32187,N32188,N32189,N32190,N32191,
  N32192,N32193,N32194,N32195,N32196,N32197,N32198,N32199,N32200,N32201,N32202,
  N32203,N32204,N32205,N32206,N32207,N32208,N32209,N32210,N32211,N32212,N32213,
  N32214,N32215,N32216,N32217,N32218,N32219,N32220,N32221,N32222,N32223,N32224,N32225,
  N32226,N32227,N32228,N32229,N32230,N32231,N32232,N32233,N32234,N32235,N32236,
  N32237,N32238,N32239,N32240,N32241,N32242,N32243,N32244,N32245,N32246,N32247,N32248,
  N32249,N32250,N32251,N32252,N32253,N32254,N32255,N32256,N32257,N32258,N32259,
  N32260,N32261,N32262,N32263,N32264,N32265,N32266,N32267,N32268,N32269,N32270,N32271,
  N32272,N32273,N32274,N32275,N32276,N32277,N32278,N32279,N32280,N32281,N32282,
  N32283,N32284,N32285,N32286,N32287,N32288,N32289,N32290,N32291,N32292,N32293,
  N32294,N32295,N32296,N32297,N32298,N32299,N32300,N32301,N32302,N32303,N32304,N32305,
  N32306,N32307,N32308,N32309,N32310,N32311,N32312,N32313,N32314,N32315,N32316,
  N32317,N32318,N32319,N32320,N32321,N32322,N32323,N32324,N32325,N32326,N32327,N32328,
  N32329,N32330,N32331,N32332,N32333,N32334,N32335,N32336,N32337,N32338,N32339,
  N32340,N32341,N32342,N32343,N32344,N32345,N32346,N32347,N32348,N32349,N32350,N32351,
  N32352,N32353,N32354,N32355,N32356,N32357,N32358,N32359,N32360,N32361,N32362,
  N32363,N32364,N32365,N32366,N32367,N32368,N32369,N32370,N32371,N32372,N32373,
  N32374,N32375,N32376,N32377,N32378,N32379,N32380,N32381,N32382,N32383,N32384,N32385,
  N32386,N32387,N32388,N32389,N32390,N32391,N32392,N32393,N32394,N32395,N32396,
  N32397,N32398,N32399,N32400,N32401,N32402,N32403,N32404,N32405,N32406,N32407,N32408,
  N32409,N32410,N32411,N32412,N32413,N32414,N32415,N32416,N32417,N32418,N32419,
  N32420,N32421,N32422,N32423,N32424,N32425,N32426,N32427,N32428,N32429,N32430,N32431,
  N32432,N32433,N32434,N32435,N32436,N32437,N32438,N32439,N32440,N32441,N32442,
  N32443,N32444,N32445,N32446,N32447,N32448,N32449,N32450,N32451,N32452,N32453,
  N32454,N32455,N32456,N32457,N32458,N32459,N32460,N32461,N32462,N32463,N32464,N32465,
  N32466,N32467,N32468,N32469,N32470,N32471,N32472,N32473,N32474,N32475,N32476,
  N32477,N32478,N32479,N32480,N32481,N32482,N32483,N32484,N32485,N32486,N32487,N32488,
  N32489,N32490,N32491,N32492,N32493,N32494,N32495,N32496,N32497,N32498,N32499,
  N32500,N32501,N32502,N32503,N32504,N32505,N32506,N32507,N32508,N32509,N32510,N32511,
  N32512,N32513,N32514,N32515,N32516,N32517,N32518,N32519,N32520,N32521,N32522,
  N32523,N32524,N32525,N32526,N32527,N32528,N32529,N32530,N32531,N32532,N32533,
  N32534,N32535,N32536,N32537,N32538,N32539,N32540,N32541,N32542,N32543,N32544,N32545,
  N32546,N32547,N32548,N32549,N32550,N32551,N32552,N32553,N32554,N32555,N32556,
  N32557,N32558,N32559,N32560,N32561,N32562,N32563,N32564,N32565,N32566,N32567,N32568,
  N32569,N32570,N32571,N32572,N32573,N32574,N32575,N32576,N32577,N32578,N32579,
  N32580,N32581,N32582,N32583,N32584,N32585,N32586,N32587,N32588,N32589,N32590,N32591,
  N32592,N32593,N32594,N32595,N32596,N32597,N32598,N32599,N32600,N32601,N32602,
  N32603,N32604,N32605,N32606,N32607,N32608,N32609,N32610,N32611,N32612,N32613,
  N32614,N32615,N32616,N32617,N32618,N32619,N32620,N32621,N32622,N32623,N32624,N32625,
  N32626,N32627,N32628,N32629,N32630,N32631,N32632,N32633,N32634,N32635,N32636,
  N32637,N32638,N32639,N32640,N32641,N32642,N32643,N32644,N32645,N32646,N32647,N32648,
  N32649,N32650,N32651,N32652,N32653,N32654,N32655,N32656,N32657,N32658,N32659,
  N32660,N32661,N32662,N32663,N32664,N32665,N32666,N32667,N32668,N32669,N32670,N32671,
  N32672,N32673,N32674,N32675,N32676,N32677,N32678,N32679,N32680,N32681,N32682,
  N32683,N32684,N32685,N32686,N32687,N32688,N32689,N32690,N32691,N32692,N32693,
  N32694,N32695,N32696,N32697,N32698,N32699,N32700,N32701,N32702,N32703,N32704,N32705,
  N32706,N32707,N32708,N32709,N32710,N32711,N32712,N32713,N32714,N32715,N32716,
  N32717,N32718,N32719,N32720,N32721,N32722,N32723,N32724,N32725,N32726,N32727,N32728,
  N32729,N32730,N32731,N32732,N32733,N32734,N32735,N32736,N32737,N32738,N32739,
  N32740,N32741,N32742,N32743,N32744,N32745,N32746,N32747,N32748,N32749,N32750,N32751,
  N32752,N32753,N32754,N32755,N32756,N32757,N32758,N32759,N32760,N32761,N32762,
  N32763,N32764,N32765,N32766,N32767,N32768,N32769,N32770,N32771,N32772,N32773,
  N32774,N32775,N32776,N32777,N32778,N32779,N32780,N32781,N32782,N32783,N32784,N32785,
  N32786,N32787,N32788,N32789,N32790,N32791,N32792,N32793,N32794,N32795,N32796,
  N32797,N32798,N32799,N32800,N32801,N32802,N32803,N32804,N32805,N32806,N32807,N32808,
  N32809,N32810,N32811,N32812,N32813,N32814,N32815,N32816,N32817,N32818,N32819,
  N32820,N32821,N32822,N32823,N32824,N32825,N32826,N32827,N32828,N32829,N32830,N32831,
  N32832,N32833,N32834,N32835,N32836,N32837,N32838,N32839,N32840,N32841,N32842,
  N32843,N32844,N32845,N32846,N32847,N32848,N32849,N32850,N32851,N32852,N32853,
  N32854,N32855,N32856,N32857,N32858,N32859,N32860,N32861,N32862,N32863,N32864,N32865,
  N32866,N32867,N32868,N32869,N32870,N32871,N32872,N32873,N32874,N32875,N32876,
  N32877,N32878,N32879,N32880,N32881,N32882,N32883,N32884,N32885,N32886,N32887,N32888,
  N32889,N32890,N32891,N32892,N32893,N32894,N32895,N32896,N32897,N32898,N32899,
  N32900,N32901,N32902,N32903,N32904,N32905,N32906,N32907,N32908,N32909,N32910,N32911,
  N32912,N32913,N32914,N32915,N32916,N32917,N32918,N32919,N32920,N32921,N32922,
  N32923,N32924,N32925,N32926,N32927,N32928,N32929,N32930,N32931,N32932,N32933,
  N32934,N32935,N32936,N32937,N32938,N32939,N32940,N32941,N32942,N32943,N32944,N32945,
  N32946,N32947,N32948,N32949,N32950,N32951,N32952,N32953,N32954,N32955,N32956,
  N32957,N32958,N32959,N32960,N32961,N32962,N32963,N32964,N32965,N32966,N32967,N32968,
  N32969,N32970,N32971,N32972,N32973,N32974,N32975,N32976,N32977,N32978,N32979,
  N32980,N32981,N32982,N32983,N32984,N32985,N32986,N32987,N32988,N32989,N32990,N32991,
  N32992,N32993,N32994,N32995,N32996,N32997,N32998,N32999,N33000,N33001,N33002,
  N33003,N33004,N33005,N33006,N33007,N33008,N33009,N33010,N33011,N33012,N33013,
  N33014,N33015,N33016,N33017,N33018,N33019,N33020,N33021,N33022,N33023,N33024,N33025,
  N33026,N33027,N33028,N33029,N33030,N33031,N33032,N33033,N33034,N33035,N33036,
  N33037,N33038,N33039,N33040,N33041,N33042,N33043,N33044,N33045,N33046,N33047,N33048,
  N33049,N33050,N33051,N33052,N33053,N33054,N33055,N33056,N33057,N33058,N33059,
  N33060,N33061,N33062,N33063,N33064,N33065,N33066,N33067,N33068,N33069,N33070,N33071,
  N33072,N33073,N33074,N33075,N33076,N33077,N33078,N33079,N33080,N33081,N33082,
  N33083,N33084,N33085,N33086,N33087,N33088,N33089,N33090,N33091,N33092,N33093,
  N33094,N33095,N33096,N33097,N33098,N33099,N33100,N33101,N33102,N33103,N33104,N33105,
  N33106,N33107,N33108,N33109,N33110,N33111,N33112,N33113,N33114,N33115,N33116,
  N33117,N33118,N33119,N33120,N33121,N33122,N33123,N33124,N33125,N33126,N33127,N33128,
  N33129,N33130,N33131,N33132,N33133,N33134,N33135,N33136,N33137,N33138,N33139,
  N33140,N33141,N33142,N33143,N33144,N33145,N33146,N33147,N33148,N33149,N33150,N33151,
  N33152,N33153,N33154,N33155,N33156,N33157,N33158,N33159,N33160,N33161,N33162,
  N33163,N33164,N33165,N33166,N33167,N33168,N33169,N33170,N33171,N33172,N33173,
  N33174,N33175,N33176,N33177,N33178,N33179,N33180,N33181,N33182,N33183,N33184,N33185,
  N33186,N33187,N33188,N33189,N33190,N33191,N33192,N33193,N33194,N33195,N33196,
  N33197,N33198,N33199,N33200,N33201,N33202,N33203,N33204,N33205,N33206,N33207,N33208,
  N33209,N33210,N33211,N33212,N33213,N33214,N33215,N33216,N33217,N33218,N33219,
  N33220,N33221,N33222,N33223,N33224,N33225,N33226,N33227,N33228,N33229,N33230,N33231,
  N33232,N33233,N33234,N33235,N33236,N33237,N33238,N33239,N33240,N33241,N33242,
  N33243,N33244,N33245,N33246,N33247,N33248,N33249,N33250,N33251,N33252,N33253,
  N33254,N33255,N33256,N33257,N33258,N33259,N33260,N33261,N33262,N33263,N33264,N33265,
  N33266,N33267,N33268,N33269,N33270,N33271,N33272,N33273,N33274,N33275,N33276,
  N33277,N33278,N33279,N33280,N33281,N33282,N33283,N33284,N33285,N33286,N33287,N33288,
  N33289,N33290,N33291,N33292,N33293,N33294,N33295,N33296,N33297,N33298,N33299,
  N33300,N33301,N33302,N33303,N33304,N33305,N33306,N33307,N33308,N33309,N33310,N33311,
  N33312,N33313,N33314,N33315,N33316,N33317,N33318,N33319,N33320,N33321,N33322,
  N33323,N33324,N33325,N33326,N33327,N33328,N33329,N33330,N33331,N33332,N33333,
  N33334,N33335,N33336,N33337,N33338,N33339,N33340,N33341,N33342,N33343,N33344,N33345,
  N33346,N33347,N33348,N33349,N33350,N33351,N33352,N33353,N33354,N33355,N33356,
  N33357,N33358,N33359,N33360,N33361,N33362,N33363,N33364,N33365,N33366,N33367,N33368,
  N33369,N33370,N33371,N33372,N33373,N33374,N33375,N33376,N33377,N33378,N33379,
  N33380,N33381,N33382,N33383,N33384,N33385,N33386,N33387,N33388,N33389,N33390,N33391,
  N33392,N33393,N33394,N33395,N33396,N33397,N33398,N33399,N33400,N33401,N33402,
  N33403,N33404,N33405,N33406,N33407,N33408,N33409,N33410,N33411,N33412,N33413,
  N33414,N33415,N33416,N33417,N33418,N33419,N33420,N33421,N33422,N33423,N33424,N33425,
  N33426,N33427,N33428,N33429,N33430,N33431,N33432,N33433,N33434,N33435,N33436,
  N33437,N33438,N33439,N33440,N33441,N33442,N33443,N33444,N33445,N33446,N33447,N33448,
  N33449,N33450,N33451,N33452,N33453,N33454,N33455,N33456,N33457,N33458,N33459,
  N33460,N33461,N33462,N33463,N33464,N33465,N33466,N33467,N33468,N33469,N33470,N33471,
  N33472,N33473,N33474,N33475,N33476,N33477,N33478,N33479,N33480,N33481,N33482,
  N33483,N33484,N33485,N33486,N33487,N33488,N33489,N33490,N33491,N33492,N33493,
  N33494,N33495,N33496,N33497,N33498,N33499,N33500,N33501,N33502,N33503,N33504,N33505,
  N33506,N33507,N33508,N33509,N33510,N33511,N33512,N33513,N33514,N33515,N33516,
  N33517,N33518,N33519,N33520,N33521,N33522,N33523,N33524,N33525,N33526,N33527,N33528,
  N33529,N33530,N33531,N33532,N33533,N33534,N33535,N33536,N33537,N33538,N33539,
  N33540,N33541,N33542,N33543,N33544,N33545,N33546,N33547,N33548,N33549,N33550,N33551,
  N33552,N33553,N33554,N33555,N33556,N33557,N33558,N33559,N33560,N33561,N33562,
  N33563,N33564,N33565,N33566,N33567,N33568,N33569,N33570,N33571,N33572,N33573,
  N33574,N33575,N33576,N33577,N33578,N33579,N33580,N33581,N33582,N33583,N33584,N33585,
  N33586,N33587,N33588,N33589,N33590,N33591,N33592,N33593,N33594,N33595,N33596,
  N33597,N33598,N33599,N33600,N33601,N33602,N33603,N33604,N33605,N33606,N33607,N33608,
  N33609,N33610,N33611,N33612,N33613,N33614,N33615,N33616,N33617,N33618,N33619,
  N33620,N33621,N33622,N33623,N33624,N33625,N33626,N33627,N33628,N33629,N33630,N33631,
  N33632,N33633,N33634,N33635,N33636,N33637,N33638,N33639,N33640,N33641,N33642,
  N33643,N33644,N33645,N33646,N33647,N33648,N33649,N33650,N33651,N33652,N33653,
  N33654,N33655,N33656,N33657,N33658,N33659,N33660,N33661,N33662,N33663,N33664,N33665,
  N33666,N33667,N33668,N33669,N33670,N33671,N33672,N33673,N33674,N33675,N33676,
  N33677,N33678,N33679,N33680,N33681,N33682,N33683,N33684,N33685,N33686,N33687,N33688,
  N33689,N33690,N33691,N33692,N33693,N33694,N33695,N33696,N33697,N33698,N33699,
  N33700,N33701,N33702,N33703,N33704,N33705,N33706,N33707,N33708,N33709,N33710,N33711,
  N33712,N33713,N33714,N33715,N33716,N33717,N33718,N33719,N33720,N33721,N33722,
  N33723,N33724,N33725,N33726,N33727,N33728,N33729,N33730,N33731,N33732,N33733,
  N33734,N33735,N33736,N33737,N33738,N33739,N33740,N33741,N33742,N33743,N33744,N33745,
  N33746,N33747,N33748,N33749,N33750,N33751,N33752,N33753,N33754,N33755,N33756,
  N33757,N33758,N33759,N33760,N33761,N33762,N33763,N33764,N33765,N33766,N33767,N33768,
  N33769,N33770,N33771,N33772,N33773,N33774,N33775,N33776,N33777,N33778,N33779,
  N33780,N33781,N33782,N33783,N33784,N33785,N33786,N33787,N33788,N33789,N33790,N33791,
  N33792,N33793,N33794,N33795,N33796,N33797,N33798,N33799,N33800,N33801,N33802,
  N33803,N33804,N33805,N33806,N33807,N33808,N33809,N33810,N33811,N33812,N33813,
  N33814,N33815,N33816,N33817,N33818,N33819,N33820,N33821,N33822,N33823,N33824,N33825,
  N33826,N33827,N33828,N33829,N33830,N33831,N33832,N33833,N33834,N33835,N33836,
  N33837,N33838,N33839,N33840,N33841,N33842,N33843,N33844,N33845,N33846,N33847,N33848,
  N33849,N33850,N33851,N33852,N33853,N33854,N33855,N33856,N33857,N33858,N33859,
  N33860,N33861,N33862,N33863,N33864,N33865,N33866,N33867,N33868,N33869,N33870,N33871,
  N33872,N33873,N33874,N33875,N33876,N33877,N33878,N33879,N33880,N33881,N33882,
  N33883,N33884,N33885,N33886,N33887,N33888,N33889,N33890,N33891,N33892,N33893,
  N33894,N33895,N33896,N33897,N33898,N33899,N33900,N33901,N33902,N33903,N33904,N33905,
  N33906,N33907,N33908,N33909,N33910,N33911,N33912,N33913,N33914,N33915,N33916,
  N33917,N33918,N33919,N33920,N33921,N33922,N33923,N33924,N33925,N33926,N33927,N33928,
  N33929,N33930,N33931,N33932,N33933,N33934,N33935,N33936,N33937,N33938,N33939,
  N33940,N33941,N33942,N33943,N33944,N33945,N33946,N33947,N33948,N33949,N33950,N33951,
  N33952,N33953,N33954,N33955,N33956,N33957,N33958,N33959,N33960,N33961,N33962,
  N33963,N33964,N33965,N33966,N33967,N33968,N33969,N33970,N33971,N33972,N33973,
  N33974,N33975,N33976,N33977,N33978,N33979,N33980,N33981,N33982,N33983,N33984,N33985,
  N33986,N33987,N33988,N33989,N33990,N33991,N33992,N33993,N33994,N33995,N33996,
  N33997,N33998,N33999,N34000,N34001,N34002,N34003,N34004,N34005,N34006,N34007,N34008,
  N34009,N34010,N34011,N34012,N34013,N34014,N34015,N34016,N34017,N34018,N34019,
  N34020,N34021,N34022,N34023,N34024,N34025,N34026,N34027,N34028,N34029,N34030,N34031,
  N34032,N34033,N34034,N34035,N34036,N34037,N34038,N34039,N34040,N34041,N34042,
  N34043,N34044,N34045,N34046,N34047,N34048,N34049,N34050,N34051,N34052,N34053,
  N34054,N34055,N34056,N34057,N34058,N34059,N34060,N34061,N34062,N34063,N34064,N34065,
  N34066,N34067,N34068,N34069,N34070,N34071,N34072,N34073,N34074,N34075,N34076,
  N34077,N34078,N34079,N34080,N34081,N34082,N34083,N34084,N34085,N34086,N34087,N34088,
  N34089,N34090,N34091,N34092,N34093,N34094,N34095,N34096,N34097,N34098,N34099,
  N34100,N34101,N34102,N34103,N34104,N34105,N34106,N34107,N34108,N34109,N34110,N34111,
  N34112,N34113,N34114,N34115,N34116,N34117,N34118,N34119,N34120,N34121,N34122,
  N34123,N34124,N34125,N34126,N34127,N34128,N34129,N34130,N34131,N34132,N34133,
  N34134,N34135,N34136,N34137,N34138,N34139,N34140,N34141,N34142,N34143,N34144,N34145,
  N34146,N34147,N34148,N34149,N34150,N34151,N34152,N34153,N34154,N34155,N34156,
  N34157,N34158,N34159,N34160,N34161,N34162,N34163,N34164,N34165,N34166,N34167,N34168,
  N34169,N34170,N34171,N34172,N34173,N34174,N34175,N34176,N34177,N34178,N34179,
  N34180,N34181,N34182,N34183,N34184,N34185,N34186,N34187,N34188,N34189,N34190,N34191,
  N34192,N34193,N34194,N34195,N34196,N34197,N34198,N34199,N34200,N34201,N34202,
  N34203,N34204,N34205,N34206,N34207,N34208,N34209,N34210,N34211,N34212,N34213,
  N34214,N34215,N34216,N34217,N34218,N34219,N34220,N34221,N34222,N34223,N34224,N34225,
  N34226,N34227,N34228,N34229,N34230,N34231,N34232,N34233,N34234,N34235,N34236,
  N34237,N34238,N34239,N34240,N34241,N34242,N34243,N34244,N34245,N34246,N34247,N34248,
  N34249,N34250,N34251,N34252,N34253,N34254,N34255,N34256,N34257,N34258,N34259,
  N34260,N34261,N34262,N34263,N34264,N34265,N34266,N34267,N34268,N34269,N34270,N34271,
  N34272,N34273,N34274,N34275,N34276,N34277,N34278,N34279,N34280,N34281,N34282,
  N34283,N34284,N34285,N34286,N34287,N34288,N34289,N34290,N34291,N34292,N34293,
  N34294,N34295,N34296,N34297,N34298,N34299,N34300,N34301,N34302,N34303,N34304,N34305,
  N34306,N34307,N34308,N34309,N34310,N34311,N34312,N34313,N34314,N34315,N34316,
  N34317,N34318,N34319,N34320,N34321,N34322,N34323,N34324,N34325,N34326,N34327,N34328,
  N34329,N34330,N34331,N34332,N34333,N34334,N34335,N34336,N34337,N34338,N34339,
  N34340,N34341,N34342,N34343,N34344,N34345,N34346,N34347,N34348,N34349,N34350,N34351,
  N34352,N34353,N34354,N34355,N34356,N34357,N34358,N34359,N34360,N34361,N34362,
  N34363,N34364,N34365,N34366,N34367,N34368,N34369,N34370,N34371,N34372,N34373,
  N34374,N34375,N34376,N34377,N34378,N34379,N34380,N34381,N34382,N34383,N34384,N34385,
  N34386,N34387,N34388,N34389,N34390,N34391,N34392,N34393,N34394,N34395,N34396,
  N34397,N34398,N34399,N34400,N34401,N34402,N34403,N34404,N34405,N34406,N34407,N34408,
  N34409,N34410,N34411,N34412,N34413,N34414,N34415,N34416,N34417,N34418,N34419,
  N34420,N34421,N34422,N34423,N34424,N34425,N34426,N34427,N34428,N34429,N34430,N34431,
  N34432,N34433,N34434,N34435,N34436,N34437,N34438,N34439,N34440,N34441,N34442,
  N34443,N34444,N34445,N34446,N34447,N34448,N34449,N34450,N34451,N34452,N34453,
  N34454,N34455,N34456,N34457,N34458,N34459,N34460,N34461,N34462,N34463,N34464,N34465,
  N34466,N34467,N34468,N34469,N34470,N34471,N34472,N34473,N34474,N34475,N34476,
  N34477,N34478,N34479,N34480,N34481,N34482,N34483,N34484,N34485,N34486,N34487,N34488,
  N34489,N34490,N34491,N34492,N34493,N34494,N34495,N34496,N34497,N34498,N34499,
  N34500,N34501,N34502,N34503,N34504,N34505,N34506,N34507,N34508,N34509,N34510,N34511,
  N34512,N34513,N34514,N34515,N34516,N34517,N34518,N34519,N34520,N34521,N34522,
  N34523,N34524,N34525,N34526,N34527,N34528,N34529,N34530,N34531,N34532,N34533,
  N34534,N34535,N34536,N34537,N34538,N34539,N34540,N34541,N34542,N34543,N34544,N34545,
  N34546,N34547,N34548,N34549,N34550,N34551,N34552,N34553,N34554,N34555,N34556,
  N34557,N34558,N34559,N34560,N34561,N34562,N34563,N34564,N34565,N34566,N34567,N34568,
  N34569,N34570,N34571,N34572,N34573,N34574,N34575,N34576,N34577,N34578,N34579,
  N34580,N34581,N34582,N34583,N34584,N34585,N34586,N34587,N34588,N34589,N34590,N34591,
  N34592,N34593,N34594,N34595,N34596,N34597,N34598,N34599,N34600,N34601,N34602,
  N34603,N34604,N34605,N34606,N34607,N34608,N34609,N34610,N34611,N34612,N34613,
  N34614,N34615,N34616,N34617,N34618,N34619,N34620,N34621,N34622,N34623,N34624,N34625,
  N34626,N34627,N34628,N34629,N34630,N34631,N34632,N34633,N34634,N34635,N34636,
  N34637,N34638,N34639,N34640,N34641,N34642,N34643,N34644,N34645,N34646,N34647,N34648,
  N34649,N34650,N34651,N34652,N34653,N34654,N34655,N34656,N34657,N34658,N34659,
  N34660,N34661,N34662,N34663,N34664,N34665,N34666,N34667,N34668,N34669,N34670,N34671,
  N34672,N34673,N34674,N34675,N34676,N34677,N34678,N34679,N34680,N34681,N34682,
  N34683,N34684,N34685,N34686,N34687,N34688,N34689,N34690,N34691,N34692,N34693,
  N34694,N34695,N34696,N34697,N34698,N34699,N34700,N34701,N34702,N34703,N34704,N34705,
  N34706,N34707,N34708,N34709,N34710,N34711,N34712,N34713,N34714,N34715,N34716,
  N34717,N34718,N34719,N34720,N34721,N34722,N34723,N34724,N34725,N34726,N34727,N34728,
  N34729,N34730,N34731,N34732,N34733,N34734,N34735,N34736,N34737,N34738,N34739,
  N34740,N34741,N34742,N34743,N34744,N34745,N34746,N34747,N34748,N34749,N34750,N34751,
  N34752,N34753,N34754,N34755,N34756,N34757,N34758,N34759,N34760,N34761,N34762,
  N34763,N34764,N34765,N34766,N34767,N34768,N34769,N34770,N34771,N34772,N34773,
  N34774,N34775,N34776,N34777,N34778,N34779,N34780,N34781,N34782,N34783,N34784,N34785,
  N34786,N34787,N34788,N34789,N34790,N34791,N34792,N34793,N34794,N34795,N34796,
  N34797,N34798,N34799,N34800,N34801,N34802,N34803,N34804,N34805,N34806,N34807,N34808,
  N34809,N34810,N34811,N34812,N34813,N34814,N34815,N34816,N34817,N34818,N34819,
  N34820,N34821,N34822,N34823,N34824,N34825,N34826,N34827,N34828,N34829,N34830,N34831,
  N34832,N34833,N34834,N34835,N34836,N34837,N34838,N34839,N34840,N34841,N34842,
  N34843,N34844,N34845,N34846,N34847,N34848,N34849,N34850,N34851,N34852,N34853,
  N34854,N34855,N34856,N34857,N34858,N34859,N34860,N34861,N34862,N34863,N34864,N34865,
  N34866,N34867,N34868,N34869,N34870,N34871,N34872,N34873,N34874,N34875,N34876,
  N34877,N34878,N34879,N34880,N34881,N34882,N34883,N34884,N34885,N34886,N34887,N34888,
  N34889,N34890,N34891,N34892,N34893,N34894,N34895,N34896,N34897,N34898,N34899,
  N34900,N34901,N34902,N34903,N34904,N34905,N34906,N34907,N34908,N34909,N34910,N34911,
  N34912,N34913,N34914,N34915,N34916,N34917,N34918,N34919,N34920,N34921,N34922,
  N34923,N34924,N34925,N34926,N34927,N34928,N34929,N34930,N34931,N34932,N34933,
  N34934,N34935,N34936,N34937,N34938,N34939,N34940,N34941,N34942,N34943,N34944,N34945,
  N34946,N34947,N34948,N34949,N34950,N34951,N34952,N34953,N34954,N34955,N34956,
  N34957,N34958,N34959,N34960,N34961,N34962,N34963,N34964,N34965,N34966,N34967,N34968,
  N34969,N34970,N34971,N34972,N34973,N34974,N34975,N34976,N34977,N34978,N34979,
  N34980,N34981,N34982,N34983,N34984,N34985,N34986,N34987,N34988,N34989,N34990,N34991,
  N34992,N34993,N34994,N34995,N34996,N34997,N34998,N34999,N35000,N35001,N35002,
  N35003,N35004,N35005,N35006,N35007,N35008,N35009,N35010,N35011,N35012,N35013,
  N35014,N35015,N35016,N35017,N35018,N35019,N35020,N35021,N35022,N35023,N35024,N35025,
  N35026,N35027,N35028,N35029,N35030,N35031,N35032,N35033,N35034,N35035,N35036,
  N35037,N35038,N35039,N35040,N35041,N35042,N35043,N35044,N35045,N35046,N35047,N35048,
  N35049,N35050,N35051,N35052,N35053,N35054,N35055,N35056,N35057,N35058,N35059,
  N35060,N35061,N35062,N35063,N35064,N35065,N35066,N35067,N35068,N35069,N35070,N35071,
  N35072,N35073,N35074,N35075,N35076,N35077,N35078,N35079,N35080,N35081,N35082,
  N35083,N35084,N35085,N35086,N35087,N35088,N35089,N35090,N35091,N35092,N35093,
  N35094,N35095,N35096,N35097,N35098,N35099,N35100,N35101,N35102,N35103,N35104,N35105,
  N35106,N35107,N35108,N35109,N35110,N35111,N35112,N35113,N35114,N35115,N35116,
  N35117,N35118,N35119,N35120,N35121,N35122,N35123,N35124,N35125,N35126,N35127,N35128,
  N35129,N35130,N35131,N35132,N35133,N35134,N35135,N35136,N35137,N35138,N35139,
  N35140,N35141,N35142,N35143,N35144,N35145,N35146,N35147,N35148,N35149,N35150,N35151,
  N35152,N35153,N35154,N35155,N35156,N35157,N35158,N35159,N35160,N35161,N35162,
  N35163,N35164,N35165,N35166,N35167,N35168,N35169,N35170,N35171,N35172,N35173,
  N35174,N35175,N35176,N35177,N35178,N35179,N35180,N35181,N35182,N35183,N35184,N35185,
  N35186,N35187,N35188,N35189,N35190,N35191,N35192,N35193,N35194,N35195,N35196,
  N35197,N35198,N35199,N35200,N35201,N35202,N35203,N35204,N35205,N35206,N35207,N35208,
  N35209,N35210,N35211,N35212,N35213,N35214,N35215,N35216,N35217,N35218,N35219,
  N35220,N35221,N35222,N35223,N35224,N35225,N35226,N35227,N35228,N35229,N35230,N35231,
  N35232,N35233,N35234,N35235,N35236,N35237,N35238,N35239,N35240,N35241,N35242,
  N35243,N35244,N35245,N35246,N35247,N35248,N35249,N35250,N35251,N35252,N35253,
  N35254,N35255,N35256,N35257,N35258,N35259,N35260,N35261,N35262,N35263,N35264,N35265,
  N35266,N35267,N35268,N35269,N35270,N35271,N35272,N35273,N35274,N35275,N35276,
  N35277,N35278,N35279,N35280,N35281,N35282,N35283,N35284,N35285,N35286,N35287,N35288,
  N35289,N35290,N35291,N35292,N35293,N35294,N35295,N35296,N35297,N35298,N35299,
  N35300,N35301,N35302,N35303,N35304,N35305,N35306,N35307,N35308,N35309,N35310,N35311,
  N35312,N35313,N35314,N35315,N35316,N35317,N35318,N35319,N35320,N35321,N35322,
  N35323,N35324,N35325,N35326,N35327,N35328,N35329,N35330,N35331,N35332,N35333,
  N35334,N35335,N35336,N35337,N35338,N35339,N35340,N35341,N35342,N35343,N35344,N35345,
  N35346,N35347,N35348,N35349,N35350,N35351,N35352,N35353,N35354,N35355,N35356,
  N35357,N35358,N35359,N35360,N35361,N35362,N35363,N35364,N35365,N35366,N35367,N35368,
  N35369,N35370,N35371,N35372,N35373,N35374,N35375,N35376,N35377,N35378,N35379,
  N35380,N35381,N35382,N35383,N35384,N35385,N35386,N35387,N35388,N35389,N35390,N35391,
  N35392,N35393,N35394,N35395,N35396,N35397,N35398,N35399,N35400,N35401,N35402,
  N35403,N35404,N35405,N35406,N35407,N35408,N35409,N35410,N35411,N35412,N35413,
  N35414,N35415,N35416,N35417,N35418,N35419,N35420,N35421,N35422,N35423,N35424,N35425,
  N35426,N35427,N35428,N35429,N35430,N35431,N35432,N35433,N35434,N35435,N35436,
  N35437,N35438,N35439,N35440,N35441,N35442,N35443,N35444,N35445,N35446,N35447,N35448,
  N35449,N35450,N35451,N35452,N35453,N35454,N35455,N35456,N35457,N35458,N35459,
  N35460,N35461,N35462,N35463,N35464,N35465,N35466,N35467,N35468,N35469,N35470,N35471,
  N35472,N35473,N35474,N35475,N35476,N35477,N35478,N35479,N35480,N35481,N35482,
  N35483,N35484,N35485,N35486,N35487,N35488,N35489,N35490,N35491,N35492,N35493,
  N35494,N35495,N35496,N35497,N35498,N35499,N35500,N35501,N35502,N35503,N35504,N35505,
  N35506,N35507,N35508,N35509,N35510,N35511,N35512,N35513,N35514,N35515,N35516,
  N35517,N35518,N35519,N35520,N35521,N35522,N35523,N35524,N35525,N35526,N35527,N35528,
  N35529,N35530,N35531,N35532,N35533,N35534,N35535,N35536,N35537,N35538,N35539,
  N35540,N35541,N35542,N35543,N35544,N35545,N35546,N35547,N35548,N35549,N35550,N35551,
  N35552,N35553,N35554,N35555,N35556,N35557,N35558,N35559,N35560,N35561,N35562,
  N35563,N35564,N35565,N35566,N35567,N35568,N35569,N35570,N35571,N35572,N35573,
  N35574,N35575,N35576,N35577,N35578,N35579,N35580,N35581,N35582,N35583,N35584,N35585,
  N35586,N35587,N35588,N35589,N35590,N35591,N35592,N35593,N35594,N35595,N35596,
  N35597,N35598,N35599,N35600,N35601,N35602,N35603,N35604,N35605,N35606,N35607,N35608,
  N35609,N35610,N35611,N35612,N35613,N35614,N35615,N35616,N35617,N35618,N35619,
  N35620,N35621,N35622,N35623,N35624,N35625,N35626,N35627,N35628,N35629,N35630,N35631,
  N35632,N35633,N35634,N35635,N35636,N35637,N35638,N35639,N35640,N35641,N35642,
  N35643,N35644,N35645,N35646,N35647,N35648,N35649,N35650,N35651,N35652,N35653,
  N35654,N35655,N35656,N35657,N35658,N35659,N35660,N35661,N35662,N35663,N35664,N35665,
  N35666,N35667,N35668,N35669,N35670,N35671,N35672,N35673,N35674,N35675,N35676,
  N35677,N35678,N35679,N35680,N35681,N35682,N35683,N35684,N35685,N35686,N35687,N35688,
  N35689,N35690,N35691,N35692,N35693,N35694,N35695,N35696,N35697,N35698,N35699,
  N35700,N35701,N35702,N35703,N35704,N35705,N35706,N35707,N35708,N35709,N35710,N35711,
  N35712,N35713,N35714,N35715,N35716,N35717,N35718,N35719,N35720,N35721,N35722,
  N35723,N35724,N35725,N35726,N35727,N35728,N35729,N35730,N35731,N35732,N35733,
  N35734,N35735,N35736,N35737,N35738,N35739,N35740,N35741,N35742,N35743,N35744,N35745,
  N35746,N35747,N35748,N35749,N35750,N35751,N35752,N35753,N35754,N35755,N35756,
  N35757,N35758,N35759,N35760,N35761,N35762,N35763,N35764,N35765,N35766,N35767,N35768,
  N35769,N35770,N35771,N35772,N35773,N35774,N35775,N35776,N35777,N35778,N35779,
  N35780,N35781,N35782,N35783,N35784,N35785,N35786,N35787,N35788,N35789,N35790,N35791,
  N35792,N35793,N35794,N35795,N35796,N35797,N35798,N35799,N35800,N35801,N35802,
  N35803,N35804,N35805,N35806,N35807,N35808,N35809,N35810,N35811,N35812,N35813,
  N35814,N35815,N35816,N35817,N35818,N35819,N35820,N35821,N35822,N35823,N35824,N35825,
  N35826,N35827,N35828,N35829,N35830,N35831,N35832,N35833,N35834,N35835,N35836,
  N35837,N35838,N35839,N35840,N35841,N35842,N35843,N35844,N35845,N35846,N35847,N35848,
  N35849,N35850,N35851,N35852,N35853,N35854,N35855,N35856,N35857,N35858,N35859,
  N35860,N35861,N35862,N35863,N35864,N35865,N35866,N35867,N35868,N35869,N35870,N35871,
  N35872,N35873,N35874,N35875,N35876,N35877,N35878,N35879,N35880,N35881,N35882,
  N35883,N35884,N35885,N35886,N35887,N35888,N35889,N35890,N35891,N35892,N35893,
  N35894,N35895,N35896,N35897,N35898,N35899,N35900,N35901,N35902,N35903,N35904,N35905,
  N35906,N35907,N35908,N35909,N35910,N35911,N35912,N35913,N35914,N35915,N35916,
  N35917,N35918,N35919,N35920,N35921,N35922,N35923,N35924,N35925,N35926,N35927,N35928,
  N35929,N35930,N35931,N35932,N35933,N35934,N35935,N35936,N35937,N35938,N35939,
  N35940,N35941,N35942,N35943,N35944,N35945,N35946,N35947,N35948,N35949,N35950,N35951,
  N35952,N35953,N35954,N35955,N35956,N35957,N35958,N35959,N35960,N35961,N35962,
  N35963,N35964,N35965,N35966,N35967,N35968,N35969,N35970,N35971,N35972,N35973,
  N35974,N35975,N35976,N35977,N35978,N35979,N35980,N35981,N35982,N35983,N35984,N35985,
  N35986,N35987,N35988,N35989,N35990,N35991,N35992,N35993,N35994,N35995,N35996,
  N35997,N35998,N35999,N36000,N36001,N36002,N36003,N36004,N36005,N36006,N36007,N36008,
  N36009,N36010,N36011,N36012,N36013,N36014,N36015,N36016,N36017,N36018,N36019,
  N36020,N36021,N36022,N36023,N36024,N36025,N36026,N36027,N36028,N36029,N36030,N36031,
  N36032,N36033,N36034,N36035,N36036,N36037,N36038,N36039,N36040,N36041,N36042,
  N36043,N36044,N36045,N36046,N36047,N36048,N36049,N36050,N36051,N36052,N36053,
  N36054,N36055,N36056,N36057,N36058,N36059,N36060,N36061,N36062,N36063,N36064,N36065,
  N36066,N36067,N36068,N36069,N36070,N36071,N36072,N36073,N36074,N36075,N36076,
  N36077,N36078,N36079,N36080,N36081,N36082,N36083,N36084,N36085,N36086,N36087,N36088,
  N36089,N36090,N36091,N36092,N36093,N36094,N36095,N36096,N36097,N36098,N36099,
  N36100,N36101,N36102,N36103,N36104,N36105,N36106,N36107,N36108,N36109,N36110,N36111,
  N36112,N36113,N36114,N36115,N36116,N36117,N36118,N36119,N36120,N36121,N36122,
  N36123,N36124,N36125,N36126,N36127,N36128,N36129,N36130,N36131,N36132,N36133,
  N36134,N36135,N36136,N36137,N36138,N36139,N36140,N36141,N36142,N36143,N36144,N36145,
  N36146,N36147,N36148,N36149,N36150,N36151,N36152,N36153,N36154,N36155,N36156,
  N36157,N36158,N36159,N36160,N36161,N36162,N36163,N36164,N36165,N36166,N36167,N36168,
  N36169,N36170,N36171,N36172,N36173,N36174,N36175,N36176,N36177,N36178,N36179,
  N36180,N36181,N36182,N36183,N36184,N36185,N36186,N36187,N36188,N36189,N36190,N36191,
  N36192,N36193,N36194,N36195,N36196,N36197,N36198,N36199,N36200,N36201,N36202,
  N36203,N36204,N36205,N36206,N36207,N36208,N36209,N36210,N36211,N36212,N36213,
  N36214,N36215,N36216,N36217,N36218,N36219,N36220,N36221,N36222,N36223,N36224,N36225,
  N36226,N36227,N36228,N36229,N36230,N36231,N36232,N36233,N36234,N36235,N36236,
  N36237,N36238,N36239,N36240,N36241,N36242,N36243,N36244,N36245,N36246,N36247,N36248,
  N36249,N36250,N36251,N36252,N36253,N36254,N36255,N36256,N36257,N36258,N36259,
  N36260,N36261,N36262,N36263,N36264,N36265,N36266,N36267,N36268,N36269,N36270,N36271,
  N36272,N36273,N36274,N36275,N36276,N36277,N36278,N36279,N36280,N36281,N36282,
  N36283,N36284,N36285,N36286,N36287,N36288,N36289,N36290,N36291,N36292,N36293,
  N36294,N36295,N36296,N36297,N36298,N36299,N36300,N36301,N36302,N36303,N36304,N36305,
  N36306,N36307,N36308,N36309,N36310,N36311,N36312,N36313,N36314,N36315,N36316,
  N36317,N36318,N36319,N36320,N36321,N36322,N36323,N36324,N36325,N36326,N36327,N36328,
  N36329,N36330,N36331,N36332,N36333,N36334,N36335,N36336,N36337,N36338,N36339,
  N36340,N36341,N36342,N36343,N36344,N36345,N36346,N36347,N36348,N36349,N36350,N36351,
  N36352,N36353,N36354,N36355,N36356,N36357,N36358,N36359,N36360,N36361,N36362,
  N36363,N36364,N36365,N36366,N36367,N36368,N36369,N36370,N36371,N36372,N36373,
  N36374,N36375,N36376,N36377,N36378,N36379,N36380,N36381,N36382,N36383,N36384,N36385,
  N36386,N36387,N36388,N36389,N36390,N36391,N36392,N36393,N36394,N36395,N36396,
  N36397,N36398,N36399,N36400,N36401,N36402,N36403,N36404,N36405,N36406,N36407,N36408,
  N36409,N36410,N36411,N36412,N36413,N36414,N36415,N36416,N36417,N36418,N36419,
  N36420,N36421,N36422,N36423,N36424,N36425,N36426,N36427,N36428,N36429,N36430,N36431,
  N36432,N36433,N36434,N36435,N36436,N36437,N36438,N36439,N36440,N36441,N36442,
  N36443,N36444,N36445,N36446,N36447,N36448,N36449,N36450,N36451,N36452,N36453,
  N36454,N36455,N36456,N36457,N36458,N36459,N36460,N36461,N36462,N36463,N36464,N36465,
  N36466,N36467,N36468,N36469,N36470,N36471,N36472,N36473,N36474,N36475,N36476,
  N36477,N36478,N36479,N36480,N36481,N36482,N36483,N36484,N36485,N36486,N36487,N36488,
  N36489,N36490,N36491,N36492,N36493,N36494,N36495,N36496,N36497,N36498,N36499,
  N36500,N36501,N36502,N36503,N36504,N36505,N36506,N36507,N36508,N36509,N36510,N36511,
  N36512,N36513,N36514,N36515,N36516,N36517,N36518,N36519,N36520,N36521,N36522,
  N36523,N36524,N36525,N36526,N36527,N36528,N36529,N36530,N36531,N36532,N36533,
  N36534,N36535,N36536,N36537,N36538,N36539,N36540,N36541,N36542,N36543,N36544,N36545,
  N36546,N36547,N36548,N36549,N36550,N36551,N36552,N36553,N36554,N36555,N36556,
  N36557,N36558,N36559,N36560,N36561,N36562,N36563,N36564,N36565,N36566,N36567,N36568,
  N36569,N36570,N36571,N36572,N36573,N36574,N36575,N36576,N36577,N36578,N36579,
  N36580,N36581,N36582,N36583,N36584,N36585,N36586,N36587,N36588,N36589,N36590,N36591,
  N36592,N36593,N36594,N36595,N36596,N36597,N36598,N36599,N36600,N36601,N36602,
  N36603,N36604,N36605,N36606,N36607,N36608,N36609,N36610,N36611,N36612,N36613,
  N36614,N36615,N36616,N36617,N36618,N36619,N36620,N36621,N36622,N36623,N36624,N36625,
  N36626,N36627,N36628,N36629,N36630,N36631,N36632,N36633,N36634,N36635,N36636,
  N36637,N36638,N36639,N36640,N36641,N36642,N36643,N36644,N36645,N36646,N36647,N36648,
  N36649,N36650,N36651,N36652,N36653,N36654,N36655,N36656,N36657,N36658,N36659,
  N36660,N36661,N36662,N36663,N36664,N36665,N36666,N36667,N36668,N36669,N36670,N36671,
  N36672,N36673,N36674,N36675,N36676,N36677,N36678,N36679,N36680,N36681,N36682,
  N36683,N36684,N36685,N36686,N36687,N36688,N36689,N36690,N36691,N36692,N36693,
  N36694,N36695,N36696,N36697,N36698,N36699,N36700,N36701,N36702,N36703,N36704,N36705,
  N36706,N36707,N36708,N36709,N36710,N36711,N36712,N36713,N36714,N36715,N36716,
  N36717,N36718,N36719,N36720,N36721,N36722,N36723,N36724,N36725,N36726,N36727,N36728,
  N36729,N36730,N36731,N36732,N36733,N36734,N36735,N36736,N36737,N36738,N36739,
  N36740,N36741,N36742,N36743,N36744,N36745,N36746,N36747,N36748,N36749,N36750,N36751,
  N36752,N36753,N36754,N36755,N36756,N36757,N36758,N36759,N36760,N36761,N36762,
  N36763,N36764,N36765,N36766,N36767,N36768,N36769,N36770,N36771,N36772,N36773,
  N36774,N36775,N36776,N36777,N36778,N36779,N36780,N36781,N36782,N36783,N36784,N36785,
  N36786,N36787,N36788,N36789,N36790,N36791,N36792,N36793,N36794,N36795,N36796,
  N36797,N36798,N36799,N36800,N36801,N36802,N36803,N36804,N36805,N36806,N36807,N36808,
  N36809,N36810,N36811,N36812,N36813,N36814,N36815,N36816,N36817,N36818,N36819,
  N36820,N36821,N36822,N36823,N36824,N36825,N36826,N36827,N36828,N36829,N36830,N36831,
  N36832,N36833,N36834,N36835,N36836,N36837,N36838,N36839,N36840,N36841,N36842,
  N36843,N36844,N36845,N36846,N36847,N36848,N36849,N36850,N36851,N36852,N36853,
  N36854,N36855,N36856,N36857,N36858,N36859,N36860,N36861,N36862,N36863,N36864,N36865,
  N36866,N36867,N36868,N36869,N36870,N36871,N36872,N36873,N36874,N36875,N36876,
  N36877,N36878,N36879,N36880,N36881,N36882,N36883,N36884,N36885,N36886,N36887,N36888,
  N36889,N36890,N36891,N36892,N36893,N36894,N36895,N36896,N36897,N36898,N36899,
  N36900,N36901,N36902,N36903,N36904,N36905,N36906,N36907,N36908,N36909,N36910,N36911,
  N36912,N36913,N36914,N36915,N36916,N36917,N36918,N36919,N36920,N36921,N36922,
  N36923,N36924,N36925,N36926,N36927,N36928,N36929,N36930,N36931,N36932,N36933,
  N36934,N36935,N36936,N36937,N36938,N36939,N36940,N36941,N36942,N36943,N36944,N36945,
  N36946,N36947,N36948,N36949,N36950,N36951,N36952,N36953,N36954,N36955,N36956,
  N36957,N36958,N36959,N36960,N36961,N36962,N36963,N36964,N36965,N36966,N36967,N36968,
  N36969,N36970,N36971,N36972,N36973,N36974,N36975,N36976,N36977,N36978,N36979,
  N36980,N36981,N36982,N36983,N36984,N36985,N36986,N36987,N36988,N36989,N36990,N36991,
  N36992,N36993,N36994,N36995,N36996,N36997,N36998,N36999,N37000,N37001,N37002,
  N37003,N37004,N37005,N37006,N37007,N37008,N37009,N37010,N37011,N37012,N37013,
  N37014,N37015,N37016,N37017,N37018,N37019,N37020,N37021,N37022,N37023,N37024,N37025,
  N37026,N37027,N37028,N37029,N37030,N37031,N37032,N37033,N37034,N37035,N37036,
  N37037,N37038,N37039,N37040,N37041,N37042,N37043,N37044,N37045,N37046,N37047,N37048,
  N37049,N37050,N37051,N37052,N37053,N37054,N37055,N37056,N37057,N37058,N37059,
  N37060,N37061,N37062,N37063,N37064,N37065,N37066,N37067,N37068,N37069,N37070,N37071,
  N37072,N37073,N37074,N37075,N37076,N37077,N37078,N37079,N37080,N37081,N37082,
  N37083,N37084,N37085,N37086,N37087,N37088,N37089,N37090,N37091,N37092,N37093,
  N37094,N37095,N37096,N37097,N37098,N37099,N37100,N37101,N37102,N37103,N37104,N37105,
  N37106,N37107,N37108,N37109,N37110,N37111,N37112,N37113,N37114,N37115,N37116,
  N37117,N37118,N37119,N37120,N37121,N37122,N37123,N37124,N37125,N37126,N37127,N37128,
  N37129,N37130,N37131,N37132,N37133,N37134,N37135,N37136,N37137,N37138,N37139,
  N37140,N37141,N37142,N37143,N37144,N37145,N37146,N37147,N37148,N37149,N37150,N37151,
  N37152,N37153,N37154,N37155,N37156,N37157,N37158,N37159,N37160,N37161,N37162,
  N37163,N37164,N37165,N37166,N37167,N37168,N37169,N37170,N37171,N37172,N37173,
  N37174,N37175,N37176,N37177,N37178,N37179,N37180,N37181,N37182,N37183,N37184,N37185,
  N37186,N37187,N37188,N37189,N37190,N37191,N37192,N37193,N37194,N37195,N37196,
  N37197,N37198,N37199,N37200,N37201,N37202,N37203,N37204,N37205,N37206,N37207,N37208,
  N37209,N37210,N37211,N37212,N37213,N37214,N37215,N37216,N37217,N37218,N37219,
  N37220,N37221,N37222,N37223,N37224,N37225,N37226,N37227,N37228,N37229,N37230,N37231,
  N37232,N37233,N37234,N37235,N37236,N37237,N37238,N37239,N37240,N37241,N37242,
  N37243,N37244,N37245,N37246,N37247,N37248,N37249,N37250,N37251,N37252,N37253,
  N37254,N37255,N37256,N37257,N37258,N37259,N37260,N37261,N37262,N37263,N37264,N37265,
  N37266,N37267,N37268,N37269,N37270,N37271,N37272,N37273,N37274,N37275,N37276,
  N37277,N37278,N37279,N37280,N37281,N37282,N37283,N37284,N37285,N37286,N37287,N37288,
  N37289,N37290,N37291,N37292,N37293,N37294,N37295,N37296,N37297,N37298,N37299,
  N37300,N37301,N37302,N37303,N37304,N37305,N37306,N37307,N37308,N37309,N37310,N37311,
  N37312,N37313,N37314,N37315,N37316,N37317,N37318,N37319,N37320,N37321,N37322,
  N37323,N37324,N37325,N37326,N37327,N37328,N37329,N37330,N37331,N37332,N37333,
  N37334,N37335,N37336,N37337,N37338,N37339,N37340,N37341,N37342,N37343,N37344,N37345,
  N37346,N37347,N37348,N37349,N37350,N37351,N37352,N37353,N37354,N37355,N37356,
  N37357,N37358,N37359,N37360,N37361,N37362,N37363,N37364,N37365,N37366,N37367,N37368,
  N37369,N37370,N37371,N37372,N37373,N37374,N37375,N37376,N37377,N37378,N37379,
  N37380,N37381,N37382,N37383,N37384,N37385,N37386,N37387,N37388,N37389,N37390,N37391,
  N37392,N37393,N37394,N37395,N37396,N37397,N37398,N37399,N37400,N37401,N37402,
  N37403,N37404,N37405,N37406,N37407,N37408,N37409,N37410,N37411,N37412,N37413,
  N37414,N37415,N37416,N37417,N37418,N37419,N37420,N37421,N37422,N37423,N37424,N37425,
  N37426,N37427,N37428,N37429,N37430,N37431,N37432,N37433,N37434,N37435,N37436,
  N37437,N37438,N37439,N37440,N37441,N37442,N37443,N37444,N37445,N37446,N37447,N37448,
  N37449,N37450,N37451,N37452,N37453,N37454,N37455,N37456,N37457,N37458,N37459,
  N37460,N37461,N37462,N37463,N37464,N37465,N37466,N37467,N37468,N37469,N37470,N37471,
  N37472,N37473,N37474,N37475,N37476,N37477,N37478,N37479,N37480,N37481,N37482,
  N37483,N37484,N37485,N37486,N37487,N37488,N37489,N37490,N37491,N37492,N37493,
  N37494,N37495,N37496,N37497,N37498,N37499,N37500,N37501,N37502,N37503,N37504,N37505,
  N37506,N37507,N37508,N37509,N37510,N37511,N37512,N37513,N37514,N37515,N37516,
  N37517,N37518,N37519,N37520,N37521,N37522,N37523,N37524,N37525,N37526,N37527,N37528,
  N37529,N37530,N37531,N37532,N37533,N37534,N37535,N37536,N37537,N37538,N37539,
  N37540,N37541,N37542,N37543,N37544,N37545,N37546,N37547,N37548,N37549,N37550,N37551,
  N37552,N37553,N37554,N37555,N37556,N37557,N37558,N37559,N37560,N37561,N37562,
  N37563,N37564,N37565,N37566,N37567,N37568,N37569,N37570,N37571,N37572,N37573,
  N37574,N37575,N37576,N37577,N37578,N37579,N37580,N37581,N37582,N37583,N37584,N37585,
  N37586,N37587,N37588,N37589,N37590,N37591,N37592,N37593,N37594,N37595,N37596,
  N37597,N37598,N37599,N37600,N37601,N37602,N37603,N37604,N37605,N37606,N37607,N37608,
  N37609,N37610,N37611,N37612,N37613,N37614,N37615,N37616,N37617,N37618,N37619,
  N37620,N37621,N37622,N37623,N37624,N37625,N37626,N37627,N37628,N37629,N37630,N37631,
  N37632,N37633,N37634,N37635,N37636,N37637,N37638,N37639,N37640,N37641,N37642,
  N37643,N37644,N37645,N37646,N37647,N37648,N37649,N37650,N37651,N37652,N37653,
  N37654,N37655,N37656,N37657,N37658,N37659,N37660,N37661,N37662,N37663,N37664,N37665,
  N37666,N37667,N37668,N37669,N37670,N37671,N37672,N37673,N37674,N37675,N37676,
  N37677,N37678,N37679,N37680,N37681,N37682,N37683,N37684,N37685,N37686,N37687,N37688,
  N37689,N37690,N37691,N37692,N37693,N37694,N37695,N37696,N37697,N37698,N37699,
  N37700,N37701,N37702,N37703,N37704,N37705,N37706,N37707,N37708,N37709,N37710,N37711,
  N37712,N37713,N37714,N37715,N37716,N37717,N37718,N37719,N37720,N37721,N37722,
  N37723,N37724,N37725,N37726,N37727,N37728,N37729,N37730,N37731,N37732,N37733,
  N37734,N37735,N37736,N37737,N37738,N37739,N37740,N37741,N37742,N37743,N37744,N37745,
  N37746,N37747,N37748,N37749,N37750,N37751,N37752,N37753,N37754,N37755,N37756,
  N37757,N37758,N37759,N37760,N37761,N37762,N37763,N37764,N37765,N37766,N37767,N37768,
  N37769,N37770,N37771,N37772,N37773,N37774,N37775,N37776,N37777,N37778,N37779,
  N37780,N37781,N37782,N37783,N37784,N37785,N37786,N37787,N37788,N37789,N37790,N37791,
  N37792,N37793,N37794,N37795,N37796,N37797,N37798,N37799,N37800,N37801,N37802,
  N37803,N37804,N37805,N37806,N37807,N37808,N37809,N37810,N37811,N37812,N37813,
  N37814,N37815,N37816,N37817,N37818,N37819,N37820,N37821,N37822,N37823,N37824,N37825,
  N37826,N37827,N37828,N37829,N37830,N37831,N37832,N37833,N37834,N37835,N37836,
  N37837,N37838,N37839,N37840,N37841,N37842,N37843,N37844,N37845,N37846,N37847,N37848,
  N37849,N37850,N37851,N37852,N37853,N37854,N37855,N37856,N37857,N37858,N37859,
  N37860,N37861,N37862,N37863,N37864,N37865,N37866,N37867,N37868,N37869,N37870,N37871,
  N37872,N37873,N37874,N37875,N37876,N37877,N37878,N37879,N37880,N37881,N37882,
  N37883,N37884,N37885,N37886,N37887,N37888,N37889,N37890,N37891,N37892,N37893,
  N37894,N37895,N37896,N37897,N37898,N37899,N37900,N37901,N37902,N37903,N37904,N37905,
  N37906,N37907,N37908,N37909,N37910,N37911,N37912,N37913,N37914,N37915,N37916,
  N37917,N37918,N37919,N37920,N37921,N37922,N37923,N37924,N37925,N37926,N37927,N37928,
  N37929,N37930,N37931,N37932,N37933,N37934,N37935,N37936,N37937,N37938,N37939,
  N37940,N37941,N37942,N37943,N37944,N37945,N37946,N37947,N37948,N37949,N37950,N37951,
  N37952,N37953,N37954,N37955,N37956,N37957,N37958,N37959,N37960,N37961,N37962,
  N37963,N37964,N37965,N37966,N37967,N37968,N37969,N37970,N37971,N37972,N37973,
  N37974,N37975,N37976,N37977,N37978,N37979,N37980,N37981,N37982,N37983,N37984,N37985,
  N37986,N37987,N37988,N37989,N37990,N37991,N37992,N37993,N37994,N37995,N37996,
  N37997,N37998,N37999,N38000,N38001,N38002,N38003,N38004,N38005,N38006,N38007,N38008,
  N38009,N38010,N38011,N38012,N38013,N38014,N38015,N38016,N38017,N38018,N38019,
  N38020,N38021,N38022,N38023,N38024,N38025,N38026,N38027,N38028,N38029,N38030,N38031,
  N38032,N38033,N38034,N38035,N38036,N38037,N38038,N38039,N38040,N38041,N38042,
  N38043,N38044,N38045,N38046,N38047,N38048,N38049,N38050,N38051,N38052,N38053,
  N38054,N38055,N38056,N38057,N38058,N38059,N38060,N38061,N38062,N38063,N38064,N38065,
  N38066,N38067,N38068,N38069,N38070,N38071,N38072,N38073,N38074,N38075,N38076,
  N38077,N38078,N38079,N38080,N38081,N38082,N38083,N38084,N38085,N38086,N38087,N38088,
  N38089,N38090,N38091,N38092,N38093,N38094,N38095,N38096,N38097,N38098,N38099,
  N38100,N38101,N38102,N38103,N38104,N38105,N38106,N38107,N38108,N38109,N38110,N38111,
  N38112,N38113,N38114,N38115,N38116,N38117,N38118,N38119,N38120,N38121,N38122,
  N38123,N38124,N38125,N38126,N38127,N38128,N38129,N38130,N38131,N38132,N38133,
  N38134,N38135,N38136,N38137,N38138,N38139,N38140,N38141,N38142,N38143,N38144,N38145,
  N38146,N38147,N38148,N38149,N38150,N38151,N38152,N38153,N38154,N38155,N38156,
  N38157,N38158,N38159,N38160,N38161,N38162,N38163,N38164,N38165,N38166,N38167,N38168,
  N38169,N38170,N38171,N38172,N38173,N38174,N38175,N38176,N38177,N38178,N38179,
  N38180,N38181,N38182,N38183,N38184,N38185,N38186,N38187,N38188,N38189,N38190,N38191,
  N38192,N38193,N38194,N38195,N38196,N38197,N38198,N38199,N38200,N38201,N38202,
  N38203,N38204,N38205,N38206,N38207,N38208,N38209,N38210,N38211,N38212,N38213,
  N38214,N38215,N38216,N38217,N38218,N38219,N38220,N38221,N38222,N38223,N38224,N38225,
  N38226,N38227,N38228,N38229,N38230,N38231,N38232,N38233,N38234,N38235,N38236,
  N38237,N38238,N38239,N38240,N38241,N38242,N38243,N38244,N38245,N38246,N38247,N38248,
  N38249,N38250,N38251,N38252,N38253,N38254,N38255,N38256,N38257,N38258,N38259,
  N38260,N38261,N38262,N38263,N38264,N38265,N38266,N38267,N38268,N38269,N38270,N38271,
  N38272,N38273,N38274,N38275,N38276,N38277,N38278,N38279,N38280,N38281,N38282,
  N38283,N38284,N38285,N38286,N38287,N38288,N38289,N38290,N38291,N38292,N38293,
  N38294,N38295,N38296,N38297,N38298,N38299,N38300,N38301,N38302,N38303,N38304,N38305,
  N38306,N38307,N38308,N38309,N38310,N38311,N38312,N38313,N38314,N38315,N38316,
  N38317,N38318,N38319,N38320,N38321,N38322,N38323,N38324,N38325,N38326,N38327,N38328,
  N38329,N38330,N38331,N38332,N38333,N38334,N38335,N38336,N38337,N38338,N38339,
  N38340,N38341,N38342,N38343,N38344,N38345,N38346,N38347,N38348,N38349,N38350,N38351,
  N38352,N38353,N38354,N38355,N38356,N38357,N38358,N38359,N38360,N38361,N38362,
  N38363,N38364,N38365,N38366,N38367,N38368,N38369,N38370,N38371,N38372,N38373,
  N38374,N38375,N38376,N38377,N38378,N38379,N38380,N38381,N38382,N38383,N38384,N38385,
  N38386,N38387,N38388,N38389,N38390,N38391,N38392,N38393,N38394,N38395,N38396,
  N38397,N38398,N38399,N38400,N38401,N38402,N38403,N38404,N38405,N38406,N38407,N38408,
  N38409,N38410,N38411,N38412,N38413,N38414,N38415,N38416,N38417,N38418,N38419,
  N38420,N38421,N38422,N38423,N38424,N38425,N38426,N38427,N38428,N38429,N38430,N38431,
  N38432,N38433,N38434,N38435,N38436,N38437,N38438,N38439,N38440,N38441,N38442,
  N38443,N38444,N38445,N38446,N38447,N38448,N38449,N38450,N38451,N38452,N38453,
  N38454,N38455,N38456,N38457,N38458,N38459,N38460,N38461,N38462,N38463,N38464,N38465,
  N38466,N38467,N38468,N38469,N38470,N38471,N38472,N38473,N38474,N38475,N38476,
  N38477,N38478,N38479,N38480,N38481,N38482,N38483,N38484,N38485,N38486,N38487,N38488,
  N38489,N38490,N38491,N38492,N38493,N38494,N38495,N38496,N38497,N38498,N38499,
  N38500,N38501,N38502,N38503,N38504,N38505,N38506,N38507,N38508,N38509,N38510,N38511,
  N38512,N38513,N38514,N38515,N38516,N38517,N38518,N38519,N38520,N38521,N38522,
  N38523,N38524,N38525,N38526,N38527,N38528,N38529,N38530,N38531,N38532,N38533,
  N38534,N38535,N38536,N38537,N38538,N38539,N38540,N38541,N38542,N38543,N38544,N38545,
  N38546,N38547,N38548,N38549,N38550,N38551,N38552,N38553,N38554,N38555,N38556,
  N38557,N38558,N38559,N38560,N38561,N38562,N38563,N38564,N38565,N38566,N38567,N38568,
  N38569,N38570,N38571,N38572,N38573,N38574,N38575,N38576,N38577,N38578,N38579,
  N38580,N38581,N38582,N38583,N38584,N38585,N38586,N38587,N38588,N38589,N38590,N38591,
  N38592,N38593,N38594,N38595,N38596,N38597,N38598,N38599,N38600,N38601,N38602,
  N38603,N38604,N38605,N38606,N38607,N38608,N38609,N38610,N38611,N38612,N38613,
  N38614,N38615,N38616,N38617,N38618,N38619,N38620,N38621,N38622,N38623,N38624,N38625,
  N38626,N38627,N38628,N38629,N38630,N38631,N38632,N38633,N38634,N38635,N38636,
  N38637,N38638,N38639,N38640,N38641,N38642,N38643,N38644,N38645,N38646,N38647,N38648,
  N38649,N38650,N38651,N38652,N38653,N38654,N38655,N38656,N38657,N38658,N38659,
  N38660,N38661,N38662,N38663,N38664,N38665,N38666,N38667,N38668,N38669,N38670,N38671,
  N38672,N38673,N38674,N38676,N38677,N38678,N38679,N38680,N38681,N38682,N38683,
  N38684,N38685,N38686,N38687,N38688,N38689,N38690,N38691,N38692,N38693,N38694,
  N38695,N38696,N38697,N38698,N38699,N38700,N38701,N38702,N38703,N38704,N38705,N38706,
  N38707,N38708,N38709,N38710,N38711,N38712,N38713,N38714,N38715,N38716,N38717,
  N38718,N38719,N38720,N38721,N38722,N38723,N38724,N38725,N38726,N38727,N38728,N38729,
  N38730,N38731,N38732,N38733,N38734,N38735,N38736,N38737,N38738,N38739,N38740,
  N38741,N38742,N38743,N38744,N38745,N38746,N38747,N38748,N38749,N38750,N38751,N38752,
  N38753,N38754,N38755,N38756,N38757,N38758,N38759,N38760,N38761,N38762,N38763,
  N38764,N38765,N38766,N38767,N38768,N38769,N38770,N38771,N38772,N38773,N38774,
  N38775,N38776,N38777,N38778,N38779,N38780,N38781,N38782,N38783,N38784,N38785,N38786,
  N38787,N38788,N38789,N38790,N38791,N38792,N38793,N38794,N38795,N38796,N38797,
  N38798,N38799,N38800,N38801,N38802,N38803,N38804,N38805,N38806,N38807,N38808,N38809,
  N38810,N38811,N38812,N38813,N38814,N38815,N38816,N38817,N38818,N38819,N38820,
  N38821,N38822,N38823,N38824,N38825,N38826,N38827,N38828,N38829,N38830,N38831,N38832,
  N38833,N38834,N38835,N38836,N38837,N38838,N38839,N38840,N38841,N38842,N38843,
  N38844,N38845,N38846,N38847,N38848,N38849,N38850,N38851,N38852,N38853,N38854,
  N38855,N38856,N38857,N38858,N38859,N38860,N38861,N38862,N38863,N38864,N38865,N38866,
  N38867,N38868,N38869,N38870,N38871,N38872,N38873,N38874,N38875,N38876,N38877,
  N38878,N38879,N38880,N38881,N38882,N38883,N38884,N38885,N38886,N38887,N38888,N38889,
  N38890,N38891,N38892,N38893,N38894,N38895,N38896,N38897,N38898,N38899,N38900,
  N38901,N38902,N38903,N38904,N38905,N38906,N38907,N38908,N38909,N38910,N38911,N38912,
  N38913,N38914,N38915,N38916,N38917,N38918,N38919,N38920,N38921,N38922,N38923,
  N38924,N38925,N38926,N38927,N38928,N38929,N38930,N38931,N38932,N38933,N38934,
  N38935,N38936,N38937,N38938,N38939,N38940,N38941,N38942,N38943,N38944,N38945,N38946,
  N38947,N38948,N38949,N38950,N38951,N38952,N38953,N38954,N38955;
  wire [2903:0] mem_n;
  wire [2:0] issue_pointer_n,issue_cnt_n,commit_pointer_n;
  reg [361:0] issue_instr_o;
  reg [2903:0] mem_q;
  reg [2:0] issue_cnt_q,commit_pointer_q;
  assign rd_clobber_fpr_o[0] = 1'b0;
  assign rd_clobber_fpr_o[1] = 1'b0;
  assign rd_clobber_fpr_o[2] = 1'b0;
  assign rd_clobber_fpr_o[3] = 1'b0;
  assign rd_clobber_fpr_o[4] = 1'b0;
  assign rd_clobber_fpr_o[5] = 1'b0;
  assign rd_clobber_fpr_o[6] = 1'b0;
  assign rd_clobber_fpr_o[7] = 1'b0;
  assign rd_clobber_fpr_o[8] = 1'b0;
  assign rd_clobber_fpr_o[9] = 1'b0;
  assign rd_clobber_fpr_o[10] = 1'b0;
  assign rd_clobber_fpr_o[11] = 1'b0;
  assign rd_clobber_fpr_o[12] = 1'b0;
  assign rd_clobber_fpr_o[13] = 1'b0;
  assign rd_clobber_fpr_o[14] = 1'b0;
  assign rd_clobber_fpr_o[15] = 1'b0;
  assign rd_clobber_fpr_o[16] = 1'b0;
  assign rd_clobber_fpr_o[17] = 1'b0;
  assign rd_clobber_fpr_o[18] = 1'b0;
  assign rd_clobber_fpr_o[19] = 1'b0;
  assign rd_clobber_fpr_o[20] = 1'b0;
  assign rd_clobber_fpr_o[21] = 1'b0;
  assign rd_clobber_fpr_o[22] = 1'b0;
  assign rd_clobber_fpr_o[23] = 1'b0;
  assign rd_clobber_fpr_o[24] = 1'b0;
  assign rd_clobber_fpr_o[25] = 1'b0;
  assign rd_clobber_fpr_o[26] = 1'b0;
  assign rd_clobber_fpr_o[27] = 1'b0;
  assign rd_clobber_fpr_o[28] = 1'b0;
  assign rd_clobber_fpr_o[29] = 1'b0;
  assign rd_clobber_fpr_o[30] = 1'b0;
  assign rd_clobber_fpr_o[31] = 1'b0;
  assign rd_clobber_fpr_o[32] = 1'b0;
  assign rd_clobber_fpr_o[33] = 1'b0;
  assign rd_clobber_fpr_o[34] = 1'b0;
  assign rd_clobber_fpr_o[35] = 1'b0;
  assign rd_clobber_fpr_o[36] = 1'b0;
  assign rd_clobber_fpr_o[37] = 1'b0;
  assign rd_clobber_fpr_o[38] = 1'b0;
  assign rd_clobber_fpr_o[39] = 1'b0;
  assign rd_clobber_fpr_o[40] = 1'b0;
  assign rd_clobber_fpr_o[41] = 1'b0;
  assign rd_clobber_fpr_o[42] = 1'b0;
  assign rd_clobber_fpr_o[43] = 1'b0;
  assign rd_clobber_fpr_o[44] = 1'b0;
  assign rd_clobber_fpr_o[45] = 1'b0;
  assign rd_clobber_fpr_o[46] = 1'b0;
  assign rd_clobber_fpr_o[47] = 1'b0;
  assign rd_clobber_fpr_o[48] = 1'b0;
  assign rd_clobber_fpr_o[49] = 1'b0;
  assign rd_clobber_fpr_o[50] = 1'b0;
  assign rd_clobber_fpr_o[51] = 1'b0;
  assign rd_clobber_fpr_o[52] = 1'b0;
  assign rd_clobber_fpr_o[53] = 1'b0;
  assign rd_clobber_fpr_o[54] = 1'b0;
  assign rd_clobber_fpr_o[55] = 1'b0;
  assign rd_clobber_fpr_o[56] = 1'b0;
  assign rd_clobber_fpr_o[57] = 1'b0;
  assign rd_clobber_fpr_o[58] = 1'b0;
  assign rd_clobber_fpr_o[59] = 1'b0;
  assign rd_clobber_fpr_o[60] = 1'b0;
  assign rd_clobber_fpr_o[61] = 1'b0;
  assign rd_clobber_fpr_o[62] = 1'b0;
  assign rd_clobber_fpr_o[63] = 1'b0;
  assign rd_clobber_fpr_o[64] = 1'b0;
  assign rd_clobber_fpr_o[65] = 1'b0;
  assign rd_clobber_fpr_o[66] = 1'b0;
  assign rd_clobber_fpr_o[67] = 1'b0;
  assign rd_clobber_fpr_o[68] = 1'b0;
  assign rd_clobber_fpr_o[69] = 1'b0;
  assign rd_clobber_fpr_o[70] = 1'b0;
  assign rd_clobber_fpr_o[71] = 1'b0;
  assign rd_clobber_fpr_o[72] = 1'b0;
  assign rd_clobber_fpr_o[73] = 1'b0;
  assign rd_clobber_fpr_o[74] = 1'b0;
  assign rd_clobber_fpr_o[75] = 1'b0;
  assign rd_clobber_fpr_o[76] = 1'b0;
  assign rd_clobber_fpr_o[77] = 1'b0;
  assign rd_clobber_fpr_o[78] = 1'b0;
  assign rd_clobber_fpr_o[79] = 1'b0;
  assign rd_clobber_fpr_o[80] = 1'b0;
  assign rd_clobber_fpr_o[81] = 1'b0;
  assign rd_clobber_fpr_o[82] = 1'b0;
  assign rd_clobber_fpr_o[83] = 1'b0;
  assign rd_clobber_fpr_o[84] = 1'b0;
  assign rd_clobber_fpr_o[85] = 1'b0;
  assign rd_clobber_fpr_o[86] = 1'b0;
  assign rd_clobber_fpr_o[87] = 1'b0;
  assign rd_clobber_fpr_o[88] = 1'b0;
  assign rd_clobber_fpr_o[89] = 1'b0;
  assign rd_clobber_fpr_o[90] = 1'b0;
  assign rd_clobber_fpr_o[91] = 1'b0;
  assign rd_clobber_fpr_o[92] = 1'b0;
  assign rd_clobber_fpr_o[93] = 1'b0;
  assign rd_clobber_fpr_o[94] = 1'b0;
  assign rd_clobber_fpr_o[95] = 1'b0;
  assign rd_clobber_fpr_o[96] = 1'b0;
  assign rd_clobber_fpr_o[97] = 1'b0;
  assign rd_clobber_fpr_o[98] = 1'b0;
  assign rd_clobber_fpr_o[99] = 1'b0;
  assign rd_clobber_fpr_o[100] = 1'b0;
  assign rd_clobber_fpr_o[101] = 1'b0;
  assign rd_clobber_fpr_o[102] = 1'b0;
  assign rd_clobber_fpr_o[103] = 1'b0;
  assign rd_clobber_fpr_o[104] = 1'b0;
  assign rd_clobber_fpr_o[105] = 1'b0;
  assign rd_clobber_fpr_o[106] = 1'b0;
  assign rd_clobber_fpr_o[107] = 1'b0;
  assign rd_clobber_fpr_o[108] = 1'b0;
  assign rd_clobber_fpr_o[109] = 1'b0;
  assign rd_clobber_fpr_o[110] = 1'b0;
  assign rd_clobber_fpr_o[111] = 1'b0;
  assign rd_clobber_fpr_o[112] = 1'b0;
  assign rd_clobber_fpr_o[113] = 1'b0;
  assign rd_clobber_fpr_o[114] = 1'b0;
  assign rd_clobber_fpr_o[115] = 1'b0;
  assign rd_clobber_fpr_o[116] = 1'b0;
  assign rd_clobber_fpr_o[117] = 1'b0;
  assign rd_clobber_fpr_o[118] = 1'b0;
  assign rd_clobber_fpr_o[119] = 1'b0;
  assign rd_clobber_fpr_o[120] = 1'b0;
  assign rd_clobber_fpr_o[121] = 1'b0;
  assign rd_clobber_fpr_o[122] = 1'b0;
  assign rd_clobber_fpr_o[123] = 1'b0;
  assign rd_clobber_fpr_o[124] = 1'b0;
  assign rd_clobber_fpr_o[125] = 1'b0;
  assign rd_clobber_fpr_o[126] = 1'b0;
  assign rd_clobber_fpr_o[127] = 1'b0;
  assign rd_clobber_fpr_o[128] = 1'b0;
  assign rd_clobber_fpr_o[129] = 1'b0;
  assign rd_clobber_fpr_o[130] = 1'b0;
  assign rd_clobber_fpr_o[131] = 1'b0;
  assign rd_clobber_fpr_o[132] = 1'b0;
  assign rd_clobber_fpr_o[133] = 1'b0;
  assign rd_clobber_fpr_o[134] = 1'b0;
  assign rd_clobber_fpr_o[135] = 1'b0;
  assign rd_clobber_fpr_o[136] = 1'b0;
  assign rd_clobber_fpr_o[137] = 1'b0;
  assign rd_clobber_fpr_o[138] = 1'b0;
  assign rd_clobber_fpr_o[139] = 1'b0;
  assign rd_clobber_fpr_o[140] = 1'b0;
  assign rd_clobber_fpr_o[141] = 1'b0;
  assign rd_clobber_fpr_o[142] = 1'b0;
  assign rd_clobber_fpr_o[143] = 1'b0;
  assign rd_clobber_fpr_o[144] = 1'b0;
  assign rd_clobber_fpr_o[145] = 1'b0;
  assign rd_clobber_fpr_o[146] = 1'b0;
  assign rd_clobber_fpr_o[147] = 1'b0;
  assign rd_clobber_fpr_o[148] = 1'b0;
  assign rd_clobber_fpr_o[149] = 1'b0;
  assign rd_clobber_fpr_o[150] = 1'b0;
  assign rd_clobber_fpr_o[151] = 1'b0;
  assign rd_clobber_fpr_o[152] = 1'b0;
  assign rd_clobber_fpr_o[153] = 1'b0;
  assign rd_clobber_fpr_o[154] = 1'b0;
  assign rd_clobber_fpr_o[155] = 1'b0;
  assign rd_clobber_fpr_o[156] = 1'b0;
  assign rd_clobber_fpr_o[157] = 1'b0;
  assign rd_clobber_fpr_o[158] = 1'b0;
  assign rd_clobber_fpr_o[159] = 1'b0;
  assign rd_clobber_fpr_o[160] = 1'b0;
  assign rd_clobber_fpr_o[161] = 1'b0;
  assign rd_clobber_fpr_o[162] = 1'b0;
  assign rd_clobber_fpr_o[163] = 1'b0;
  assign rd_clobber_fpr_o[164] = 1'b0;
  assign rd_clobber_fpr_o[165] = 1'b0;
  assign rd_clobber_fpr_o[166] = 1'b0;
  assign rd_clobber_fpr_o[167] = 1'b0;
  assign rd_clobber_fpr_o[168] = 1'b0;
  assign rd_clobber_fpr_o[169] = 1'b0;
  assign rd_clobber_fpr_o[170] = 1'b0;
  assign rd_clobber_fpr_o[171] = 1'b0;
  assign rd_clobber_fpr_o[172] = 1'b0;
  assign rd_clobber_fpr_o[173] = 1'b0;
  assign rd_clobber_fpr_o[174] = 1'b0;
  assign rd_clobber_fpr_o[175] = 1'b0;
  assign rd_clobber_fpr_o[176] = 1'b0;
  assign rd_clobber_fpr_o[177] = 1'b0;
  assign rd_clobber_fpr_o[178] = 1'b0;
  assign rd_clobber_fpr_o[179] = 1'b0;
  assign rd_clobber_fpr_o[180] = 1'b0;
  assign rd_clobber_fpr_o[181] = 1'b0;
  assign rd_clobber_fpr_o[182] = 1'b0;
  assign rd_clobber_fpr_o[183] = 1'b0;
  assign rd_clobber_fpr_o[184] = 1'b0;
  assign rd_clobber_fpr_o[185] = 1'b0;
  assign rd_clobber_fpr_o[186] = 1'b0;
  assign rd_clobber_fpr_o[187] = 1'b0;
  assign rd_clobber_fpr_o[188] = 1'b0;
  assign rd_clobber_fpr_o[189] = 1'b0;
  assign rd_clobber_fpr_o[190] = 1'b0;
  assign rd_clobber_fpr_o[191] = 1'b0;
  assign rd_clobber_fpr_o[192] = 1'b0;
  assign rd_clobber_fpr_o[193] = 1'b0;
  assign rd_clobber_fpr_o[194] = 1'b0;
  assign rd_clobber_fpr_o[195] = 1'b0;
  assign rd_clobber_fpr_o[196] = 1'b0;
  assign rd_clobber_fpr_o[197] = 1'b0;
  assign rd_clobber_fpr_o[198] = 1'b0;
  assign rd_clobber_fpr_o[199] = 1'b0;
  assign rd_clobber_fpr_o[200] = 1'b0;
  assign rd_clobber_fpr_o[201] = 1'b0;
  assign rd_clobber_fpr_o[202] = 1'b0;
  assign rd_clobber_fpr_o[203] = 1'b0;
  assign rd_clobber_fpr_o[204] = 1'b0;
  assign rd_clobber_fpr_o[205] = 1'b0;
  assign rd_clobber_fpr_o[206] = 1'b0;
  assign rd_clobber_fpr_o[207] = 1'b0;
  assign rd_clobber_fpr_o[208] = 1'b0;
  assign rd_clobber_fpr_o[209] = 1'b0;
  assign rd_clobber_fpr_o[210] = 1'b0;
  assign rd_clobber_fpr_o[211] = 1'b0;
  assign rd_clobber_fpr_o[212] = 1'b0;
  assign rd_clobber_fpr_o[213] = 1'b0;
  assign rd_clobber_fpr_o[214] = 1'b0;
  assign rd_clobber_fpr_o[215] = 1'b0;
  assign rd_clobber_fpr_o[216] = 1'b0;
  assign rd_clobber_fpr_o[217] = 1'b0;
  assign rd_clobber_fpr_o[218] = 1'b0;
  assign rd_clobber_fpr_o[219] = 1'b0;
  assign rd_clobber_fpr_o[220] = 1'b0;
  assign rd_clobber_fpr_o[221] = 1'b0;
  assign rd_clobber_fpr_o[222] = 1'b0;
  assign rd_clobber_fpr_o[223] = 1'b0;
  assign rd_clobber_fpr_o[224] = 1'b0;
  assign rd_clobber_fpr_o[225] = 1'b0;
  assign rd_clobber_fpr_o[226] = 1'b0;
  assign rd_clobber_fpr_o[227] = 1'b0;
  assign rd_clobber_fpr_o[228] = 1'b0;
  assign rd_clobber_fpr_o[229] = 1'b0;
  assign rd_clobber_fpr_o[230] = 1'b0;
  assign rd_clobber_fpr_o[231] = 1'b0;
  assign rd_clobber_fpr_o[232] = 1'b0;
  assign rd_clobber_fpr_o[233] = 1'b0;
  assign rd_clobber_fpr_o[234] = 1'b0;
  assign rd_clobber_fpr_o[235] = 1'b0;
  assign rd_clobber_fpr_o[236] = 1'b0;
  assign rd_clobber_fpr_o[237] = 1'b0;
  assign rd_clobber_fpr_o[238] = 1'b0;
  assign rd_clobber_fpr_o[239] = 1'b0;
  assign rd_clobber_fpr_o[240] = 1'b0;
  assign rd_clobber_fpr_o[241] = 1'b0;
  assign rd_clobber_fpr_o[242] = 1'b0;
  assign rd_clobber_fpr_o[243] = 1'b0;
  assign rd_clobber_fpr_o[244] = 1'b0;
  assign rd_clobber_fpr_o[245] = 1'b0;
  assign rd_clobber_fpr_o[246] = 1'b0;
  assign rd_clobber_fpr_o[247] = 1'b0;
  assign rd_clobber_fpr_o[248] = 1'b0;
  assign rd_clobber_fpr_o[249] = 1'b0;
  assign rd_clobber_fpr_o[250] = 1'b0;
  assign rd_clobber_fpr_o[251] = 1'b0;
  assign rd_clobber_fpr_o[252] = 1'b0;
  assign rd_clobber_fpr_o[253] = 1'b0;
  assign rd_clobber_fpr_o[254] = 1'b0;
  assign rd_clobber_fpr_o[255] = 1'b0;
  assign rd_clobber_fpr_o[256] = 1'b0;
  assign rd_clobber_fpr_o[257] = 1'b0;
  assign rd_clobber_fpr_o[258] = 1'b0;
  assign rd_clobber_fpr_o[259] = 1'b0;
  assign rd_clobber_gpr_o[0] = 1'b0;
  assign rd_clobber_gpr_o[1] = 1'b0;
  assign rd_clobber_gpr_o[2] = 1'b0;
  assign rd_clobber_gpr_o[3] = 1'b0;
  assign rd_clobber_gpr_o[256] = 1'b0;
  assign rd_clobber_gpr_o[257] = 1'b0;
  assign rd_clobber_gpr_o[258] = 1'b0;
  assign rd_clobber_gpr_o[259] = 1'b0;
  assign issue_instr_o[361] = decoded_instr_i[361];
  assign issue_instr_o[360] = decoded_instr_i[360];
  assign issue_instr_o[359] = decoded_instr_i[359];
  assign issue_instr_o[358] = decoded_instr_i[358];
  assign issue_instr_o[357] = decoded_instr_i[357];
  assign issue_instr_o[356] = decoded_instr_i[356];
  assign issue_instr_o[355] = decoded_instr_i[355];
  assign issue_instr_o[354] = decoded_instr_i[354];
  assign issue_instr_o[353] = decoded_instr_i[353];
  assign issue_instr_o[352] = decoded_instr_i[352];
  assign issue_instr_o[351] = decoded_instr_i[351];
  assign issue_instr_o[350] = decoded_instr_i[350];
  assign issue_instr_o[349] = decoded_instr_i[349];
  assign issue_instr_o[348] = decoded_instr_i[348];
  assign issue_instr_o[347] = decoded_instr_i[347];
  assign issue_instr_o[346] = decoded_instr_i[346];
  assign issue_instr_o[345] = decoded_instr_i[345];
  assign issue_instr_o[344] = decoded_instr_i[344];
  assign issue_instr_o[343] = decoded_instr_i[343];
  assign issue_instr_o[342] = decoded_instr_i[342];
  assign issue_instr_o[341] = decoded_instr_i[341];
  assign issue_instr_o[340] = decoded_instr_i[340];
  assign issue_instr_o[339] = decoded_instr_i[339];
  assign issue_instr_o[338] = decoded_instr_i[338];
  assign issue_instr_o[337] = decoded_instr_i[337];
  assign issue_instr_o[336] = decoded_instr_i[336];
  assign issue_instr_o[335] = decoded_instr_i[335];
  assign issue_instr_o[334] = decoded_instr_i[334];
  assign issue_instr_o[333] = decoded_instr_i[333];
  assign issue_instr_o[332] = decoded_instr_i[332];
  assign issue_instr_o[331] = decoded_instr_i[331];
  assign issue_instr_o[330] = decoded_instr_i[330];
  assign issue_instr_o[329] = decoded_instr_i[329];
  assign issue_instr_o[328] = decoded_instr_i[328];
  assign issue_instr_o[327] = decoded_instr_i[327];
  assign issue_instr_o[326] = decoded_instr_i[326];
  assign issue_instr_o[325] = decoded_instr_i[325];
  assign issue_instr_o[324] = decoded_instr_i[324];
  assign issue_instr_o[323] = decoded_instr_i[323];
  assign issue_instr_o[322] = decoded_instr_i[322];
  assign issue_instr_o[321] = decoded_instr_i[321];
  assign issue_instr_o[320] = decoded_instr_i[320];
  assign issue_instr_o[319] = decoded_instr_i[319];
  assign issue_instr_o[318] = decoded_instr_i[318];
  assign issue_instr_o[317] = decoded_instr_i[317];
  assign issue_instr_o[316] = decoded_instr_i[316];
  assign issue_instr_o[315] = decoded_instr_i[315];
  assign issue_instr_o[314] = decoded_instr_i[314];
  assign issue_instr_o[313] = decoded_instr_i[313];
  assign issue_instr_o[312] = decoded_instr_i[312];
  assign issue_instr_o[311] = decoded_instr_i[311];
  assign issue_instr_o[310] = decoded_instr_i[310];
  assign issue_instr_o[309] = decoded_instr_i[309];
  assign issue_instr_o[308] = decoded_instr_i[308];
  assign issue_instr_o[307] = decoded_instr_i[307];
  assign issue_instr_o[306] = decoded_instr_i[306];
  assign issue_instr_o[305] = decoded_instr_i[305];
  assign issue_instr_o[304] = decoded_instr_i[304];
  assign issue_instr_o[303] = decoded_instr_i[303];
  assign issue_instr_o[302] = decoded_instr_i[302];
  assign issue_instr_o[301] = decoded_instr_i[301];
  assign issue_instr_o[300] = decoded_instr_i[300];
  assign issue_instr_o[299] = decoded_instr_i[299];
  assign issue_instr_o[298] = decoded_instr_i[298];
  assign issue_instr_o[294] = decoded_instr_i[294];
  assign issue_instr_o[293] = decoded_instr_i[293];
  assign issue_instr_o[292] = decoded_instr_i[292];
  assign issue_instr_o[291] = decoded_instr_i[291];
  assign issue_instr_o[290] = decoded_instr_i[290];
  assign issue_instr_o[289] = decoded_instr_i[289];
  assign issue_instr_o[288] = decoded_instr_i[288];
  assign issue_instr_o[287] = decoded_instr_i[287];
  assign issue_instr_o[286] = decoded_instr_i[286];
  assign issue_instr_o[285] = decoded_instr_i[285];
  assign issue_instr_o[284] = decoded_instr_i[284];
  assign issue_instr_o[283] = decoded_instr_i[283];
  assign issue_instr_o[282] = decoded_instr_i[282];
  assign issue_instr_o[281] = decoded_instr_i[281];
  assign issue_instr_o[280] = decoded_instr_i[280];
  assign issue_instr_o[279] = decoded_instr_i[279];
  assign issue_instr_o[278] = decoded_instr_i[278];
  assign issue_instr_o[277] = decoded_instr_i[277];
  assign issue_instr_o[276] = decoded_instr_i[276];
  assign issue_instr_o[275] = decoded_instr_i[275];
  assign issue_instr_o[274] = decoded_instr_i[274];
  assign issue_instr_o[273] = decoded_instr_i[273];
  assign issue_instr_o[272] = decoded_instr_i[272];
  assign issue_instr_o[271] = decoded_instr_i[271];
  assign issue_instr_o[270] = decoded_instr_i[270];
  assign issue_instr_o[269] = decoded_instr_i[269];
  assign issue_instr_o[268] = decoded_instr_i[268];
  assign issue_instr_o[267] = decoded_instr_i[267];
  assign issue_instr_o[266] = decoded_instr_i[266];
  assign issue_instr_o[265] = decoded_instr_i[265];
  assign issue_instr_o[264] = decoded_instr_i[264];
  assign issue_instr_o[263] = decoded_instr_i[263];
  assign issue_instr_o[262] = decoded_instr_i[262];
  assign issue_instr_o[261] = decoded_instr_i[261];
  assign issue_instr_o[260] = decoded_instr_i[260];
  assign issue_instr_o[259] = decoded_instr_i[259];
  assign issue_instr_o[258] = decoded_instr_i[258];
  assign issue_instr_o[257] = decoded_instr_i[257];
  assign issue_instr_o[256] = decoded_instr_i[256];
  assign issue_instr_o[255] = decoded_instr_i[255];
  assign issue_instr_o[254] = decoded_instr_i[254];
  assign issue_instr_o[253] = decoded_instr_i[253];
  assign issue_instr_o[252] = decoded_instr_i[252];
  assign issue_instr_o[251] = decoded_instr_i[251];
  assign issue_instr_o[250] = decoded_instr_i[250];
  assign issue_instr_o[249] = decoded_instr_i[249];
  assign issue_instr_o[248] = decoded_instr_i[248];
  assign issue_instr_o[247] = decoded_instr_i[247];
  assign issue_instr_o[246] = decoded_instr_i[246];
  assign issue_instr_o[245] = decoded_instr_i[245];
  assign issue_instr_o[244] = decoded_instr_i[244];
  assign issue_instr_o[243] = decoded_instr_i[243];
  assign issue_instr_o[242] = decoded_instr_i[242];
  assign issue_instr_o[241] = decoded_instr_i[241];
  assign issue_instr_o[240] = decoded_instr_i[240];
  assign issue_instr_o[239] = decoded_instr_i[239];
  assign issue_instr_o[238] = decoded_instr_i[238];
  assign issue_instr_o[237] = decoded_instr_i[237];
  assign issue_instr_o[236] = decoded_instr_i[236];
  assign issue_instr_o[235] = decoded_instr_i[235];
  assign issue_instr_o[234] = decoded_instr_i[234];
  assign issue_instr_o[233] = decoded_instr_i[233];
  assign issue_instr_o[232] = decoded_instr_i[232];
  assign issue_instr_o[231] = decoded_instr_i[231];
  assign issue_instr_o[230] = decoded_instr_i[230];
  assign issue_instr_o[229] = decoded_instr_i[229];
  assign issue_instr_o[228] = decoded_instr_i[228];
  assign issue_instr_o[227] = decoded_instr_i[227];
  assign issue_instr_o[226] = decoded_instr_i[226];
  assign issue_instr_o[225] = decoded_instr_i[225];
  assign issue_instr_o[224] = decoded_instr_i[224];
  assign issue_instr_o[223] = decoded_instr_i[223];
  assign issue_instr_o[222] = decoded_instr_i[222];
  assign issue_instr_o[221] = decoded_instr_i[221];
  assign issue_instr_o[220] = decoded_instr_i[220];
  assign issue_instr_o[219] = decoded_instr_i[219];
  assign issue_instr_o[218] = decoded_instr_i[218];
  assign issue_instr_o[217] = decoded_instr_i[217];
  assign issue_instr_o[216] = decoded_instr_i[216];
  assign issue_instr_o[215] = decoded_instr_i[215];
  assign issue_instr_o[214] = decoded_instr_i[214];
  assign issue_instr_o[213] = decoded_instr_i[213];
  assign issue_instr_o[212] = decoded_instr_i[212];
  assign issue_instr_o[211] = decoded_instr_i[211];
  assign issue_instr_o[210] = decoded_instr_i[210];
  assign issue_instr_o[209] = decoded_instr_i[209];
  assign issue_instr_o[208] = decoded_instr_i[208];
  assign issue_instr_o[207] = decoded_instr_i[207];
  assign issue_instr_o[206] = decoded_instr_i[206];
  assign issue_instr_o[205] = decoded_instr_i[205];
  assign issue_instr_o[204] = decoded_instr_i[204];
  assign issue_instr_o[203] = decoded_instr_i[203];
  assign issue_instr_o[202] = decoded_instr_i[202];
  assign issue_instr_o[201] = decoded_instr_i[201];
  assign issue_instr_o[200] = decoded_instr_i[200];
  assign issue_instr_o[199] = decoded_instr_i[199];
  assign issue_instr_o[198] = decoded_instr_i[198];
  assign issue_instr_o[197] = decoded_instr_i[197];
  assign issue_instr_o[196] = decoded_instr_i[196];
  assign issue_instr_o[195] = decoded_instr_i[195];
  assign issue_instr_o[194] = decoded_instr_i[194];
  assign issue_instr_o[193] = decoded_instr_i[193];
  assign issue_instr_o[192] = decoded_instr_i[192];
  assign issue_instr_o[191] = decoded_instr_i[191];
  assign issue_instr_o[190] = decoded_instr_i[190];
  assign issue_instr_o[189] = decoded_instr_i[189];
  assign issue_instr_o[188] = decoded_instr_i[188];
  assign issue_instr_o[187] = decoded_instr_i[187];
  assign issue_instr_o[186] = decoded_instr_i[186];
  assign issue_instr_o[185] = decoded_instr_i[185];
  assign issue_instr_o[184] = decoded_instr_i[184];
  assign issue_instr_o[183] = decoded_instr_i[183];
  assign issue_instr_o[182] = decoded_instr_i[182];
  assign issue_instr_o[181] = decoded_instr_i[181];
  assign issue_instr_o[180] = decoded_instr_i[180];
  assign issue_instr_o[179] = decoded_instr_i[179];
  assign issue_instr_o[178] = decoded_instr_i[178];
  assign issue_instr_o[177] = decoded_instr_i[177];
  assign issue_instr_o[176] = decoded_instr_i[176];
  assign issue_instr_o[175] = decoded_instr_i[175];
  assign issue_instr_o[174] = decoded_instr_i[174];
  assign issue_instr_o[173] = decoded_instr_i[173];
  assign issue_instr_o[172] = decoded_instr_i[172];
  assign issue_instr_o[171] = decoded_instr_i[171];
  assign issue_instr_o[170] = decoded_instr_i[170];
  assign issue_instr_o[169] = decoded_instr_i[169];
  assign issue_instr_o[168] = decoded_instr_i[168];
  assign issue_instr_o[167] = decoded_instr_i[167];
  assign issue_instr_o[166] = decoded_instr_i[166];
  assign issue_instr_o[165] = decoded_instr_i[165];
  assign issue_instr_o[164] = decoded_instr_i[164];
  assign issue_instr_o[163] = decoded_instr_i[163];
  assign issue_instr_o[162] = decoded_instr_i[162];
  assign issue_instr_o[161] = decoded_instr_i[161];
  assign issue_instr_o[160] = decoded_instr_i[160];
  assign issue_instr_o[159] = decoded_instr_i[159];
  assign issue_instr_o[158] = decoded_instr_i[158];
  assign issue_instr_o[157] = decoded_instr_i[157];
  assign issue_instr_o[156] = decoded_instr_i[156];
  assign issue_instr_o[155] = decoded_instr_i[155];
  assign issue_instr_o[154] = decoded_instr_i[154];
  assign issue_instr_o[153] = decoded_instr_i[153];
  assign issue_instr_o[152] = decoded_instr_i[152];
  assign issue_instr_o[151] = decoded_instr_i[151];
  assign issue_instr_o[150] = decoded_instr_i[150];
  assign issue_instr_o[149] = decoded_instr_i[149];
  assign issue_instr_o[148] = decoded_instr_i[148];
  assign issue_instr_o[147] = decoded_instr_i[147];
  assign issue_instr_o[146] = decoded_instr_i[146];
  assign issue_instr_o[145] = decoded_instr_i[145];
  assign issue_instr_o[144] = decoded_instr_i[144];
  assign issue_instr_o[143] = decoded_instr_i[143];
  assign issue_instr_o[142] = decoded_instr_i[142];
  assign issue_instr_o[141] = decoded_instr_i[141];
  assign issue_instr_o[140] = decoded_instr_i[140];
  assign issue_instr_o[139] = decoded_instr_i[139];
  assign issue_instr_o[138] = decoded_instr_i[138];
  assign issue_instr_o[137] = decoded_instr_i[137];
  assign issue_instr_o[136] = decoded_instr_i[136];
  assign issue_instr_o[135] = decoded_instr_i[135];
  assign issue_instr_o[134] = decoded_instr_i[134];
  assign issue_instr_o[133] = decoded_instr_i[133];
  assign issue_instr_o[132] = decoded_instr_i[132];
  assign issue_instr_o[131] = decoded_instr_i[131];
  assign issue_instr_o[130] = decoded_instr_i[130];
  assign issue_instr_o[129] = decoded_instr_i[129];
  assign issue_instr_o[128] = decoded_instr_i[128];
  assign issue_instr_o[127] = decoded_instr_i[127];
  assign issue_instr_o[126] = decoded_instr_i[126];
  assign issue_instr_o[125] = decoded_instr_i[125];
  assign issue_instr_o[124] = decoded_instr_i[124];
  assign issue_instr_o[123] = decoded_instr_i[123];
  assign issue_instr_o[122] = decoded_instr_i[122];
  assign issue_instr_o[121] = decoded_instr_i[121];
  assign issue_instr_o[120] = decoded_instr_i[120];
  assign issue_instr_o[119] = decoded_instr_i[119];
  assign issue_instr_o[118] = decoded_instr_i[118];
  assign issue_instr_o[117] = decoded_instr_i[117];
  assign issue_instr_o[116] = decoded_instr_i[116];
  assign issue_instr_o[115] = decoded_instr_i[115];
  assign issue_instr_o[114] = decoded_instr_i[114];
  assign issue_instr_o[113] = decoded_instr_i[113];
  assign issue_instr_o[112] = decoded_instr_i[112];
  assign issue_instr_o[111] = decoded_instr_i[111];
  assign issue_instr_o[110] = decoded_instr_i[110];
  assign issue_instr_o[109] = decoded_instr_i[109];
  assign issue_instr_o[108] = decoded_instr_i[108];
  assign issue_instr_o[107] = decoded_instr_i[107];
  assign issue_instr_o[106] = decoded_instr_i[106];
  assign issue_instr_o[105] = decoded_instr_i[105];
  assign issue_instr_o[104] = decoded_instr_i[104];
  assign issue_instr_o[103] = decoded_instr_i[103];
  assign issue_instr_o[102] = decoded_instr_i[102];
  assign issue_instr_o[101] = decoded_instr_i[101];
  assign issue_instr_o[100] = decoded_instr_i[100];
  assign issue_instr_o[99] = decoded_instr_i[99];
  assign issue_instr_o[98] = decoded_instr_i[98];
  assign issue_instr_o[97] = decoded_instr_i[97];
  assign issue_instr_o[96] = decoded_instr_i[96];
  assign issue_instr_o[95] = decoded_instr_i[95];
  assign issue_instr_o[94] = decoded_instr_i[94];
  assign issue_instr_o[93] = decoded_instr_i[93];
  assign issue_instr_o[92] = decoded_instr_i[92];
  assign issue_instr_o[91] = decoded_instr_i[91];
  assign issue_instr_o[90] = decoded_instr_i[90];
  assign issue_instr_o[89] = decoded_instr_i[89];
  assign issue_instr_o[88] = decoded_instr_i[88];
  assign issue_instr_o[87] = decoded_instr_i[87];
  assign issue_instr_o[86] = decoded_instr_i[86];
  assign issue_instr_o[85] = decoded_instr_i[85];
  assign issue_instr_o[84] = decoded_instr_i[84];
  assign issue_instr_o[83] = decoded_instr_i[83];
  assign issue_instr_o[82] = decoded_instr_i[82];
  assign issue_instr_o[81] = decoded_instr_i[81];
  assign issue_instr_o[80] = decoded_instr_i[80];
  assign issue_instr_o[79] = decoded_instr_i[79];
  assign issue_instr_o[78] = decoded_instr_i[78];
  assign issue_instr_o[77] = decoded_instr_i[77];
  assign issue_instr_o[76] = decoded_instr_i[76];
  assign issue_instr_o[75] = decoded_instr_i[75];
  assign issue_instr_o[74] = decoded_instr_i[74];
  assign issue_instr_o[73] = decoded_instr_i[73];
  assign issue_instr_o[72] = decoded_instr_i[72];
  assign issue_instr_o[71] = decoded_instr_i[71];
  assign issue_instr_o[70] = decoded_instr_i[70];
  assign issue_instr_o[69] = decoded_instr_i[69];
  assign issue_instr_o[68] = decoded_instr_i[68];
  assign issue_instr_o[67] = decoded_instr_i[67];
  assign issue_instr_o[66] = decoded_instr_i[66];
  assign issue_instr_o[65] = decoded_instr_i[65];
  assign issue_instr_o[64] = decoded_instr_i[64];
  assign issue_instr_o[63] = decoded_instr_i[63];
  assign issue_instr_o[62] = decoded_instr_i[62];
  assign issue_instr_o[61] = decoded_instr_i[61];
  assign issue_instr_o[60] = decoded_instr_i[60];
  assign issue_instr_o[59] = decoded_instr_i[59];
  assign issue_instr_o[58] = decoded_instr_i[58];
  assign issue_instr_o[57] = decoded_instr_i[57];
  assign issue_instr_o[56] = decoded_instr_i[56];
  assign issue_instr_o[55] = decoded_instr_i[55];
  assign issue_instr_o[54] = decoded_instr_i[54];
  assign issue_instr_o[53] = decoded_instr_i[53];
  assign issue_instr_o[52] = decoded_instr_i[52];
  assign issue_instr_o[51] = decoded_instr_i[51];
  assign issue_instr_o[50] = decoded_instr_i[50];
  assign issue_instr_o[49] = decoded_instr_i[49];
  assign issue_instr_o[48] = decoded_instr_i[48];
  assign issue_instr_o[47] = decoded_instr_i[47];
  assign issue_instr_o[46] = decoded_instr_i[46];
  assign issue_instr_o[45] = decoded_instr_i[45];
  assign issue_instr_o[44] = decoded_instr_i[44];
  assign issue_instr_o[43] = decoded_instr_i[43];
  assign issue_instr_o[42] = decoded_instr_i[42];
  assign issue_instr_o[41] = decoded_instr_i[41];
  assign issue_instr_o[40] = decoded_instr_i[40];
  assign issue_instr_o[39] = decoded_instr_i[39];
  assign issue_instr_o[38] = decoded_instr_i[38];
  assign issue_instr_o[37] = decoded_instr_i[37];
  assign issue_instr_o[36] = decoded_instr_i[36];
  assign issue_instr_o[35] = decoded_instr_i[35];
  assign issue_instr_o[34] = decoded_instr_i[34];
  assign issue_instr_o[33] = decoded_instr_i[33];
  assign issue_instr_o[32] = decoded_instr_i[32];
  assign issue_instr_o[31] = decoded_instr_i[31];
  assign issue_instr_o[30] = decoded_instr_i[30];
  assign issue_instr_o[29] = decoded_instr_i[29];
  assign issue_instr_o[28] = decoded_instr_i[28];
  assign issue_instr_o[27] = decoded_instr_i[27];
  assign issue_instr_o[26] = decoded_instr_i[26];
  assign issue_instr_o[25] = decoded_instr_i[25];
  assign issue_instr_o[24] = decoded_instr_i[24];
  assign issue_instr_o[23] = decoded_instr_i[23];
  assign issue_instr_o[22] = decoded_instr_i[22];
  assign issue_instr_o[21] = decoded_instr_i[21];
  assign issue_instr_o[20] = decoded_instr_i[20];
  assign issue_instr_o[19] = decoded_instr_i[19];
  assign issue_instr_o[18] = decoded_instr_i[18];
  assign issue_instr_o[17] = decoded_instr_i[17];
  assign issue_instr_o[16] = decoded_instr_i[16];
  assign issue_instr_o[15] = decoded_instr_i[15];
  assign issue_instr_o[14] = decoded_instr_i[14];
  assign issue_instr_o[13] = decoded_instr_i[13];
  assign issue_instr_o[12] = decoded_instr_i[12];
  assign issue_instr_o[11] = decoded_instr_i[11];
  assign issue_instr_o[10] = decoded_instr_i[10];
  assign issue_instr_o[9] = decoded_instr_i[9];
  assign issue_instr_o[8] = decoded_instr_i[8];
  assign issue_instr_o[7] = decoded_instr_i[7];
  assign issue_instr_o[6] = decoded_instr_i[6];
  assign issue_instr_o[5] = decoded_instr_i[5];
  assign issue_instr_o[4] = decoded_instr_i[4];
  assign issue_instr_o[3] = decoded_instr_i[3];
  assign issue_instr_o[2] = decoded_instr_i[2];
  assign issue_instr_o[1] = decoded_instr_i[1];
  assign issue_instr_o[0] = decoded_instr_i[0];
  assign commit_instr_o[361] = (N856)? mem_q[361] : 
                               (N858)? mem_q[724] : 
                               (N860)? mem_q[1087] : 
                               (N862)? mem_q[1450] : 
                               (N857)? mem_q[1813] : 
                               (N859)? mem_q[2176] : 
                               (N861)? mem_q[2539] : 
                               (N863)? mem_q[2902] : 1'b0;
  assign commit_instr_o[360] = (N856)? mem_q[360] : 
                               (N858)? mem_q[723] : 
                               (N860)? mem_q[1086] : 
                               (N862)? mem_q[1449] : 
                               (N857)? mem_q[1812] : 
                               (N859)? mem_q[2175] : 
                               (N861)? mem_q[2538] : 
                               (N863)? mem_q[2901] : 1'b0;
  assign commit_instr_o[359] = (N856)? mem_q[359] : 
                               (N858)? mem_q[722] : 
                               (N860)? mem_q[1085] : 
                               (N862)? mem_q[1448] : 
                               (N857)? mem_q[1811] : 
                               (N859)? mem_q[2174] : 
                               (N861)? mem_q[2537] : 
                               (N863)? mem_q[2900] : 1'b0;
  assign commit_instr_o[358] = (N856)? mem_q[358] : 
                               (N858)? mem_q[721] : 
                               (N860)? mem_q[1084] : 
                               (N862)? mem_q[1447] : 
                               (N857)? mem_q[1810] : 
                               (N859)? mem_q[2173] : 
                               (N861)? mem_q[2536] : 
                               (N863)? mem_q[2899] : 1'b0;
  assign commit_instr_o[357] = (N856)? mem_q[357] : 
                               (N858)? mem_q[720] : 
                               (N860)? mem_q[1083] : 
                               (N862)? mem_q[1446] : 
                               (N857)? mem_q[1809] : 
                               (N859)? mem_q[2172] : 
                               (N861)? mem_q[2535] : 
                               (N863)? mem_q[2898] : 1'b0;
  assign commit_instr_o[356] = (N856)? mem_q[356] : 
                               (N858)? mem_q[719] : 
                               (N860)? mem_q[1082] : 
                               (N862)? mem_q[1445] : 
                               (N857)? mem_q[1808] : 
                               (N859)? mem_q[2171] : 
                               (N861)? mem_q[2534] : 
                               (N863)? mem_q[2897] : 1'b0;
  assign commit_instr_o[355] = (N856)? mem_q[355] : 
                               (N858)? mem_q[718] : 
                               (N860)? mem_q[1081] : 
                               (N862)? mem_q[1444] : 
                               (N857)? mem_q[1807] : 
                               (N859)? mem_q[2170] : 
                               (N861)? mem_q[2533] : 
                               (N863)? mem_q[2896] : 1'b0;
  assign commit_instr_o[354] = (N856)? mem_q[354] : 
                               (N858)? mem_q[717] : 
                               (N860)? mem_q[1080] : 
                               (N862)? mem_q[1443] : 
                               (N857)? mem_q[1806] : 
                               (N859)? mem_q[2169] : 
                               (N861)? mem_q[2532] : 
                               (N863)? mem_q[2895] : 1'b0;
  assign commit_instr_o[353] = (N856)? mem_q[353] : 
                               (N858)? mem_q[716] : 
                               (N860)? mem_q[1079] : 
                               (N862)? mem_q[1442] : 
                               (N857)? mem_q[1805] : 
                               (N859)? mem_q[2168] : 
                               (N861)? mem_q[2531] : 
                               (N863)? mem_q[2894] : 1'b0;
  assign commit_instr_o[352] = (N856)? mem_q[352] : 
                               (N858)? mem_q[715] : 
                               (N860)? mem_q[1078] : 
                               (N862)? mem_q[1441] : 
                               (N857)? mem_q[1804] : 
                               (N859)? mem_q[2167] : 
                               (N861)? mem_q[2530] : 
                               (N863)? mem_q[2893] : 1'b0;
  assign commit_instr_o[351] = (N856)? mem_q[351] : 
                               (N858)? mem_q[714] : 
                               (N860)? mem_q[1077] : 
                               (N862)? mem_q[1440] : 
                               (N857)? mem_q[1803] : 
                               (N859)? mem_q[2166] : 
                               (N861)? mem_q[2529] : 
                               (N863)? mem_q[2892] : 1'b0;
  assign commit_instr_o[350] = (N856)? mem_q[350] : 
                               (N858)? mem_q[713] : 
                               (N860)? mem_q[1076] : 
                               (N862)? mem_q[1439] : 
                               (N857)? mem_q[1802] : 
                               (N859)? mem_q[2165] : 
                               (N861)? mem_q[2528] : 
                               (N863)? mem_q[2891] : 1'b0;
  assign commit_instr_o[349] = (N856)? mem_q[349] : 
                               (N858)? mem_q[712] : 
                               (N860)? mem_q[1075] : 
                               (N862)? mem_q[1438] : 
                               (N857)? mem_q[1801] : 
                               (N859)? mem_q[2164] : 
                               (N861)? mem_q[2527] : 
                               (N863)? mem_q[2890] : 1'b0;
  assign commit_instr_o[348] = (N856)? mem_q[348] : 
                               (N858)? mem_q[711] : 
                               (N860)? mem_q[1074] : 
                               (N862)? mem_q[1437] : 
                               (N857)? mem_q[1800] : 
                               (N859)? mem_q[2163] : 
                               (N861)? mem_q[2526] : 
                               (N863)? mem_q[2889] : 1'b0;
  assign commit_instr_o[347] = (N856)? mem_q[347] : 
                               (N858)? mem_q[710] : 
                               (N860)? mem_q[1073] : 
                               (N862)? mem_q[1436] : 
                               (N857)? mem_q[1799] : 
                               (N859)? mem_q[2162] : 
                               (N861)? mem_q[2525] : 
                               (N863)? mem_q[2888] : 1'b0;
  assign commit_instr_o[346] = (N856)? mem_q[346] : 
                               (N858)? mem_q[709] : 
                               (N860)? mem_q[1072] : 
                               (N862)? mem_q[1435] : 
                               (N857)? mem_q[1798] : 
                               (N859)? mem_q[2161] : 
                               (N861)? mem_q[2524] : 
                               (N863)? mem_q[2887] : 1'b0;
  assign commit_instr_o[345] = (N856)? mem_q[345] : 
                               (N858)? mem_q[708] : 
                               (N860)? mem_q[1071] : 
                               (N862)? mem_q[1434] : 
                               (N857)? mem_q[1797] : 
                               (N859)? mem_q[2160] : 
                               (N861)? mem_q[2523] : 
                               (N863)? mem_q[2886] : 1'b0;
  assign commit_instr_o[344] = (N856)? mem_q[344] : 
                               (N858)? mem_q[707] : 
                               (N860)? mem_q[1070] : 
                               (N862)? mem_q[1433] : 
                               (N857)? mem_q[1796] : 
                               (N859)? mem_q[2159] : 
                               (N861)? mem_q[2522] : 
                               (N863)? mem_q[2885] : 1'b0;
  assign commit_instr_o[343] = (N856)? mem_q[343] : 
                               (N858)? mem_q[706] : 
                               (N860)? mem_q[1069] : 
                               (N862)? mem_q[1432] : 
                               (N857)? mem_q[1795] : 
                               (N859)? mem_q[2158] : 
                               (N861)? mem_q[2521] : 
                               (N863)? mem_q[2884] : 1'b0;
  assign commit_instr_o[342] = (N856)? mem_q[342] : 
                               (N858)? mem_q[705] : 
                               (N860)? mem_q[1068] : 
                               (N862)? mem_q[1431] : 
                               (N857)? mem_q[1794] : 
                               (N859)? mem_q[2157] : 
                               (N861)? mem_q[2520] : 
                               (N863)? mem_q[2883] : 1'b0;
  assign commit_instr_o[341] = (N856)? mem_q[341] : 
                               (N858)? mem_q[704] : 
                               (N860)? mem_q[1067] : 
                               (N862)? mem_q[1430] : 
                               (N857)? mem_q[1793] : 
                               (N859)? mem_q[2156] : 
                               (N861)? mem_q[2519] : 
                               (N863)? mem_q[2882] : 1'b0;
  assign commit_instr_o[340] = (N856)? mem_q[340] : 
                               (N858)? mem_q[703] : 
                               (N860)? mem_q[1066] : 
                               (N862)? mem_q[1429] : 
                               (N857)? mem_q[1792] : 
                               (N859)? mem_q[2155] : 
                               (N861)? mem_q[2518] : 
                               (N863)? mem_q[2881] : 1'b0;
  assign commit_instr_o[339] = (N856)? mem_q[339] : 
                               (N858)? mem_q[702] : 
                               (N860)? mem_q[1065] : 
                               (N862)? mem_q[1428] : 
                               (N857)? mem_q[1791] : 
                               (N859)? mem_q[2154] : 
                               (N861)? mem_q[2517] : 
                               (N863)? mem_q[2880] : 1'b0;
  assign commit_instr_o[338] = (N856)? mem_q[338] : 
                               (N858)? mem_q[701] : 
                               (N860)? mem_q[1064] : 
                               (N862)? mem_q[1427] : 
                               (N857)? mem_q[1790] : 
                               (N859)? mem_q[2153] : 
                               (N861)? mem_q[2516] : 
                               (N863)? mem_q[2879] : 1'b0;
  assign commit_instr_o[337] = (N856)? mem_q[337] : 
                               (N858)? mem_q[700] : 
                               (N860)? mem_q[1063] : 
                               (N862)? mem_q[1426] : 
                               (N857)? mem_q[1789] : 
                               (N859)? mem_q[2152] : 
                               (N861)? mem_q[2515] : 
                               (N863)? mem_q[2878] : 1'b0;
  assign commit_instr_o[336] = (N856)? mem_q[336] : 
                               (N858)? mem_q[699] : 
                               (N860)? mem_q[1062] : 
                               (N862)? mem_q[1425] : 
                               (N857)? mem_q[1788] : 
                               (N859)? mem_q[2151] : 
                               (N861)? mem_q[2514] : 
                               (N863)? mem_q[2877] : 1'b0;
  assign commit_instr_o[335] = (N856)? mem_q[335] : 
                               (N858)? mem_q[698] : 
                               (N860)? mem_q[1061] : 
                               (N862)? mem_q[1424] : 
                               (N857)? mem_q[1787] : 
                               (N859)? mem_q[2150] : 
                               (N861)? mem_q[2513] : 
                               (N863)? mem_q[2876] : 1'b0;
  assign commit_instr_o[334] = (N856)? mem_q[334] : 
                               (N858)? mem_q[697] : 
                               (N860)? mem_q[1060] : 
                               (N862)? mem_q[1423] : 
                               (N857)? mem_q[1786] : 
                               (N859)? mem_q[2149] : 
                               (N861)? mem_q[2512] : 
                               (N863)? mem_q[2875] : 1'b0;
  assign commit_instr_o[333] = (N856)? mem_q[333] : 
                               (N858)? mem_q[696] : 
                               (N860)? mem_q[1059] : 
                               (N862)? mem_q[1422] : 
                               (N857)? mem_q[1785] : 
                               (N859)? mem_q[2148] : 
                               (N861)? mem_q[2511] : 
                               (N863)? mem_q[2874] : 1'b0;
  assign commit_instr_o[332] = (N856)? mem_q[332] : 
                               (N858)? mem_q[695] : 
                               (N860)? mem_q[1058] : 
                               (N862)? mem_q[1421] : 
                               (N857)? mem_q[1784] : 
                               (N859)? mem_q[2147] : 
                               (N861)? mem_q[2510] : 
                               (N863)? mem_q[2873] : 1'b0;
  assign commit_instr_o[331] = (N856)? mem_q[331] : 
                               (N858)? mem_q[694] : 
                               (N860)? mem_q[1057] : 
                               (N862)? mem_q[1420] : 
                               (N857)? mem_q[1783] : 
                               (N859)? mem_q[2146] : 
                               (N861)? mem_q[2509] : 
                               (N863)? mem_q[2872] : 1'b0;
  assign commit_instr_o[330] = (N856)? mem_q[330] : 
                               (N858)? mem_q[693] : 
                               (N860)? mem_q[1056] : 
                               (N862)? mem_q[1419] : 
                               (N857)? mem_q[1782] : 
                               (N859)? mem_q[2145] : 
                               (N861)? mem_q[2508] : 
                               (N863)? mem_q[2871] : 1'b0;
  assign commit_instr_o[329] = (N856)? mem_q[329] : 
                               (N858)? mem_q[692] : 
                               (N860)? mem_q[1055] : 
                               (N862)? mem_q[1418] : 
                               (N857)? mem_q[1781] : 
                               (N859)? mem_q[2144] : 
                               (N861)? mem_q[2507] : 
                               (N863)? mem_q[2870] : 1'b0;
  assign commit_instr_o[328] = (N856)? mem_q[328] : 
                               (N858)? mem_q[691] : 
                               (N860)? mem_q[1054] : 
                               (N862)? mem_q[1417] : 
                               (N857)? mem_q[1780] : 
                               (N859)? mem_q[2143] : 
                               (N861)? mem_q[2506] : 
                               (N863)? mem_q[2869] : 1'b0;
  assign commit_instr_o[327] = (N856)? mem_q[327] : 
                               (N858)? mem_q[690] : 
                               (N860)? mem_q[1053] : 
                               (N862)? mem_q[1416] : 
                               (N857)? mem_q[1779] : 
                               (N859)? mem_q[2142] : 
                               (N861)? mem_q[2505] : 
                               (N863)? mem_q[2868] : 1'b0;
  assign commit_instr_o[326] = (N856)? mem_q[326] : 
                               (N858)? mem_q[689] : 
                               (N860)? mem_q[1052] : 
                               (N862)? mem_q[1415] : 
                               (N857)? mem_q[1778] : 
                               (N859)? mem_q[2141] : 
                               (N861)? mem_q[2504] : 
                               (N863)? mem_q[2867] : 1'b0;
  assign commit_instr_o[325] = (N856)? mem_q[325] : 
                               (N858)? mem_q[688] : 
                               (N860)? mem_q[1051] : 
                               (N862)? mem_q[1414] : 
                               (N857)? mem_q[1777] : 
                               (N859)? mem_q[2140] : 
                               (N861)? mem_q[2503] : 
                               (N863)? mem_q[2866] : 1'b0;
  assign commit_instr_o[324] = (N856)? mem_q[324] : 
                               (N858)? mem_q[687] : 
                               (N860)? mem_q[1050] : 
                               (N862)? mem_q[1413] : 
                               (N857)? mem_q[1776] : 
                               (N859)? mem_q[2139] : 
                               (N861)? mem_q[2502] : 
                               (N863)? mem_q[2865] : 1'b0;
  assign commit_instr_o[323] = (N856)? mem_q[323] : 
                               (N858)? mem_q[686] : 
                               (N860)? mem_q[1049] : 
                               (N862)? mem_q[1412] : 
                               (N857)? mem_q[1775] : 
                               (N859)? mem_q[2138] : 
                               (N861)? mem_q[2501] : 
                               (N863)? mem_q[2864] : 1'b0;
  assign commit_instr_o[322] = (N856)? mem_q[322] : 
                               (N858)? mem_q[685] : 
                               (N860)? mem_q[1048] : 
                               (N862)? mem_q[1411] : 
                               (N857)? mem_q[1774] : 
                               (N859)? mem_q[2137] : 
                               (N861)? mem_q[2500] : 
                               (N863)? mem_q[2863] : 1'b0;
  assign commit_instr_o[321] = (N856)? mem_q[321] : 
                               (N858)? mem_q[684] : 
                               (N860)? mem_q[1047] : 
                               (N862)? mem_q[1410] : 
                               (N857)? mem_q[1773] : 
                               (N859)? mem_q[2136] : 
                               (N861)? mem_q[2499] : 
                               (N863)? mem_q[2862] : 1'b0;
  assign commit_instr_o[320] = (N856)? mem_q[320] : 
                               (N858)? mem_q[683] : 
                               (N860)? mem_q[1046] : 
                               (N862)? mem_q[1409] : 
                               (N857)? mem_q[1772] : 
                               (N859)? mem_q[2135] : 
                               (N861)? mem_q[2498] : 
                               (N863)? mem_q[2861] : 1'b0;
  assign commit_instr_o[319] = (N856)? mem_q[319] : 
                               (N858)? mem_q[682] : 
                               (N860)? mem_q[1045] : 
                               (N862)? mem_q[1408] : 
                               (N857)? mem_q[1771] : 
                               (N859)? mem_q[2134] : 
                               (N861)? mem_q[2497] : 
                               (N863)? mem_q[2860] : 1'b0;
  assign commit_instr_o[318] = (N856)? mem_q[318] : 
                               (N858)? mem_q[681] : 
                               (N860)? mem_q[1044] : 
                               (N862)? mem_q[1407] : 
                               (N857)? mem_q[1770] : 
                               (N859)? mem_q[2133] : 
                               (N861)? mem_q[2496] : 
                               (N863)? mem_q[2859] : 1'b0;
  assign commit_instr_o[317] = (N856)? mem_q[317] : 
                               (N858)? mem_q[680] : 
                               (N860)? mem_q[1043] : 
                               (N862)? mem_q[1406] : 
                               (N857)? mem_q[1769] : 
                               (N859)? mem_q[2132] : 
                               (N861)? mem_q[2495] : 
                               (N863)? mem_q[2858] : 1'b0;
  assign commit_instr_o[316] = (N856)? mem_q[316] : 
                               (N858)? mem_q[679] : 
                               (N860)? mem_q[1042] : 
                               (N862)? mem_q[1405] : 
                               (N857)? mem_q[1768] : 
                               (N859)? mem_q[2131] : 
                               (N861)? mem_q[2494] : 
                               (N863)? mem_q[2857] : 1'b0;
  assign commit_instr_o[315] = (N856)? mem_q[315] : 
                               (N858)? mem_q[678] : 
                               (N860)? mem_q[1041] : 
                               (N862)? mem_q[1404] : 
                               (N857)? mem_q[1767] : 
                               (N859)? mem_q[2130] : 
                               (N861)? mem_q[2493] : 
                               (N863)? mem_q[2856] : 1'b0;
  assign commit_instr_o[314] = (N856)? mem_q[314] : 
                               (N858)? mem_q[677] : 
                               (N860)? mem_q[1040] : 
                               (N862)? mem_q[1403] : 
                               (N857)? mem_q[1766] : 
                               (N859)? mem_q[2129] : 
                               (N861)? mem_q[2492] : 
                               (N863)? mem_q[2855] : 1'b0;
  assign commit_instr_o[313] = (N856)? mem_q[313] : 
                               (N858)? mem_q[676] : 
                               (N860)? mem_q[1039] : 
                               (N862)? mem_q[1402] : 
                               (N857)? mem_q[1765] : 
                               (N859)? mem_q[2128] : 
                               (N861)? mem_q[2491] : 
                               (N863)? mem_q[2854] : 1'b0;
  assign commit_instr_o[312] = (N856)? mem_q[312] : 
                               (N858)? mem_q[675] : 
                               (N860)? mem_q[1038] : 
                               (N862)? mem_q[1401] : 
                               (N857)? mem_q[1764] : 
                               (N859)? mem_q[2127] : 
                               (N861)? mem_q[2490] : 
                               (N863)? mem_q[2853] : 1'b0;
  assign commit_instr_o[311] = (N856)? mem_q[311] : 
                               (N858)? mem_q[674] : 
                               (N860)? mem_q[1037] : 
                               (N862)? mem_q[1400] : 
                               (N857)? mem_q[1763] : 
                               (N859)? mem_q[2126] : 
                               (N861)? mem_q[2489] : 
                               (N863)? mem_q[2852] : 1'b0;
  assign commit_instr_o[310] = (N856)? mem_q[310] : 
                               (N858)? mem_q[673] : 
                               (N860)? mem_q[1036] : 
                               (N862)? mem_q[1399] : 
                               (N857)? mem_q[1762] : 
                               (N859)? mem_q[2125] : 
                               (N861)? mem_q[2488] : 
                               (N863)? mem_q[2851] : 1'b0;
  assign commit_instr_o[309] = (N856)? mem_q[309] : 
                               (N858)? mem_q[672] : 
                               (N860)? mem_q[1035] : 
                               (N862)? mem_q[1398] : 
                               (N857)? mem_q[1761] : 
                               (N859)? mem_q[2124] : 
                               (N861)? mem_q[2487] : 
                               (N863)? mem_q[2850] : 1'b0;
  assign commit_instr_o[308] = (N856)? mem_q[308] : 
                               (N858)? mem_q[671] : 
                               (N860)? mem_q[1034] : 
                               (N862)? mem_q[1397] : 
                               (N857)? mem_q[1760] : 
                               (N859)? mem_q[2123] : 
                               (N861)? mem_q[2486] : 
                               (N863)? mem_q[2849] : 1'b0;
  assign commit_instr_o[307] = (N856)? mem_q[307] : 
                               (N858)? mem_q[670] : 
                               (N860)? mem_q[1033] : 
                               (N862)? mem_q[1396] : 
                               (N857)? mem_q[1759] : 
                               (N859)? mem_q[2122] : 
                               (N861)? mem_q[2485] : 
                               (N863)? mem_q[2848] : 1'b0;
  assign commit_instr_o[306] = (N856)? mem_q[306] : 
                               (N858)? mem_q[669] : 
                               (N860)? mem_q[1032] : 
                               (N862)? mem_q[1395] : 
                               (N857)? mem_q[1758] : 
                               (N859)? mem_q[2121] : 
                               (N861)? mem_q[2484] : 
                               (N863)? mem_q[2847] : 1'b0;
  assign commit_instr_o[305] = (N856)? mem_q[305] : 
                               (N858)? mem_q[668] : 
                               (N860)? mem_q[1031] : 
                               (N862)? mem_q[1394] : 
                               (N857)? mem_q[1757] : 
                               (N859)? mem_q[2120] : 
                               (N861)? mem_q[2483] : 
                               (N863)? mem_q[2846] : 1'b0;
  assign commit_instr_o[304] = (N856)? mem_q[304] : 
                               (N858)? mem_q[667] : 
                               (N860)? mem_q[1030] : 
                               (N862)? mem_q[1393] : 
                               (N857)? mem_q[1756] : 
                               (N859)? mem_q[2119] : 
                               (N861)? mem_q[2482] : 
                               (N863)? mem_q[2845] : 1'b0;
  assign commit_instr_o[303] = (N856)? mem_q[303] : 
                               (N858)? mem_q[666] : 
                               (N860)? mem_q[1029] : 
                               (N862)? mem_q[1392] : 
                               (N857)? mem_q[1755] : 
                               (N859)? mem_q[2118] : 
                               (N861)? mem_q[2481] : 
                               (N863)? mem_q[2844] : 1'b0;
  assign commit_instr_o[302] = (N856)? mem_q[302] : 
                               (N858)? mem_q[665] : 
                               (N860)? mem_q[1028] : 
                               (N862)? mem_q[1391] : 
                               (N857)? mem_q[1754] : 
                               (N859)? mem_q[2117] : 
                               (N861)? mem_q[2480] : 
                               (N863)? mem_q[2843] : 1'b0;
  assign commit_instr_o[301] = (N856)? mem_q[301] : 
                               (N858)? mem_q[664] : 
                               (N860)? mem_q[1027] : 
                               (N862)? mem_q[1390] : 
                               (N857)? mem_q[1753] : 
                               (N859)? mem_q[2116] : 
                               (N861)? mem_q[2479] : 
                               (N863)? mem_q[2842] : 1'b0;
  assign commit_instr_o[300] = (N856)? mem_q[300] : 
                               (N858)? mem_q[663] : 
                               (N860)? mem_q[1026] : 
                               (N862)? mem_q[1389] : 
                               (N857)? mem_q[1752] : 
                               (N859)? mem_q[2115] : 
                               (N861)? mem_q[2478] : 
                               (N863)? mem_q[2841] : 1'b0;
  assign commit_instr_o[299] = (N856)? mem_q[299] : 
                               (N858)? mem_q[662] : 
                               (N860)? mem_q[1025] : 
                               (N862)? mem_q[1388] : 
                               (N857)? mem_q[1751] : 
                               (N859)? mem_q[2114] : 
                               (N861)? mem_q[2477] : 
                               (N863)? mem_q[2840] : 1'b0;
  assign commit_instr_o[298] = (N856)? mem_q[298] : 
                               (N858)? mem_q[661] : 
                               (N860)? mem_q[1024] : 
                               (N862)? mem_q[1387] : 
                               (N857)? mem_q[1750] : 
                               (N859)? mem_q[2113] : 
                               (N861)? mem_q[2476] : 
                               (N863)? mem_q[2839] : 1'b0;
  assign commit_instr_o[297] = (N856)? mem_q[297] : 
                               (N858)? mem_q[660] : 
                               (N860)? mem_q[1023] : 
                               (N862)? mem_q[1386] : 
                               (N857)? mem_q[1749] : 
                               (N859)? mem_q[2112] : 
                               (N861)? mem_q[2475] : 
                               (N863)? mem_q[2838] : 1'b0;
  assign commit_instr_o[296] = (N856)? mem_q[296] : 
                               (N858)? mem_q[659] : 
                               (N860)? mem_q[1022] : 
                               (N862)? mem_q[1385] : 
                               (N857)? mem_q[1748] : 
                               (N859)? mem_q[2111] : 
                               (N861)? mem_q[2474] : 
                               (N863)? mem_q[2837] : 1'b0;
  assign commit_instr_o[295] = (N856)? mem_q[295] : 
                               (N858)? mem_q[658] : 
                               (N860)? mem_q[1021] : 
                               (N862)? mem_q[1384] : 
                               (N857)? mem_q[1747] : 
                               (N859)? mem_q[2110] : 
                               (N861)? mem_q[2473] : 
                               (N863)? mem_q[2836] : 1'b0;
  assign commit_instr_o[294] = (N856)? mem_q[294] : 
                               (N858)? mem_q[657] : 
                               (N860)? mem_q[1020] : 
                               (N862)? mem_q[1383] : 
                               (N857)? mem_q[1746] : 
                               (N859)? mem_q[2109] : 
                               (N861)? mem_q[2472] : 
                               (N863)? mem_q[2835] : 1'b0;
  assign commit_instr_o[293] = (N856)? mem_q[293] : 
                               (N858)? mem_q[656] : 
                               (N860)? mem_q[1019] : 
                               (N862)? mem_q[1382] : 
                               (N857)? mem_q[1745] : 
                               (N859)? mem_q[2108] : 
                               (N861)? mem_q[2471] : 
                               (N863)? mem_q[2834] : 1'b0;
  assign commit_instr_o[292] = (N856)? mem_q[292] : 
                               (N858)? mem_q[655] : 
                               (N860)? mem_q[1018] : 
                               (N862)? mem_q[1381] : 
                               (N857)? mem_q[1744] : 
                               (N859)? mem_q[2107] : 
                               (N861)? mem_q[2470] : 
                               (N863)? mem_q[2833] : 1'b0;
  assign commit_instr_o[291] = (N856)? mem_q[291] : 
                               (N858)? mem_q[654] : 
                               (N860)? mem_q[1017] : 
                               (N862)? mem_q[1380] : 
                               (N857)? mem_q[1743] : 
                               (N859)? mem_q[2106] : 
                               (N861)? mem_q[2469] : 
                               (N863)? mem_q[2832] : 1'b0;
  assign commit_instr_o[290] = (N856)? mem_q[290] : 
                               (N858)? mem_q[653] : 
                               (N860)? mem_q[1016] : 
                               (N862)? mem_q[1379] : 
                               (N857)? mem_q[1742] : 
                               (N859)? mem_q[2105] : 
                               (N861)? mem_q[2468] : 
                               (N863)? mem_q[2831] : 1'b0;
  assign commit_instr_o[289] = (N856)? mem_q[289] : 
                               (N858)? mem_q[652] : 
                               (N860)? mem_q[1015] : 
                               (N862)? mem_q[1378] : 
                               (N857)? mem_q[1741] : 
                               (N859)? mem_q[2104] : 
                               (N861)? mem_q[2467] : 
                               (N863)? mem_q[2830] : 1'b0;
  assign commit_instr_o[288] = (N856)? mem_q[288] : 
                               (N858)? mem_q[651] : 
                               (N860)? mem_q[1014] : 
                               (N862)? mem_q[1377] : 
                               (N857)? mem_q[1740] : 
                               (N859)? mem_q[2103] : 
                               (N861)? mem_q[2466] : 
                               (N863)? mem_q[2829] : 1'b0;
  assign commit_instr_o[287] = (N856)? mem_q[287] : 
                               (N858)? mem_q[650] : 
                               (N860)? mem_q[1013] : 
                               (N862)? mem_q[1376] : 
                               (N857)? mem_q[1739] : 
                               (N859)? mem_q[2102] : 
                               (N861)? mem_q[2465] : 
                               (N863)? mem_q[2828] : 1'b0;
  assign commit_instr_o[286] = (N856)? mem_q[286] : 
                               (N858)? mem_q[649] : 
                               (N860)? mem_q[1012] : 
                               (N862)? mem_q[1375] : 
                               (N857)? mem_q[1738] : 
                               (N859)? mem_q[2101] : 
                               (N861)? mem_q[2464] : 
                               (N863)? mem_q[2827] : 1'b0;
  assign commit_instr_o[285] = (N856)? mem_q[285] : 
                               (N858)? mem_q[648] : 
                               (N860)? mem_q[1011] : 
                               (N862)? mem_q[1374] : 
                               (N857)? mem_q[1737] : 
                               (N859)? mem_q[2100] : 
                               (N861)? mem_q[2463] : 
                               (N863)? mem_q[2826] : 1'b0;
  assign commit_instr_o[284] = (N856)? mem_q[284] : 
                               (N858)? mem_q[647] : 
                               (N860)? mem_q[1010] : 
                               (N862)? mem_q[1373] : 
                               (N857)? mem_q[1736] : 
                               (N859)? mem_q[2099] : 
                               (N861)? mem_q[2462] : 
                               (N863)? mem_q[2825] : 1'b0;
  assign commit_instr_o[283] = (N856)? mem_q[283] : 
                               (N858)? mem_q[646] : 
                               (N860)? mem_q[1009] : 
                               (N862)? mem_q[1372] : 
                               (N857)? mem_q[1735] : 
                               (N859)? mem_q[2098] : 
                               (N861)? mem_q[2461] : 
                               (N863)? mem_q[2824] : 1'b0;
  assign commit_instr_o[282] = (N856)? mem_q[282] : 
                               (N858)? mem_q[645] : 
                               (N860)? mem_q[1008] : 
                               (N862)? mem_q[1371] : 
                               (N857)? mem_q[1734] : 
                               (N859)? mem_q[2097] : 
                               (N861)? mem_q[2460] : 
                               (N863)? mem_q[2823] : 1'b0;
  assign commit_instr_o[281] = (N856)? mem_q[281] : 
                               (N858)? mem_q[644] : 
                               (N860)? mem_q[1007] : 
                               (N862)? mem_q[1370] : 
                               (N857)? mem_q[1733] : 
                               (N859)? mem_q[2096] : 
                               (N861)? mem_q[2459] : 
                               (N863)? mem_q[2822] : 1'b0;
  assign commit_instr_o[280] = (N856)? mem_q[280] : 
                               (N858)? mem_q[643] : 
                               (N860)? mem_q[1006] : 
                               (N862)? mem_q[1369] : 
                               (N857)? mem_q[1732] : 
                               (N859)? mem_q[2095] : 
                               (N861)? mem_q[2458] : 
                               (N863)? mem_q[2821] : 1'b0;
  assign commit_instr_o[279] = (N856)? mem_q[279] : 
                               (N858)? mem_q[642] : 
                               (N860)? mem_q[1005] : 
                               (N862)? mem_q[1368] : 
                               (N857)? mem_q[1731] : 
                               (N859)? mem_q[2094] : 
                               (N861)? mem_q[2457] : 
                               (N863)? mem_q[2820] : 1'b0;
  assign commit_instr_o[278] = (N856)? mem_q[278] : 
                               (N858)? mem_q[641] : 
                               (N860)? mem_q[1004] : 
                               (N862)? mem_q[1367] : 
                               (N857)? mem_q[1730] : 
                               (N859)? mem_q[2093] : 
                               (N861)? mem_q[2456] : 
                               (N863)? mem_q[2819] : 1'b0;
  assign commit_instr_o[277] = (N856)? mem_q[277] : 
                               (N858)? mem_q[640] : 
                               (N860)? mem_q[1003] : 
                               (N862)? mem_q[1366] : 
                               (N857)? mem_q[1729] : 
                               (N859)? mem_q[2092] : 
                               (N861)? mem_q[2455] : 
                               (N863)? mem_q[2818] : 1'b0;
  assign commit_instr_o[276] = (N856)? mem_q[276] : 
                               (N858)? mem_q[639] : 
                               (N860)? mem_q[1002] : 
                               (N862)? mem_q[1365] : 
                               (N857)? mem_q[1728] : 
                               (N859)? mem_q[2091] : 
                               (N861)? mem_q[2454] : 
                               (N863)? mem_q[2817] : 1'b0;
  assign commit_instr_o[275] = (N856)? mem_q[275] : 
                               (N858)? mem_q[638] : 
                               (N860)? mem_q[1001] : 
                               (N862)? mem_q[1364] : 
                               (N857)? mem_q[1727] : 
                               (N859)? mem_q[2090] : 
                               (N861)? mem_q[2453] : 
                               (N863)? mem_q[2816] : 1'b0;
  assign commit_instr_o[274] = (N856)? mem_q[274] : 
                               (N858)? mem_q[637] : 
                               (N860)? mem_q[1000] : 
                               (N862)? mem_q[1363] : 
                               (N857)? mem_q[1726] : 
                               (N859)? mem_q[2089] : 
                               (N861)? mem_q[2452] : 
                               (N863)? mem_q[2815] : 1'b0;
  assign commit_instr_o[273] = (N856)? mem_q[273] : 
                               (N858)? mem_q[636] : 
                               (N860)? mem_q[999] : 
                               (N862)? mem_q[1362] : 
                               (N857)? mem_q[1725] : 
                               (N859)? mem_q[2088] : 
                               (N861)? mem_q[2451] : 
                               (N863)? mem_q[2814] : 1'b0;
  assign commit_instr_o[272] = (N856)? mem_q[272] : 
                               (N858)? mem_q[635] : 
                               (N860)? mem_q[998] : 
                               (N862)? mem_q[1361] : 
                               (N857)? mem_q[1724] : 
                               (N859)? mem_q[2087] : 
                               (N861)? mem_q[2450] : 
                               (N863)? mem_q[2813] : 1'b0;
  assign commit_instr_o[271] = (N856)? mem_q[271] : 
                               (N858)? mem_q[634] : 
                               (N860)? mem_q[997] : 
                               (N862)? mem_q[1360] : 
                               (N857)? mem_q[1723] : 
                               (N859)? mem_q[2086] : 
                               (N861)? mem_q[2449] : 
                               (N863)? mem_q[2812] : 1'b0;
  assign commit_instr_o[270] = (N856)? mem_q[270] : 
                               (N858)? mem_q[633] : 
                               (N860)? mem_q[996] : 
                               (N862)? mem_q[1359] : 
                               (N857)? mem_q[1722] : 
                               (N859)? mem_q[2085] : 
                               (N861)? mem_q[2448] : 
                               (N863)? mem_q[2811] : 1'b0;
  assign commit_instr_o[269] = (N856)? mem_q[269] : 
                               (N858)? mem_q[632] : 
                               (N860)? mem_q[995] : 
                               (N862)? mem_q[1358] : 
                               (N857)? mem_q[1721] : 
                               (N859)? mem_q[2084] : 
                               (N861)? mem_q[2447] : 
                               (N863)? mem_q[2810] : 1'b0;
  assign commit_instr_o[268] = (N856)? mem_q[268] : 
                               (N858)? mem_q[631] : 
                               (N860)? mem_q[994] : 
                               (N862)? mem_q[1357] : 
                               (N857)? mem_q[1720] : 
                               (N859)? mem_q[2083] : 
                               (N861)? mem_q[2446] : 
                               (N863)? mem_q[2809] : 1'b0;
  assign commit_instr_o[267] = (N856)? mem_q[267] : 
                               (N858)? mem_q[630] : 
                               (N860)? mem_q[993] : 
                               (N862)? mem_q[1356] : 
                               (N857)? mem_q[1719] : 
                               (N859)? mem_q[2082] : 
                               (N861)? mem_q[2445] : 
                               (N863)? mem_q[2808] : 1'b0;
  assign commit_instr_o[266] = (N856)? mem_q[266] : 
                               (N858)? mem_q[629] : 
                               (N860)? mem_q[992] : 
                               (N862)? mem_q[1355] : 
                               (N857)? mem_q[1718] : 
                               (N859)? mem_q[2081] : 
                               (N861)? mem_q[2444] : 
                               (N863)? mem_q[2807] : 1'b0;
  assign commit_instr_o[265] = (N856)? mem_q[265] : 
                               (N858)? mem_q[628] : 
                               (N860)? mem_q[991] : 
                               (N862)? mem_q[1354] : 
                               (N857)? mem_q[1717] : 
                               (N859)? mem_q[2080] : 
                               (N861)? mem_q[2443] : 
                               (N863)? mem_q[2806] : 1'b0;
  assign commit_instr_o[264] = (N856)? mem_q[264] : 
                               (N858)? mem_q[627] : 
                               (N860)? mem_q[990] : 
                               (N862)? mem_q[1353] : 
                               (N857)? mem_q[1716] : 
                               (N859)? mem_q[2079] : 
                               (N861)? mem_q[2442] : 
                               (N863)? mem_q[2805] : 1'b0;
  assign commit_instr_o[263] = (N856)? mem_q[263] : 
                               (N858)? mem_q[626] : 
                               (N860)? mem_q[989] : 
                               (N862)? mem_q[1352] : 
                               (N857)? mem_q[1715] : 
                               (N859)? mem_q[2078] : 
                               (N861)? mem_q[2441] : 
                               (N863)? mem_q[2804] : 1'b0;
  assign commit_instr_o[262] = (N856)? mem_q[262] : 
                               (N858)? mem_q[625] : 
                               (N860)? mem_q[988] : 
                               (N862)? mem_q[1351] : 
                               (N857)? mem_q[1714] : 
                               (N859)? mem_q[2077] : 
                               (N861)? mem_q[2440] : 
                               (N863)? mem_q[2803] : 1'b0;
  assign commit_instr_o[261] = (N856)? mem_q[261] : 
                               (N858)? mem_q[624] : 
                               (N860)? mem_q[987] : 
                               (N862)? mem_q[1350] : 
                               (N857)? mem_q[1713] : 
                               (N859)? mem_q[2076] : 
                               (N861)? mem_q[2439] : 
                               (N863)? mem_q[2802] : 1'b0;
  assign commit_instr_o[260] = (N856)? mem_q[260] : 
                               (N858)? mem_q[623] : 
                               (N860)? mem_q[986] : 
                               (N862)? mem_q[1349] : 
                               (N857)? mem_q[1712] : 
                               (N859)? mem_q[2075] : 
                               (N861)? mem_q[2438] : 
                               (N863)? mem_q[2801] : 1'b0;
  assign commit_instr_o[259] = (N856)? mem_q[259] : 
                               (N858)? mem_q[622] : 
                               (N860)? mem_q[985] : 
                               (N862)? mem_q[1348] : 
                               (N857)? mem_q[1711] : 
                               (N859)? mem_q[2074] : 
                               (N861)? mem_q[2437] : 
                               (N863)? mem_q[2800] : 1'b0;
  assign commit_instr_o[258] = (N856)? mem_q[258] : 
                               (N858)? mem_q[621] : 
                               (N860)? mem_q[984] : 
                               (N862)? mem_q[1347] : 
                               (N857)? mem_q[1710] : 
                               (N859)? mem_q[2073] : 
                               (N861)? mem_q[2436] : 
                               (N863)? mem_q[2799] : 1'b0;
  assign commit_instr_o[257] = (N856)? mem_q[257] : 
                               (N858)? mem_q[620] : 
                               (N860)? mem_q[983] : 
                               (N862)? mem_q[1346] : 
                               (N857)? mem_q[1709] : 
                               (N859)? mem_q[2072] : 
                               (N861)? mem_q[2435] : 
                               (N863)? mem_q[2798] : 1'b0;
  assign commit_instr_o[256] = (N856)? mem_q[256] : 
                               (N858)? mem_q[619] : 
                               (N860)? mem_q[982] : 
                               (N862)? mem_q[1345] : 
                               (N857)? mem_q[1708] : 
                               (N859)? mem_q[2071] : 
                               (N861)? mem_q[2434] : 
                               (N863)? mem_q[2797] : 1'b0;
  assign commit_instr_o[255] = (N856)? mem_q[255] : 
                               (N858)? mem_q[618] : 
                               (N860)? mem_q[981] : 
                               (N862)? mem_q[1344] : 
                               (N857)? mem_q[1707] : 
                               (N859)? mem_q[2070] : 
                               (N861)? mem_q[2433] : 
                               (N863)? mem_q[2796] : 1'b0;
  assign commit_instr_o[254] = (N856)? mem_q[254] : 
                               (N858)? mem_q[617] : 
                               (N860)? mem_q[980] : 
                               (N862)? mem_q[1343] : 
                               (N857)? mem_q[1706] : 
                               (N859)? mem_q[2069] : 
                               (N861)? mem_q[2432] : 
                               (N863)? mem_q[2795] : 1'b0;
  assign commit_instr_o[253] = (N856)? mem_q[253] : 
                               (N858)? mem_q[616] : 
                               (N860)? mem_q[979] : 
                               (N862)? mem_q[1342] : 
                               (N857)? mem_q[1705] : 
                               (N859)? mem_q[2068] : 
                               (N861)? mem_q[2431] : 
                               (N863)? mem_q[2794] : 1'b0;
  assign commit_instr_o[252] = (N856)? mem_q[252] : 
                               (N858)? mem_q[615] : 
                               (N860)? mem_q[978] : 
                               (N862)? mem_q[1341] : 
                               (N857)? mem_q[1704] : 
                               (N859)? mem_q[2067] : 
                               (N861)? mem_q[2430] : 
                               (N863)? mem_q[2793] : 1'b0;
  assign commit_instr_o[251] = (N856)? mem_q[251] : 
                               (N858)? mem_q[614] : 
                               (N860)? mem_q[977] : 
                               (N862)? mem_q[1340] : 
                               (N857)? mem_q[1703] : 
                               (N859)? mem_q[2066] : 
                               (N861)? mem_q[2429] : 
                               (N863)? mem_q[2792] : 1'b0;
  assign commit_instr_o[250] = (N856)? mem_q[250] : 
                               (N858)? mem_q[613] : 
                               (N860)? mem_q[976] : 
                               (N862)? mem_q[1339] : 
                               (N857)? mem_q[1702] : 
                               (N859)? mem_q[2065] : 
                               (N861)? mem_q[2428] : 
                               (N863)? mem_q[2791] : 1'b0;
  assign commit_instr_o[249] = (N856)? mem_q[249] : 
                               (N858)? mem_q[612] : 
                               (N860)? mem_q[975] : 
                               (N862)? mem_q[1338] : 
                               (N857)? mem_q[1701] : 
                               (N859)? mem_q[2064] : 
                               (N861)? mem_q[2427] : 
                               (N863)? mem_q[2790] : 1'b0;
  assign commit_instr_o[248] = (N856)? mem_q[248] : 
                               (N858)? mem_q[611] : 
                               (N860)? mem_q[974] : 
                               (N862)? mem_q[1337] : 
                               (N857)? mem_q[1700] : 
                               (N859)? mem_q[2063] : 
                               (N861)? mem_q[2426] : 
                               (N863)? mem_q[2789] : 1'b0;
  assign commit_instr_o[247] = (N856)? mem_q[247] : 
                               (N858)? mem_q[610] : 
                               (N860)? mem_q[973] : 
                               (N862)? mem_q[1336] : 
                               (N857)? mem_q[1699] : 
                               (N859)? mem_q[2062] : 
                               (N861)? mem_q[2425] : 
                               (N863)? mem_q[2788] : 1'b0;
  assign commit_instr_o[246] = (N856)? mem_q[246] : 
                               (N858)? mem_q[609] : 
                               (N860)? mem_q[972] : 
                               (N862)? mem_q[1335] : 
                               (N857)? mem_q[1698] : 
                               (N859)? mem_q[2061] : 
                               (N861)? mem_q[2424] : 
                               (N863)? mem_q[2787] : 1'b0;
  assign commit_instr_o[245] = (N856)? mem_q[245] : 
                               (N858)? mem_q[608] : 
                               (N860)? mem_q[971] : 
                               (N862)? mem_q[1334] : 
                               (N857)? mem_q[1697] : 
                               (N859)? mem_q[2060] : 
                               (N861)? mem_q[2423] : 
                               (N863)? mem_q[2786] : 1'b0;
  assign commit_instr_o[244] = (N856)? mem_q[244] : 
                               (N858)? mem_q[607] : 
                               (N860)? mem_q[970] : 
                               (N862)? mem_q[1333] : 
                               (N857)? mem_q[1696] : 
                               (N859)? mem_q[2059] : 
                               (N861)? mem_q[2422] : 
                               (N863)? mem_q[2785] : 1'b0;
  assign commit_instr_o[243] = (N856)? mem_q[243] : 
                               (N858)? mem_q[606] : 
                               (N860)? mem_q[969] : 
                               (N862)? mem_q[1332] : 
                               (N857)? mem_q[1695] : 
                               (N859)? mem_q[2058] : 
                               (N861)? mem_q[2421] : 
                               (N863)? mem_q[2784] : 1'b0;
  assign commit_instr_o[242] = (N856)? mem_q[242] : 
                               (N858)? mem_q[605] : 
                               (N860)? mem_q[968] : 
                               (N862)? mem_q[1331] : 
                               (N857)? mem_q[1694] : 
                               (N859)? mem_q[2057] : 
                               (N861)? mem_q[2420] : 
                               (N863)? mem_q[2783] : 1'b0;
  assign commit_instr_o[241] = (N856)? mem_q[241] : 
                               (N858)? mem_q[604] : 
                               (N860)? mem_q[967] : 
                               (N862)? mem_q[1330] : 
                               (N857)? mem_q[1693] : 
                               (N859)? mem_q[2056] : 
                               (N861)? mem_q[2419] : 
                               (N863)? mem_q[2782] : 1'b0;
  assign commit_instr_o[240] = (N856)? mem_q[240] : 
                               (N858)? mem_q[603] : 
                               (N860)? mem_q[966] : 
                               (N862)? mem_q[1329] : 
                               (N857)? mem_q[1692] : 
                               (N859)? mem_q[2055] : 
                               (N861)? mem_q[2418] : 
                               (N863)? mem_q[2781] : 1'b0;
  assign commit_instr_o[239] = (N856)? mem_q[239] : 
                               (N858)? mem_q[602] : 
                               (N860)? mem_q[965] : 
                               (N862)? mem_q[1328] : 
                               (N857)? mem_q[1691] : 
                               (N859)? mem_q[2054] : 
                               (N861)? mem_q[2417] : 
                               (N863)? mem_q[2780] : 1'b0;
  assign commit_instr_o[238] = (N856)? mem_q[238] : 
                               (N858)? mem_q[601] : 
                               (N860)? mem_q[964] : 
                               (N862)? mem_q[1327] : 
                               (N857)? mem_q[1690] : 
                               (N859)? mem_q[2053] : 
                               (N861)? mem_q[2416] : 
                               (N863)? mem_q[2779] : 1'b0;
  assign commit_instr_o[237] = (N856)? mem_q[237] : 
                               (N858)? mem_q[600] : 
                               (N860)? mem_q[963] : 
                               (N862)? mem_q[1326] : 
                               (N857)? mem_q[1689] : 
                               (N859)? mem_q[2052] : 
                               (N861)? mem_q[2415] : 
                               (N863)? mem_q[2778] : 1'b0;
  assign commit_instr_o[236] = (N856)? mem_q[236] : 
                               (N858)? mem_q[599] : 
                               (N860)? mem_q[962] : 
                               (N862)? mem_q[1325] : 
                               (N857)? mem_q[1688] : 
                               (N859)? mem_q[2051] : 
                               (N861)? mem_q[2414] : 
                               (N863)? mem_q[2777] : 1'b0;
  assign commit_instr_o[235] = (N856)? mem_q[235] : 
                               (N858)? mem_q[598] : 
                               (N860)? mem_q[961] : 
                               (N862)? mem_q[1324] : 
                               (N857)? mem_q[1687] : 
                               (N859)? mem_q[2050] : 
                               (N861)? mem_q[2413] : 
                               (N863)? mem_q[2776] : 1'b0;
  assign commit_instr_o[234] = (N856)? mem_q[234] : 
                               (N858)? mem_q[597] : 
                               (N860)? mem_q[960] : 
                               (N862)? mem_q[1323] : 
                               (N857)? mem_q[1686] : 
                               (N859)? mem_q[2049] : 
                               (N861)? mem_q[2412] : 
                               (N863)? mem_q[2775] : 1'b0;
  assign commit_instr_o[233] = (N856)? mem_q[233] : 
                               (N858)? mem_q[596] : 
                               (N860)? mem_q[959] : 
                               (N862)? mem_q[1322] : 
                               (N857)? mem_q[1685] : 
                               (N859)? mem_q[2048] : 
                               (N861)? mem_q[2411] : 
                               (N863)? mem_q[2774] : 1'b0;
  assign commit_instr_o[232] = (N856)? mem_q[232] : 
                               (N858)? mem_q[595] : 
                               (N860)? mem_q[958] : 
                               (N862)? mem_q[1321] : 
                               (N857)? mem_q[1684] : 
                               (N859)? mem_q[2047] : 
                               (N861)? mem_q[2410] : 
                               (N863)? mem_q[2773] : 1'b0;
  assign commit_instr_o[231] = (N856)? mem_q[231] : 
                               (N858)? mem_q[594] : 
                               (N860)? mem_q[957] : 
                               (N862)? mem_q[1320] : 
                               (N857)? mem_q[1683] : 
                               (N859)? mem_q[2046] : 
                               (N861)? mem_q[2409] : 
                               (N863)? mem_q[2772] : 1'b0;
  assign commit_instr_o[230] = (N856)? mem_q[230] : 
                               (N858)? mem_q[593] : 
                               (N860)? mem_q[956] : 
                               (N862)? mem_q[1319] : 
                               (N857)? mem_q[1682] : 
                               (N859)? mem_q[2045] : 
                               (N861)? mem_q[2408] : 
                               (N863)? mem_q[2771] : 1'b0;
  assign commit_instr_o[229] = (N856)? mem_q[229] : 
                               (N858)? mem_q[592] : 
                               (N860)? mem_q[955] : 
                               (N862)? mem_q[1318] : 
                               (N857)? mem_q[1681] : 
                               (N859)? mem_q[2044] : 
                               (N861)? mem_q[2407] : 
                               (N863)? mem_q[2770] : 1'b0;
  assign commit_instr_o[228] = (N856)? mem_q[228] : 
                               (N858)? mem_q[591] : 
                               (N860)? mem_q[954] : 
                               (N862)? mem_q[1317] : 
                               (N857)? mem_q[1680] : 
                               (N859)? mem_q[2043] : 
                               (N861)? mem_q[2406] : 
                               (N863)? mem_q[2769] : 1'b0;
  assign commit_instr_o[227] = (N856)? mem_q[227] : 
                               (N858)? mem_q[590] : 
                               (N860)? mem_q[953] : 
                               (N862)? mem_q[1316] : 
                               (N857)? mem_q[1679] : 
                               (N859)? mem_q[2042] : 
                               (N861)? mem_q[2405] : 
                               (N863)? mem_q[2768] : 1'b0;
  assign commit_instr_o[226] = (N856)? mem_q[226] : 
                               (N858)? mem_q[589] : 
                               (N860)? mem_q[952] : 
                               (N862)? mem_q[1315] : 
                               (N857)? mem_q[1678] : 
                               (N859)? mem_q[2041] : 
                               (N861)? mem_q[2404] : 
                               (N863)? mem_q[2767] : 1'b0;
  assign commit_instr_o[225] = (N856)? mem_q[225] : 
                               (N858)? mem_q[588] : 
                               (N860)? mem_q[951] : 
                               (N862)? mem_q[1314] : 
                               (N857)? mem_q[1677] : 
                               (N859)? mem_q[2040] : 
                               (N861)? mem_q[2403] : 
                               (N863)? mem_q[2766] : 1'b0;
  assign commit_instr_o[224] = (N856)? mem_q[224] : 
                               (N858)? mem_q[587] : 
                               (N860)? mem_q[950] : 
                               (N862)? mem_q[1313] : 
                               (N857)? mem_q[1676] : 
                               (N859)? mem_q[2039] : 
                               (N861)? mem_q[2402] : 
                               (N863)? mem_q[2765] : 1'b0;
  assign commit_instr_o[223] = (N856)? mem_q[223] : 
                               (N858)? mem_q[586] : 
                               (N860)? mem_q[949] : 
                               (N862)? mem_q[1312] : 
                               (N857)? mem_q[1675] : 
                               (N859)? mem_q[2038] : 
                               (N861)? mem_q[2401] : 
                               (N863)? mem_q[2764] : 1'b0;
  assign commit_instr_o[222] = (N856)? mem_q[222] : 
                               (N858)? mem_q[585] : 
                               (N860)? mem_q[948] : 
                               (N862)? mem_q[1311] : 
                               (N857)? mem_q[1674] : 
                               (N859)? mem_q[2037] : 
                               (N861)? mem_q[2400] : 
                               (N863)? mem_q[2763] : 1'b0;
  assign commit_instr_o[221] = (N856)? mem_q[221] : 
                               (N858)? mem_q[584] : 
                               (N860)? mem_q[947] : 
                               (N862)? mem_q[1310] : 
                               (N857)? mem_q[1673] : 
                               (N859)? mem_q[2036] : 
                               (N861)? mem_q[2399] : 
                               (N863)? mem_q[2762] : 1'b0;
  assign commit_instr_o[220] = (N856)? mem_q[220] : 
                               (N858)? mem_q[583] : 
                               (N860)? mem_q[946] : 
                               (N862)? mem_q[1309] : 
                               (N857)? mem_q[1672] : 
                               (N859)? mem_q[2035] : 
                               (N861)? mem_q[2398] : 
                               (N863)? mem_q[2761] : 1'b0;
  assign commit_instr_o[219] = (N856)? mem_q[219] : 
                               (N858)? mem_q[582] : 
                               (N860)? mem_q[945] : 
                               (N862)? mem_q[1308] : 
                               (N857)? mem_q[1671] : 
                               (N859)? mem_q[2034] : 
                               (N861)? mem_q[2397] : 
                               (N863)? mem_q[2760] : 1'b0;
  assign commit_instr_o[218] = (N856)? mem_q[218] : 
                               (N858)? mem_q[581] : 
                               (N860)? mem_q[944] : 
                               (N862)? mem_q[1307] : 
                               (N857)? mem_q[1670] : 
                               (N859)? mem_q[2033] : 
                               (N861)? mem_q[2396] : 
                               (N863)? mem_q[2759] : 1'b0;
  assign commit_instr_o[217] = (N856)? mem_q[217] : 
                               (N858)? mem_q[580] : 
                               (N860)? mem_q[943] : 
                               (N862)? mem_q[1306] : 
                               (N857)? mem_q[1669] : 
                               (N859)? mem_q[2032] : 
                               (N861)? mem_q[2395] : 
                               (N863)? mem_q[2758] : 1'b0;
  assign commit_instr_o[216] = (N856)? mem_q[216] : 
                               (N858)? mem_q[579] : 
                               (N860)? mem_q[942] : 
                               (N862)? mem_q[1305] : 
                               (N857)? mem_q[1668] : 
                               (N859)? mem_q[2031] : 
                               (N861)? mem_q[2394] : 
                               (N863)? mem_q[2757] : 1'b0;
  assign commit_instr_o[215] = (N856)? mem_q[215] : 
                               (N858)? mem_q[578] : 
                               (N860)? mem_q[941] : 
                               (N862)? mem_q[1304] : 
                               (N857)? mem_q[1667] : 
                               (N859)? mem_q[2030] : 
                               (N861)? mem_q[2393] : 
                               (N863)? mem_q[2756] : 1'b0;
  assign commit_instr_o[214] = (N856)? mem_q[214] : 
                               (N858)? mem_q[577] : 
                               (N860)? mem_q[940] : 
                               (N862)? mem_q[1303] : 
                               (N857)? mem_q[1666] : 
                               (N859)? mem_q[2029] : 
                               (N861)? mem_q[2392] : 
                               (N863)? mem_q[2755] : 1'b0;
  assign commit_instr_o[213] = (N856)? mem_q[213] : 
                               (N858)? mem_q[576] : 
                               (N860)? mem_q[939] : 
                               (N862)? mem_q[1302] : 
                               (N857)? mem_q[1665] : 
                               (N859)? mem_q[2028] : 
                               (N861)? mem_q[2391] : 
                               (N863)? mem_q[2754] : 1'b0;
  assign commit_instr_o[212] = (N856)? mem_q[212] : 
                               (N858)? mem_q[575] : 
                               (N860)? mem_q[938] : 
                               (N862)? mem_q[1301] : 
                               (N857)? mem_q[1664] : 
                               (N859)? mem_q[2027] : 
                               (N861)? mem_q[2390] : 
                               (N863)? mem_q[2753] : 1'b0;
  assign commit_instr_o[211] = (N856)? mem_q[211] : 
                               (N858)? mem_q[574] : 
                               (N860)? mem_q[937] : 
                               (N862)? mem_q[1300] : 
                               (N857)? mem_q[1663] : 
                               (N859)? mem_q[2026] : 
                               (N861)? mem_q[2389] : 
                               (N863)? mem_q[2752] : 1'b0;
  assign commit_instr_o[210] = (N856)? mem_q[210] : 
                               (N858)? mem_q[573] : 
                               (N860)? mem_q[936] : 
                               (N862)? mem_q[1299] : 
                               (N857)? mem_q[1662] : 
                               (N859)? mem_q[2025] : 
                               (N861)? mem_q[2388] : 
                               (N863)? mem_q[2751] : 1'b0;
  assign commit_instr_o[209] = (N856)? mem_q[209] : 
                               (N858)? mem_q[572] : 
                               (N860)? mem_q[935] : 
                               (N862)? mem_q[1298] : 
                               (N857)? mem_q[1661] : 
                               (N859)? mem_q[2024] : 
                               (N861)? mem_q[2387] : 
                               (N863)? mem_q[2750] : 1'b0;
  assign commit_instr_o[208] = (N856)? mem_q[208] : 
                               (N858)? mem_q[571] : 
                               (N860)? mem_q[934] : 
                               (N862)? mem_q[1297] : 
                               (N857)? mem_q[1660] : 
                               (N859)? mem_q[2023] : 
                               (N861)? mem_q[2386] : 
                               (N863)? mem_q[2749] : 1'b0;
  assign commit_instr_o[207] = (N856)? mem_q[207] : 
                               (N858)? mem_q[570] : 
                               (N860)? mem_q[933] : 
                               (N862)? mem_q[1296] : 
                               (N857)? mem_q[1659] : 
                               (N859)? mem_q[2022] : 
                               (N861)? mem_q[2385] : 
                               (N863)? mem_q[2748] : 1'b0;
  assign commit_instr_o[206] = (N856)? mem_q[206] : 
                               (N858)? mem_q[569] : 
                               (N860)? mem_q[932] : 
                               (N862)? mem_q[1295] : 
                               (N857)? mem_q[1658] : 
                               (N859)? mem_q[2021] : 
                               (N861)? mem_q[2384] : 
                               (N863)? mem_q[2747] : 1'b0;
  assign commit_instr_o[205] = (N856)? mem_q[205] : 
                               (N858)? mem_q[568] : 
                               (N860)? mem_q[931] : 
                               (N862)? mem_q[1294] : 
                               (N857)? mem_q[1657] : 
                               (N859)? mem_q[2020] : 
                               (N861)? mem_q[2383] : 
                               (N863)? mem_q[2746] : 1'b0;
  assign commit_instr_o[204] = (N856)? mem_q[204] : 
                               (N858)? mem_q[567] : 
                               (N860)? mem_q[930] : 
                               (N862)? mem_q[1293] : 
                               (N857)? mem_q[1656] : 
                               (N859)? mem_q[2019] : 
                               (N861)? mem_q[2382] : 
                               (N863)? mem_q[2745] : 1'b0;
  assign commit_instr_o[203] = (N856)? mem_q[203] : 
                               (N858)? mem_q[566] : 
                               (N860)? mem_q[929] : 
                               (N862)? mem_q[1292] : 
                               (N857)? mem_q[1655] : 
                               (N859)? mem_q[2018] : 
                               (N861)? mem_q[2381] : 
                               (N863)? mem_q[2744] : 1'b0;
  assign commit_instr_o[202] = (N856)? mem_q[202] : 
                               (N858)? mem_q[565] : 
                               (N860)? mem_q[928] : 
                               (N862)? mem_q[1291] : 
                               (N857)? mem_q[1654] : 
                               (N859)? mem_q[2017] : 
                               (N861)? mem_q[2380] : 
                               (N863)? mem_q[2743] : 1'b0;
  assign commit_instr_o[201] = (N856)? mem_q[201] : 
                               (N858)? mem_q[564] : 
                               (N860)? mem_q[927] : 
                               (N862)? mem_q[1290] : 
                               (N857)? mem_q[1653] : 
                               (N859)? mem_q[2016] : 
                               (N861)? mem_q[2379] : 
                               (N863)? mem_q[2742] : 1'b0;
  assign commit_instr_o[200] = (N856)? mem_q[200] : 
                               (N858)? mem_q[563] : 
                               (N860)? mem_q[926] : 
                               (N862)? mem_q[1289] : 
                               (N857)? mem_q[1652] : 
                               (N859)? mem_q[2015] : 
                               (N861)? mem_q[2378] : 
                               (N863)? mem_q[2741] : 1'b0;
  assign commit_instr_o[199] = (N856)? mem_q[199] : 
                               (N858)? mem_q[562] : 
                               (N860)? mem_q[925] : 
                               (N862)? mem_q[1288] : 
                               (N857)? mem_q[1651] : 
                               (N859)? mem_q[2014] : 
                               (N861)? mem_q[2377] : 
                               (N863)? mem_q[2740] : 1'b0;
  assign commit_instr_o[198] = (N856)? mem_q[198] : 
                               (N858)? mem_q[561] : 
                               (N860)? mem_q[924] : 
                               (N862)? mem_q[1287] : 
                               (N857)? mem_q[1650] : 
                               (N859)? mem_q[2013] : 
                               (N861)? mem_q[2376] : 
                               (N863)? mem_q[2739] : 1'b0;
  assign commit_instr_o[197] = (N856)? mem_q[197] : 
                               (N858)? mem_q[560] : 
                               (N860)? mem_q[923] : 
                               (N862)? mem_q[1286] : 
                               (N857)? mem_q[1649] : 
                               (N859)? mem_q[2012] : 
                               (N861)? mem_q[2375] : 
                               (N863)? mem_q[2738] : 1'b0;
  assign commit_instr_o[196] = (N856)? mem_q[196] : 
                               (N858)? mem_q[559] : 
                               (N860)? mem_q[922] : 
                               (N862)? mem_q[1285] : 
                               (N857)? mem_q[1648] : 
                               (N859)? mem_q[2011] : 
                               (N861)? mem_q[2374] : 
                               (N863)? mem_q[2737] : 1'b0;
  assign commit_instr_o[195] = (N856)? mem_q[195] : 
                               (N858)? mem_q[558] : 
                               (N860)? mem_q[921] : 
                               (N862)? mem_q[1284] : 
                               (N857)? mem_q[1647] : 
                               (N859)? mem_q[2010] : 
                               (N861)? mem_q[2373] : 
                               (N863)? mem_q[2736] : 1'b0;
  assign commit_instr_o[194] = (N856)? mem_q[194] : 
                               (N858)? mem_q[557] : 
                               (N860)? mem_q[920] : 
                               (N862)? mem_q[1283] : 
                               (N857)? mem_q[1646] : 
                               (N859)? mem_q[2009] : 
                               (N861)? mem_q[2372] : 
                               (N863)? mem_q[2735] : 1'b0;
  assign commit_instr_o[193] = (N856)? mem_q[193] : 
                               (N858)? mem_q[556] : 
                               (N860)? mem_q[919] : 
                               (N862)? mem_q[1282] : 
                               (N857)? mem_q[1645] : 
                               (N859)? mem_q[2008] : 
                               (N861)? mem_q[2371] : 
                               (N863)? mem_q[2734] : 1'b0;
  assign commit_instr_o[192] = (N856)? mem_q[192] : 
                               (N858)? mem_q[555] : 
                               (N860)? mem_q[918] : 
                               (N862)? mem_q[1281] : 
                               (N857)? mem_q[1644] : 
                               (N859)? mem_q[2007] : 
                               (N861)? mem_q[2370] : 
                               (N863)? mem_q[2733] : 1'b0;
  assign commit_instr_o[191] = (N856)? mem_q[191] : 
                               (N858)? mem_q[554] : 
                               (N860)? mem_q[917] : 
                               (N862)? mem_q[1280] : 
                               (N857)? mem_q[1643] : 
                               (N859)? mem_q[2006] : 
                               (N861)? mem_q[2369] : 
                               (N863)? mem_q[2732] : 1'b0;
  assign commit_instr_o[190] = (N856)? mem_q[190] : 
                               (N858)? mem_q[553] : 
                               (N860)? mem_q[916] : 
                               (N862)? mem_q[1279] : 
                               (N857)? mem_q[1642] : 
                               (N859)? mem_q[2005] : 
                               (N861)? mem_q[2368] : 
                               (N863)? mem_q[2731] : 1'b0;
  assign commit_instr_o[189] = (N856)? mem_q[189] : 
                               (N858)? mem_q[552] : 
                               (N860)? mem_q[915] : 
                               (N862)? mem_q[1278] : 
                               (N857)? mem_q[1641] : 
                               (N859)? mem_q[2004] : 
                               (N861)? mem_q[2367] : 
                               (N863)? mem_q[2730] : 1'b0;
  assign commit_instr_o[188] = (N856)? mem_q[188] : 
                               (N858)? mem_q[551] : 
                               (N860)? mem_q[914] : 
                               (N862)? mem_q[1277] : 
                               (N857)? mem_q[1640] : 
                               (N859)? mem_q[2003] : 
                               (N861)? mem_q[2366] : 
                               (N863)? mem_q[2729] : 1'b0;
  assign commit_instr_o[187] = (N856)? mem_q[187] : 
                               (N858)? mem_q[550] : 
                               (N860)? mem_q[913] : 
                               (N862)? mem_q[1276] : 
                               (N857)? mem_q[1639] : 
                               (N859)? mem_q[2002] : 
                               (N861)? mem_q[2365] : 
                               (N863)? mem_q[2728] : 1'b0;
  assign commit_instr_o[186] = (N856)? mem_q[186] : 
                               (N858)? mem_q[549] : 
                               (N860)? mem_q[912] : 
                               (N862)? mem_q[1275] : 
                               (N857)? mem_q[1638] : 
                               (N859)? mem_q[2001] : 
                               (N861)? mem_q[2364] : 
                               (N863)? mem_q[2727] : 1'b0;
  assign commit_instr_o[185] = (N856)? mem_q[185] : 
                               (N858)? mem_q[548] : 
                               (N860)? mem_q[911] : 
                               (N862)? mem_q[1274] : 
                               (N857)? mem_q[1637] : 
                               (N859)? mem_q[2000] : 
                               (N861)? mem_q[2363] : 
                               (N863)? mem_q[2726] : 1'b0;
  assign commit_instr_o[184] = (N856)? mem_q[184] : 
                               (N858)? mem_q[547] : 
                               (N860)? mem_q[910] : 
                               (N862)? mem_q[1273] : 
                               (N857)? mem_q[1636] : 
                               (N859)? mem_q[1999] : 
                               (N861)? mem_q[2362] : 
                               (N863)? mem_q[2725] : 1'b0;
  assign commit_instr_o[183] = (N856)? mem_q[183] : 
                               (N858)? mem_q[546] : 
                               (N860)? mem_q[909] : 
                               (N862)? mem_q[1272] : 
                               (N857)? mem_q[1635] : 
                               (N859)? mem_q[1998] : 
                               (N861)? mem_q[2361] : 
                               (N863)? mem_q[2724] : 1'b0;
  assign commit_instr_o[182] = (N856)? mem_q[182] : 
                               (N858)? mem_q[545] : 
                               (N860)? mem_q[908] : 
                               (N862)? mem_q[1271] : 
                               (N857)? mem_q[1634] : 
                               (N859)? mem_q[1997] : 
                               (N861)? mem_q[2360] : 
                               (N863)? mem_q[2723] : 1'b0;
  assign commit_instr_o[181] = (N856)? mem_q[181] : 
                               (N858)? mem_q[544] : 
                               (N860)? mem_q[907] : 
                               (N862)? mem_q[1270] : 
                               (N857)? mem_q[1633] : 
                               (N859)? mem_q[1996] : 
                               (N861)? mem_q[2359] : 
                               (N863)? mem_q[2722] : 1'b0;
  assign commit_instr_o[180] = (N856)? mem_q[180] : 
                               (N858)? mem_q[543] : 
                               (N860)? mem_q[906] : 
                               (N862)? mem_q[1269] : 
                               (N857)? mem_q[1632] : 
                               (N859)? mem_q[1995] : 
                               (N861)? mem_q[2358] : 
                               (N863)? mem_q[2721] : 1'b0;
  assign commit_instr_o[179] = (N856)? mem_q[179] : 
                               (N858)? mem_q[542] : 
                               (N860)? mem_q[905] : 
                               (N862)? mem_q[1268] : 
                               (N857)? mem_q[1631] : 
                               (N859)? mem_q[1994] : 
                               (N861)? mem_q[2357] : 
                               (N863)? mem_q[2720] : 1'b0;
  assign commit_instr_o[178] = (N856)? mem_q[178] : 
                               (N858)? mem_q[541] : 
                               (N860)? mem_q[904] : 
                               (N862)? mem_q[1267] : 
                               (N857)? mem_q[1630] : 
                               (N859)? mem_q[1993] : 
                               (N861)? mem_q[2356] : 
                               (N863)? mem_q[2719] : 1'b0;
  assign commit_instr_o[177] = (N856)? mem_q[177] : 
                               (N858)? mem_q[540] : 
                               (N860)? mem_q[903] : 
                               (N862)? mem_q[1266] : 
                               (N857)? mem_q[1629] : 
                               (N859)? mem_q[1992] : 
                               (N861)? mem_q[2355] : 
                               (N863)? mem_q[2718] : 1'b0;
  assign commit_instr_o[176] = (N856)? mem_q[176] : 
                               (N858)? mem_q[539] : 
                               (N860)? mem_q[902] : 
                               (N862)? mem_q[1265] : 
                               (N857)? mem_q[1628] : 
                               (N859)? mem_q[1991] : 
                               (N861)? mem_q[2354] : 
                               (N863)? mem_q[2717] : 1'b0;
  assign commit_instr_o[175] = (N856)? mem_q[175] : 
                               (N858)? mem_q[538] : 
                               (N860)? mem_q[901] : 
                               (N862)? mem_q[1264] : 
                               (N857)? mem_q[1627] : 
                               (N859)? mem_q[1990] : 
                               (N861)? mem_q[2353] : 
                               (N863)? mem_q[2716] : 1'b0;
  assign commit_instr_o[174] = (N856)? mem_q[174] : 
                               (N858)? mem_q[537] : 
                               (N860)? mem_q[900] : 
                               (N862)? mem_q[1263] : 
                               (N857)? mem_q[1626] : 
                               (N859)? mem_q[1989] : 
                               (N861)? mem_q[2352] : 
                               (N863)? mem_q[2715] : 1'b0;
  assign commit_instr_o[173] = (N856)? mem_q[173] : 
                               (N858)? mem_q[536] : 
                               (N860)? mem_q[899] : 
                               (N862)? mem_q[1262] : 
                               (N857)? mem_q[1625] : 
                               (N859)? mem_q[1988] : 
                               (N861)? mem_q[2351] : 
                               (N863)? mem_q[2714] : 1'b0;
  assign commit_instr_o[172] = (N856)? mem_q[172] : 
                               (N858)? mem_q[535] : 
                               (N860)? mem_q[898] : 
                               (N862)? mem_q[1261] : 
                               (N857)? mem_q[1624] : 
                               (N859)? mem_q[1987] : 
                               (N861)? mem_q[2350] : 
                               (N863)? mem_q[2713] : 1'b0;
  assign commit_instr_o[171] = (N856)? mem_q[171] : 
                               (N858)? mem_q[534] : 
                               (N860)? mem_q[897] : 
                               (N862)? mem_q[1260] : 
                               (N857)? mem_q[1623] : 
                               (N859)? mem_q[1986] : 
                               (N861)? mem_q[2349] : 
                               (N863)? mem_q[2712] : 1'b0;
  assign commit_instr_o[170] = (N856)? mem_q[170] : 
                               (N858)? mem_q[533] : 
                               (N860)? mem_q[896] : 
                               (N862)? mem_q[1259] : 
                               (N857)? mem_q[1622] : 
                               (N859)? mem_q[1985] : 
                               (N861)? mem_q[2348] : 
                               (N863)? mem_q[2711] : 1'b0;
  assign commit_instr_o[169] = (N856)? mem_q[169] : 
                               (N858)? mem_q[532] : 
                               (N860)? mem_q[895] : 
                               (N862)? mem_q[1258] : 
                               (N857)? mem_q[1621] : 
                               (N859)? mem_q[1984] : 
                               (N861)? mem_q[2347] : 
                               (N863)? mem_q[2710] : 1'b0;
  assign commit_instr_o[168] = (N856)? mem_q[168] : 
                               (N858)? mem_q[531] : 
                               (N860)? mem_q[894] : 
                               (N862)? mem_q[1257] : 
                               (N857)? mem_q[1620] : 
                               (N859)? mem_q[1983] : 
                               (N861)? mem_q[2346] : 
                               (N863)? mem_q[2709] : 1'b0;
  assign commit_instr_o[167] = (N856)? mem_q[167] : 
                               (N858)? mem_q[530] : 
                               (N860)? mem_q[893] : 
                               (N862)? mem_q[1256] : 
                               (N857)? mem_q[1619] : 
                               (N859)? mem_q[1982] : 
                               (N861)? mem_q[2345] : 
                               (N863)? mem_q[2708] : 1'b0;
  assign commit_instr_o[166] = (N856)? mem_q[166] : 
                               (N858)? mem_q[529] : 
                               (N860)? mem_q[892] : 
                               (N862)? mem_q[1255] : 
                               (N857)? mem_q[1618] : 
                               (N859)? mem_q[1981] : 
                               (N861)? mem_q[2344] : 
                               (N863)? mem_q[2707] : 1'b0;
  assign commit_instr_o[165] = (N856)? mem_q[165] : 
                               (N858)? mem_q[528] : 
                               (N860)? mem_q[891] : 
                               (N862)? mem_q[1254] : 
                               (N857)? mem_q[1617] : 
                               (N859)? mem_q[1980] : 
                               (N861)? mem_q[2343] : 
                               (N863)? mem_q[2706] : 1'b0;
  assign commit_instr_o[164] = (N856)? mem_q[164] : 
                               (N858)? mem_q[527] : 
                               (N860)? mem_q[890] : 
                               (N862)? mem_q[1253] : 
                               (N857)? mem_q[1616] : 
                               (N859)? mem_q[1979] : 
                               (N861)? mem_q[2342] : 
                               (N863)? mem_q[2705] : 1'b0;
  assign commit_instr_o[163] = (N856)? mem_q[163] : 
                               (N858)? mem_q[526] : 
                               (N860)? mem_q[889] : 
                               (N862)? mem_q[1252] : 
                               (N857)? mem_q[1615] : 
                               (N859)? mem_q[1978] : 
                               (N861)? mem_q[2341] : 
                               (N863)? mem_q[2704] : 1'b0;
  assign commit_instr_o[162] = (N856)? mem_q[162] : 
                               (N858)? mem_q[525] : 
                               (N860)? mem_q[888] : 
                               (N862)? mem_q[1251] : 
                               (N857)? mem_q[1614] : 
                               (N859)? mem_q[1977] : 
                               (N861)? mem_q[2340] : 
                               (N863)? mem_q[2703] : 1'b0;
  assign commit_instr_o[161] = (N856)? mem_q[161] : 
                               (N858)? mem_q[524] : 
                               (N860)? mem_q[887] : 
                               (N862)? mem_q[1250] : 
                               (N857)? mem_q[1613] : 
                               (N859)? mem_q[1976] : 
                               (N861)? mem_q[2339] : 
                               (N863)? mem_q[2702] : 1'b0;
  assign commit_instr_o[160] = (N856)? mem_q[160] : 
                               (N858)? mem_q[523] : 
                               (N860)? mem_q[886] : 
                               (N862)? mem_q[1249] : 
                               (N857)? mem_q[1612] : 
                               (N859)? mem_q[1975] : 
                               (N861)? mem_q[2338] : 
                               (N863)? mem_q[2701] : 1'b0;
  assign commit_instr_o[159] = (N856)? mem_q[159] : 
                               (N858)? mem_q[522] : 
                               (N860)? mem_q[885] : 
                               (N862)? mem_q[1248] : 
                               (N857)? mem_q[1611] : 
                               (N859)? mem_q[1974] : 
                               (N861)? mem_q[2337] : 
                               (N863)? mem_q[2700] : 1'b0;
  assign commit_instr_o[158] = (N856)? mem_q[158] : 
                               (N858)? mem_q[521] : 
                               (N860)? mem_q[884] : 
                               (N862)? mem_q[1247] : 
                               (N857)? mem_q[1610] : 
                               (N859)? mem_q[1973] : 
                               (N861)? mem_q[2336] : 
                               (N863)? mem_q[2699] : 1'b0;
  assign commit_instr_o[157] = (N856)? mem_q[157] : 
                               (N858)? mem_q[520] : 
                               (N860)? mem_q[883] : 
                               (N862)? mem_q[1246] : 
                               (N857)? mem_q[1609] : 
                               (N859)? mem_q[1972] : 
                               (N861)? mem_q[2335] : 
                               (N863)? mem_q[2698] : 1'b0;
  assign commit_instr_o[156] = (N856)? mem_q[156] : 
                               (N858)? mem_q[519] : 
                               (N860)? mem_q[882] : 
                               (N862)? mem_q[1245] : 
                               (N857)? mem_q[1608] : 
                               (N859)? mem_q[1971] : 
                               (N861)? mem_q[2334] : 
                               (N863)? mem_q[2697] : 1'b0;
  assign commit_instr_o[155] = (N856)? mem_q[155] : 
                               (N858)? mem_q[518] : 
                               (N860)? mem_q[881] : 
                               (N862)? mem_q[1244] : 
                               (N857)? mem_q[1607] : 
                               (N859)? mem_q[1970] : 
                               (N861)? mem_q[2333] : 
                               (N863)? mem_q[2696] : 1'b0;
  assign commit_instr_o[154] = (N856)? mem_q[154] : 
                               (N858)? mem_q[517] : 
                               (N860)? mem_q[880] : 
                               (N862)? mem_q[1243] : 
                               (N857)? mem_q[1606] : 
                               (N859)? mem_q[1969] : 
                               (N861)? mem_q[2332] : 
                               (N863)? mem_q[2695] : 1'b0;
  assign commit_instr_o[153] = (N856)? mem_q[153] : 
                               (N858)? mem_q[516] : 
                               (N860)? mem_q[879] : 
                               (N862)? mem_q[1242] : 
                               (N857)? mem_q[1605] : 
                               (N859)? mem_q[1968] : 
                               (N861)? mem_q[2331] : 
                               (N863)? mem_q[2694] : 1'b0;
  assign commit_instr_o[152] = (N856)? mem_q[152] : 
                               (N858)? mem_q[515] : 
                               (N860)? mem_q[878] : 
                               (N862)? mem_q[1241] : 
                               (N857)? mem_q[1604] : 
                               (N859)? mem_q[1967] : 
                               (N861)? mem_q[2330] : 
                               (N863)? mem_q[2693] : 1'b0;
  assign commit_instr_o[151] = (N856)? mem_q[151] : 
                               (N858)? mem_q[514] : 
                               (N860)? mem_q[877] : 
                               (N862)? mem_q[1240] : 
                               (N857)? mem_q[1603] : 
                               (N859)? mem_q[1966] : 
                               (N861)? mem_q[2329] : 
                               (N863)? mem_q[2692] : 1'b0;
  assign commit_instr_o[150] = (N856)? mem_q[150] : 
                               (N858)? mem_q[513] : 
                               (N860)? mem_q[876] : 
                               (N862)? mem_q[1239] : 
                               (N857)? mem_q[1602] : 
                               (N859)? mem_q[1965] : 
                               (N861)? mem_q[2328] : 
                               (N863)? mem_q[2691] : 1'b0;
  assign commit_instr_o[149] = (N856)? mem_q[149] : 
                               (N858)? mem_q[512] : 
                               (N860)? mem_q[875] : 
                               (N862)? mem_q[1238] : 
                               (N857)? mem_q[1601] : 
                               (N859)? mem_q[1964] : 
                               (N861)? mem_q[2327] : 
                               (N863)? mem_q[2690] : 1'b0;
  assign commit_instr_o[148] = (N856)? mem_q[148] : 
                               (N858)? mem_q[511] : 
                               (N860)? mem_q[874] : 
                               (N862)? mem_q[1237] : 
                               (N857)? mem_q[1600] : 
                               (N859)? mem_q[1963] : 
                               (N861)? mem_q[2326] : 
                               (N863)? mem_q[2689] : 1'b0;
  assign commit_instr_o[147] = (N856)? mem_q[147] : 
                               (N858)? mem_q[510] : 
                               (N860)? mem_q[873] : 
                               (N862)? mem_q[1236] : 
                               (N857)? mem_q[1599] : 
                               (N859)? mem_q[1962] : 
                               (N861)? mem_q[2325] : 
                               (N863)? mem_q[2688] : 1'b0;
  assign commit_instr_o[146] = (N856)? mem_q[146] : 
                               (N858)? mem_q[509] : 
                               (N860)? mem_q[872] : 
                               (N862)? mem_q[1235] : 
                               (N857)? mem_q[1598] : 
                               (N859)? mem_q[1961] : 
                               (N861)? mem_q[2324] : 
                               (N863)? mem_q[2687] : 1'b0;
  assign commit_instr_o[145] = (N856)? mem_q[145] : 
                               (N858)? mem_q[508] : 
                               (N860)? mem_q[871] : 
                               (N862)? mem_q[1234] : 
                               (N857)? mem_q[1597] : 
                               (N859)? mem_q[1960] : 
                               (N861)? mem_q[2323] : 
                               (N863)? mem_q[2686] : 1'b0;
  assign commit_instr_o[144] = (N856)? mem_q[144] : 
                               (N858)? mem_q[507] : 
                               (N860)? mem_q[870] : 
                               (N862)? mem_q[1233] : 
                               (N857)? mem_q[1596] : 
                               (N859)? mem_q[1959] : 
                               (N861)? mem_q[2322] : 
                               (N863)? mem_q[2685] : 1'b0;
  assign commit_instr_o[143] = (N856)? mem_q[143] : 
                               (N858)? mem_q[506] : 
                               (N860)? mem_q[869] : 
                               (N862)? mem_q[1232] : 
                               (N857)? mem_q[1595] : 
                               (N859)? mem_q[1958] : 
                               (N861)? mem_q[2321] : 
                               (N863)? mem_q[2684] : 1'b0;
  assign commit_instr_o[142] = (N856)? mem_q[142] : 
                               (N858)? mem_q[505] : 
                               (N860)? mem_q[868] : 
                               (N862)? mem_q[1231] : 
                               (N857)? mem_q[1594] : 
                               (N859)? mem_q[1957] : 
                               (N861)? mem_q[2320] : 
                               (N863)? mem_q[2683] : 1'b0;
  assign commit_instr_o[141] = (N856)? mem_q[141] : 
                               (N858)? mem_q[504] : 
                               (N860)? mem_q[867] : 
                               (N862)? mem_q[1230] : 
                               (N857)? mem_q[1593] : 
                               (N859)? mem_q[1956] : 
                               (N861)? mem_q[2319] : 
                               (N863)? mem_q[2682] : 1'b0;
  assign commit_instr_o[140] = (N856)? mem_q[140] : 
                               (N858)? mem_q[503] : 
                               (N860)? mem_q[866] : 
                               (N862)? mem_q[1229] : 
                               (N857)? mem_q[1592] : 
                               (N859)? mem_q[1955] : 
                               (N861)? mem_q[2318] : 
                               (N863)? mem_q[2681] : 1'b0;
  assign commit_instr_o[139] = (N856)? mem_q[139] : 
                               (N858)? mem_q[502] : 
                               (N860)? mem_q[865] : 
                               (N862)? mem_q[1228] : 
                               (N857)? mem_q[1591] : 
                               (N859)? mem_q[1954] : 
                               (N861)? mem_q[2317] : 
                               (N863)? mem_q[2680] : 1'b0;
  assign commit_instr_o[138] = (N856)? mem_q[138] : 
                               (N858)? mem_q[501] : 
                               (N860)? mem_q[864] : 
                               (N862)? mem_q[1227] : 
                               (N857)? mem_q[1590] : 
                               (N859)? mem_q[1953] : 
                               (N861)? mem_q[2316] : 
                               (N863)? mem_q[2679] : 1'b0;
  assign commit_instr_o[137] = (N856)? mem_q[137] : 
                               (N858)? mem_q[500] : 
                               (N860)? mem_q[863] : 
                               (N862)? mem_q[1226] : 
                               (N857)? mem_q[1589] : 
                               (N859)? mem_q[1952] : 
                               (N861)? mem_q[2315] : 
                               (N863)? mem_q[2678] : 1'b0;
  assign commit_instr_o[136] = (N856)? mem_q[136] : 
                               (N858)? mem_q[499] : 
                               (N860)? mem_q[862] : 
                               (N862)? mem_q[1225] : 
                               (N857)? mem_q[1588] : 
                               (N859)? mem_q[1951] : 
                               (N861)? mem_q[2314] : 
                               (N863)? mem_q[2677] : 1'b0;
  assign commit_instr_o[135] = (N856)? mem_q[135] : 
                               (N858)? mem_q[498] : 
                               (N860)? mem_q[861] : 
                               (N862)? mem_q[1224] : 
                               (N857)? mem_q[1587] : 
                               (N859)? mem_q[1950] : 
                               (N861)? mem_q[2313] : 
                               (N863)? mem_q[2676] : 1'b0;
  assign commit_instr_o[134] = (N856)? mem_q[134] : 
                               (N858)? mem_q[497] : 
                               (N860)? mem_q[860] : 
                               (N862)? mem_q[1223] : 
                               (N857)? mem_q[1586] : 
                               (N859)? mem_q[1949] : 
                               (N861)? mem_q[2312] : 
                               (N863)? mem_q[2675] : 1'b0;
  assign commit_instr_o[133] = (N856)? mem_q[133] : 
                               (N858)? mem_q[496] : 
                               (N860)? mem_q[859] : 
                               (N862)? mem_q[1222] : 
                               (N857)? mem_q[1585] : 
                               (N859)? mem_q[1948] : 
                               (N861)? mem_q[2311] : 
                               (N863)? mem_q[2674] : 1'b0;
  assign commit_instr_o[132] = (N856)? mem_q[132] : 
                               (N858)? mem_q[495] : 
                               (N860)? mem_q[858] : 
                               (N862)? mem_q[1221] : 
                               (N857)? mem_q[1584] : 
                               (N859)? mem_q[1947] : 
                               (N861)? mem_q[2310] : 
                               (N863)? mem_q[2673] : 1'b0;
  assign commit_instr_o[131] = (N856)? mem_q[131] : 
                               (N858)? mem_q[494] : 
                               (N860)? mem_q[857] : 
                               (N862)? mem_q[1220] : 
                               (N857)? mem_q[1583] : 
                               (N859)? mem_q[1946] : 
                               (N861)? mem_q[2309] : 
                               (N863)? mem_q[2672] : 1'b0;
  assign commit_instr_o[130] = (N856)? mem_q[130] : 
                               (N858)? mem_q[493] : 
                               (N860)? mem_q[856] : 
                               (N862)? mem_q[1219] : 
                               (N857)? mem_q[1582] : 
                               (N859)? mem_q[1945] : 
                               (N861)? mem_q[2308] : 
                               (N863)? mem_q[2671] : 1'b0;
  assign commit_instr_o[129] = (N856)? mem_q[129] : 
                               (N858)? mem_q[492] : 
                               (N860)? mem_q[855] : 
                               (N862)? mem_q[1218] : 
                               (N857)? mem_q[1581] : 
                               (N859)? mem_q[1944] : 
                               (N861)? mem_q[2307] : 
                               (N863)? mem_q[2670] : 1'b0;
  assign commit_instr_o[128] = (N856)? mem_q[128] : 
                               (N858)? mem_q[491] : 
                               (N860)? mem_q[854] : 
                               (N862)? mem_q[1217] : 
                               (N857)? mem_q[1580] : 
                               (N859)? mem_q[1943] : 
                               (N861)? mem_q[2306] : 
                               (N863)? mem_q[2669] : 1'b0;
  assign commit_instr_o[127] = (N856)? mem_q[127] : 
                               (N858)? mem_q[490] : 
                               (N860)? mem_q[853] : 
                               (N862)? mem_q[1216] : 
                               (N857)? mem_q[1579] : 
                               (N859)? mem_q[1942] : 
                               (N861)? mem_q[2305] : 
                               (N863)? mem_q[2668] : 1'b0;
  assign commit_instr_o[126] = (N856)? mem_q[126] : 
                               (N858)? mem_q[489] : 
                               (N860)? mem_q[852] : 
                               (N862)? mem_q[1215] : 
                               (N857)? mem_q[1578] : 
                               (N859)? mem_q[1941] : 
                               (N861)? mem_q[2304] : 
                               (N863)? mem_q[2667] : 1'b0;
  assign commit_instr_o[125] = (N856)? mem_q[125] : 
                               (N858)? mem_q[488] : 
                               (N860)? mem_q[851] : 
                               (N862)? mem_q[1214] : 
                               (N857)? mem_q[1577] : 
                               (N859)? mem_q[1940] : 
                               (N861)? mem_q[2303] : 
                               (N863)? mem_q[2666] : 1'b0;
  assign commit_instr_o[124] = (N856)? mem_q[124] : 
                               (N858)? mem_q[487] : 
                               (N860)? mem_q[850] : 
                               (N862)? mem_q[1213] : 
                               (N857)? mem_q[1576] : 
                               (N859)? mem_q[1939] : 
                               (N861)? mem_q[2302] : 
                               (N863)? mem_q[2665] : 1'b0;
  assign commit_instr_o[123] = (N856)? mem_q[123] : 
                               (N858)? mem_q[486] : 
                               (N860)? mem_q[849] : 
                               (N862)? mem_q[1212] : 
                               (N857)? mem_q[1575] : 
                               (N859)? mem_q[1938] : 
                               (N861)? mem_q[2301] : 
                               (N863)? mem_q[2664] : 1'b0;
  assign commit_instr_o[122] = (N856)? mem_q[122] : 
                               (N858)? mem_q[485] : 
                               (N860)? mem_q[848] : 
                               (N862)? mem_q[1211] : 
                               (N857)? mem_q[1574] : 
                               (N859)? mem_q[1937] : 
                               (N861)? mem_q[2300] : 
                               (N863)? mem_q[2663] : 1'b0;
  assign commit_instr_o[121] = (N856)? mem_q[121] : 
                               (N858)? mem_q[484] : 
                               (N860)? mem_q[847] : 
                               (N862)? mem_q[1210] : 
                               (N857)? mem_q[1573] : 
                               (N859)? mem_q[1936] : 
                               (N861)? mem_q[2299] : 
                               (N863)? mem_q[2662] : 1'b0;
  assign commit_instr_o[120] = (N856)? mem_q[120] : 
                               (N858)? mem_q[483] : 
                               (N860)? mem_q[846] : 
                               (N862)? mem_q[1209] : 
                               (N857)? mem_q[1572] : 
                               (N859)? mem_q[1935] : 
                               (N861)? mem_q[2298] : 
                               (N863)? mem_q[2661] : 1'b0;
  assign commit_instr_o[119] = (N856)? mem_q[119] : 
                               (N858)? mem_q[482] : 
                               (N860)? mem_q[845] : 
                               (N862)? mem_q[1208] : 
                               (N857)? mem_q[1571] : 
                               (N859)? mem_q[1934] : 
                               (N861)? mem_q[2297] : 
                               (N863)? mem_q[2660] : 1'b0;
  assign commit_instr_o[118] = (N856)? mem_q[118] : 
                               (N858)? mem_q[481] : 
                               (N860)? mem_q[844] : 
                               (N862)? mem_q[1207] : 
                               (N857)? mem_q[1570] : 
                               (N859)? mem_q[1933] : 
                               (N861)? mem_q[2296] : 
                               (N863)? mem_q[2659] : 1'b0;
  assign commit_instr_o[117] = (N856)? mem_q[117] : 
                               (N858)? mem_q[480] : 
                               (N860)? mem_q[843] : 
                               (N862)? mem_q[1206] : 
                               (N857)? mem_q[1569] : 
                               (N859)? mem_q[1932] : 
                               (N861)? mem_q[2295] : 
                               (N863)? mem_q[2658] : 1'b0;
  assign commit_instr_o[116] = (N856)? mem_q[116] : 
                               (N858)? mem_q[479] : 
                               (N860)? mem_q[842] : 
                               (N862)? mem_q[1205] : 
                               (N857)? mem_q[1568] : 
                               (N859)? mem_q[1931] : 
                               (N861)? mem_q[2294] : 
                               (N863)? mem_q[2657] : 1'b0;
  assign commit_instr_o[115] = (N856)? mem_q[115] : 
                               (N858)? mem_q[478] : 
                               (N860)? mem_q[841] : 
                               (N862)? mem_q[1204] : 
                               (N857)? mem_q[1567] : 
                               (N859)? mem_q[1930] : 
                               (N861)? mem_q[2293] : 
                               (N863)? mem_q[2656] : 1'b0;
  assign commit_instr_o[114] = (N856)? mem_q[114] : 
                               (N858)? mem_q[477] : 
                               (N860)? mem_q[840] : 
                               (N862)? mem_q[1203] : 
                               (N857)? mem_q[1566] : 
                               (N859)? mem_q[1929] : 
                               (N861)? mem_q[2292] : 
                               (N863)? mem_q[2655] : 1'b0;
  assign commit_instr_o[113] = (N856)? mem_q[113] : 
                               (N858)? mem_q[476] : 
                               (N860)? mem_q[839] : 
                               (N862)? mem_q[1202] : 
                               (N857)? mem_q[1565] : 
                               (N859)? mem_q[1928] : 
                               (N861)? mem_q[2291] : 
                               (N863)? mem_q[2654] : 1'b0;
  assign commit_instr_o[112] = (N856)? mem_q[112] : 
                               (N858)? mem_q[475] : 
                               (N860)? mem_q[838] : 
                               (N862)? mem_q[1201] : 
                               (N857)? mem_q[1564] : 
                               (N859)? mem_q[1927] : 
                               (N861)? mem_q[2290] : 
                               (N863)? mem_q[2653] : 1'b0;
  assign commit_instr_o[111] = (N856)? mem_q[111] : 
                               (N858)? mem_q[474] : 
                               (N860)? mem_q[837] : 
                               (N862)? mem_q[1200] : 
                               (N857)? mem_q[1563] : 
                               (N859)? mem_q[1926] : 
                               (N861)? mem_q[2289] : 
                               (N863)? mem_q[2652] : 1'b0;
  assign commit_instr_o[110] = (N856)? mem_q[110] : 
                               (N858)? mem_q[473] : 
                               (N860)? mem_q[836] : 
                               (N862)? mem_q[1199] : 
                               (N857)? mem_q[1562] : 
                               (N859)? mem_q[1925] : 
                               (N861)? mem_q[2288] : 
                               (N863)? mem_q[2651] : 1'b0;
  assign commit_instr_o[109] = (N856)? mem_q[109] : 
                               (N858)? mem_q[472] : 
                               (N860)? mem_q[835] : 
                               (N862)? mem_q[1198] : 
                               (N857)? mem_q[1561] : 
                               (N859)? mem_q[1924] : 
                               (N861)? mem_q[2287] : 
                               (N863)? mem_q[2650] : 1'b0;
  assign commit_instr_o[108] = (N856)? mem_q[108] : 
                               (N858)? mem_q[471] : 
                               (N860)? mem_q[834] : 
                               (N862)? mem_q[1197] : 
                               (N857)? mem_q[1560] : 
                               (N859)? mem_q[1923] : 
                               (N861)? mem_q[2286] : 
                               (N863)? mem_q[2649] : 1'b0;
  assign commit_instr_o[107] = (N856)? mem_q[107] : 
                               (N858)? mem_q[470] : 
                               (N860)? mem_q[833] : 
                               (N862)? mem_q[1196] : 
                               (N857)? mem_q[1559] : 
                               (N859)? mem_q[1922] : 
                               (N861)? mem_q[2285] : 
                               (N863)? mem_q[2648] : 1'b0;
  assign commit_instr_o[106] = (N856)? mem_q[106] : 
                               (N858)? mem_q[469] : 
                               (N860)? mem_q[832] : 
                               (N862)? mem_q[1195] : 
                               (N857)? mem_q[1558] : 
                               (N859)? mem_q[1921] : 
                               (N861)? mem_q[2284] : 
                               (N863)? mem_q[2647] : 1'b0;
  assign commit_instr_o[105] = (N856)? mem_q[105] : 
                               (N858)? mem_q[468] : 
                               (N860)? mem_q[831] : 
                               (N862)? mem_q[1194] : 
                               (N857)? mem_q[1557] : 
                               (N859)? mem_q[1920] : 
                               (N861)? mem_q[2283] : 
                               (N863)? mem_q[2646] : 1'b0;
  assign commit_instr_o[104] = (N856)? mem_q[104] : 
                               (N858)? mem_q[467] : 
                               (N860)? mem_q[830] : 
                               (N862)? mem_q[1193] : 
                               (N857)? mem_q[1556] : 
                               (N859)? mem_q[1919] : 
                               (N861)? mem_q[2282] : 
                               (N863)? mem_q[2645] : 1'b0;
  assign commit_instr_o[103] = (N856)? mem_q[103] : 
                               (N858)? mem_q[466] : 
                               (N860)? mem_q[829] : 
                               (N862)? mem_q[1192] : 
                               (N857)? mem_q[1555] : 
                               (N859)? mem_q[1918] : 
                               (N861)? mem_q[2281] : 
                               (N863)? mem_q[2644] : 1'b0;
  assign commit_instr_o[102] = (N856)? mem_q[102] : 
                               (N858)? mem_q[465] : 
                               (N860)? mem_q[828] : 
                               (N862)? mem_q[1191] : 
                               (N857)? mem_q[1554] : 
                               (N859)? mem_q[1917] : 
                               (N861)? mem_q[2280] : 
                               (N863)? mem_q[2643] : 1'b0;
  assign commit_instr_o[101] = (N856)? mem_q[101] : 
                               (N858)? mem_q[464] : 
                               (N860)? mem_q[827] : 
                               (N862)? mem_q[1190] : 
                               (N857)? mem_q[1553] : 
                               (N859)? mem_q[1916] : 
                               (N861)? mem_q[2279] : 
                               (N863)? mem_q[2642] : 1'b0;
  assign commit_instr_o[100] = (N856)? mem_q[100] : 
                               (N858)? mem_q[463] : 
                               (N860)? mem_q[826] : 
                               (N862)? mem_q[1189] : 
                               (N857)? mem_q[1552] : 
                               (N859)? mem_q[1915] : 
                               (N861)? mem_q[2278] : 
                               (N863)? mem_q[2641] : 1'b0;
  assign commit_instr_o[99] = (N856)? mem_q[99] : 
                              (N858)? mem_q[462] : 
                              (N860)? mem_q[825] : 
                              (N862)? mem_q[1188] : 
                              (N857)? mem_q[1551] : 
                              (N859)? mem_q[1914] : 
                              (N861)? mem_q[2277] : 
                              (N863)? mem_q[2640] : 1'b0;
  assign commit_instr_o[98] = (N856)? mem_q[98] : 
                              (N858)? mem_q[461] : 
                              (N860)? mem_q[824] : 
                              (N862)? mem_q[1187] : 
                              (N857)? mem_q[1550] : 
                              (N859)? mem_q[1913] : 
                              (N861)? mem_q[2276] : 
                              (N863)? mem_q[2639] : 1'b0;
  assign commit_instr_o[97] = (N856)? mem_q[97] : 
                              (N858)? mem_q[460] : 
                              (N860)? mem_q[823] : 
                              (N862)? mem_q[1186] : 
                              (N857)? mem_q[1549] : 
                              (N859)? mem_q[1912] : 
                              (N861)? mem_q[2275] : 
                              (N863)? mem_q[2638] : 1'b0;
  assign commit_instr_o[96] = (N856)? mem_q[96] : 
                              (N858)? mem_q[459] : 
                              (N860)? mem_q[822] : 
                              (N862)? mem_q[1185] : 
                              (N857)? mem_q[1548] : 
                              (N859)? mem_q[1911] : 
                              (N861)? mem_q[2274] : 
                              (N863)? mem_q[2637] : 1'b0;
  assign commit_instr_o[95] = (N856)? mem_q[95] : 
                              (N858)? mem_q[458] : 
                              (N860)? mem_q[821] : 
                              (N862)? mem_q[1184] : 
                              (N857)? mem_q[1547] : 
                              (N859)? mem_q[1910] : 
                              (N861)? mem_q[2273] : 
                              (N863)? mem_q[2636] : 1'b0;
  assign commit_instr_o[94] = (N856)? mem_q[94] : 
                              (N858)? mem_q[457] : 
                              (N860)? mem_q[820] : 
                              (N862)? mem_q[1183] : 
                              (N857)? mem_q[1546] : 
                              (N859)? mem_q[1909] : 
                              (N861)? mem_q[2272] : 
                              (N863)? mem_q[2635] : 1'b0;
  assign commit_instr_o[93] = (N856)? mem_q[93] : 
                              (N858)? mem_q[456] : 
                              (N860)? mem_q[819] : 
                              (N862)? mem_q[1182] : 
                              (N857)? mem_q[1545] : 
                              (N859)? mem_q[1908] : 
                              (N861)? mem_q[2271] : 
                              (N863)? mem_q[2634] : 1'b0;
  assign commit_instr_o[92] = (N856)? mem_q[92] : 
                              (N858)? mem_q[455] : 
                              (N860)? mem_q[818] : 
                              (N862)? mem_q[1181] : 
                              (N857)? mem_q[1544] : 
                              (N859)? mem_q[1907] : 
                              (N861)? mem_q[2270] : 
                              (N863)? mem_q[2633] : 1'b0;
  assign commit_instr_o[91] = (N856)? mem_q[91] : 
                              (N858)? mem_q[454] : 
                              (N860)? mem_q[817] : 
                              (N862)? mem_q[1180] : 
                              (N857)? mem_q[1543] : 
                              (N859)? mem_q[1906] : 
                              (N861)? mem_q[2269] : 
                              (N863)? mem_q[2632] : 1'b0;
  assign commit_instr_o[90] = (N856)? mem_q[90] : 
                              (N858)? mem_q[453] : 
                              (N860)? mem_q[816] : 
                              (N862)? mem_q[1179] : 
                              (N857)? mem_q[1542] : 
                              (N859)? mem_q[1905] : 
                              (N861)? mem_q[2268] : 
                              (N863)? mem_q[2631] : 1'b0;
  assign commit_instr_o[89] = (N856)? mem_q[89] : 
                              (N858)? mem_q[452] : 
                              (N860)? mem_q[815] : 
                              (N862)? mem_q[1178] : 
                              (N857)? mem_q[1541] : 
                              (N859)? mem_q[1904] : 
                              (N861)? mem_q[2267] : 
                              (N863)? mem_q[2630] : 1'b0;
  assign commit_instr_o[88] = (N856)? mem_q[88] : 
                              (N858)? mem_q[451] : 
                              (N860)? mem_q[814] : 
                              (N862)? mem_q[1177] : 
                              (N857)? mem_q[1540] : 
                              (N859)? mem_q[1903] : 
                              (N861)? mem_q[2266] : 
                              (N863)? mem_q[2629] : 1'b0;
  assign commit_instr_o[87] = (N856)? mem_q[87] : 
                              (N858)? mem_q[450] : 
                              (N860)? mem_q[813] : 
                              (N862)? mem_q[1176] : 
                              (N857)? mem_q[1539] : 
                              (N859)? mem_q[1902] : 
                              (N861)? mem_q[2265] : 
                              (N863)? mem_q[2628] : 1'b0;
  assign commit_instr_o[86] = (N856)? mem_q[86] : 
                              (N858)? mem_q[449] : 
                              (N860)? mem_q[812] : 
                              (N862)? mem_q[1175] : 
                              (N857)? mem_q[1538] : 
                              (N859)? mem_q[1901] : 
                              (N861)? mem_q[2264] : 
                              (N863)? mem_q[2627] : 1'b0;
  assign commit_instr_o[85] = (N856)? mem_q[85] : 
                              (N858)? mem_q[448] : 
                              (N860)? mem_q[811] : 
                              (N862)? mem_q[1174] : 
                              (N857)? mem_q[1537] : 
                              (N859)? mem_q[1900] : 
                              (N861)? mem_q[2263] : 
                              (N863)? mem_q[2626] : 1'b0;
  assign commit_instr_o[84] = (N856)? mem_q[84] : 
                              (N858)? mem_q[447] : 
                              (N860)? mem_q[810] : 
                              (N862)? mem_q[1173] : 
                              (N857)? mem_q[1536] : 
                              (N859)? mem_q[1899] : 
                              (N861)? mem_q[2262] : 
                              (N863)? mem_q[2625] : 1'b0;
  assign commit_instr_o[83] = (N856)? mem_q[83] : 
                              (N858)? mem_q[446] : 
                              (N860)? mem_q[809] : 
                              (N862)? mem_q[1172] : 
                              (N857)? mem_q[1535] : 
                              (N859)? mem_q[1898] : 
                              (N861)? mem_q[2261] : 
                              (N863)? mem_q[2624] : 1'b0;
  assign commit_instr_o[82] = (N856)? mem_q[82] : 
                              (N858)? mem_q[445] : 
                              (N860)? mem_q[808] : 
                              (N862)? mem_q[1171] : 
                              (N857)? mem_q[1534] : 
                              (N859)? mem_q[1897] : 
                              (N861)? mem_q[2260] : 
                              (N863)? mem_q[2623] : 1'b0;
  assign commit_instr_o[81] = (N856)? mem_q[81] : 
                              (N858)? mem_q[444] : 
                              (N860)? mem_q[807] : 
                              (N862)? mem_q[1170] : 
                              (N857)? mem_q[1533] : 
                              (N859)? mem_q[1896] : 
                              (N861)? mem_q[2259] : 
                              (N863)? mem_q[2622] : 1'b0;
  assign commit_instr_o[80] = (N856)? mem_q[80] : 
                              (N858)? mem_q[443] : 
                              (N860)? mem_q[806] : 
                              (N862)? mem_q[1169] : 
                              (N857)? mem_q[1532] : 
                              (N859)? mem_q[1895] : 
                              (N861)? mem_q[2258] : 
                              (N863)? mem_q[2621] : 1'b0;
  assign commit_instr_o[79] = (N856)? mem_q[79] : 
                              (N858)? mem_q[442] : 
                              (N860)? mem_q[805] : 
                              (N862)? mem_q[1168] : 
                              (N857)? mem_q[1531] : 
                              (N859)? mem_q[1894] : 
                              (N861)? mem_q[2257] : 
                              (N863)? mem_q[2620] : 1'b0;
  assign commit_instr_o[78] = (N856)? mem_q[78] : 
                              (N858)? mem_q[441] : 
                              (N860)? mem_q[804] : 
                              (N862)? mem_q[1167] : 
                              (N857)? mem_q[1530] : 
                              (N859)? mem_q[1893] : 
                              (N861)? mem_q[2256] : 
                              (N863)? mem_q[2619] : 1'b0;
  assign commit_instr_o[77] = (N856)? mem_q[77] : 
                              (N858)? mem_q[440] : 
                              (N860)? mem_q[803] : 
                              (N862)? mem_q[1166] : 
                              (N857)? mem_q[1529] : 
                              (N859)? mem_q[1892] : 
                              (N861)? mem_q[2255] : 
                              (N863)? mem_q[2618] : 1'b0;
  assign commit_instr_o[76] = (N856)? mem_q[76] : 
                              (N858)? mem_q[439] : 
                              (N860)? mem_q[802] : 
                              (N862)? mem_q[1165] : 
                              (N857)? mem_q[1528] : 
                              (N859)? mem_q[1891] : 
                              (N861)? mem_q[2254] : 
                              (N863)? mem_q[2617] : 1'b0;
  assign commit_instr_o[75] = (N856)? mem_q[75] : 
                              (N858)? mem_q[438] : 
                              (N860)? mem_q[801] : 
                              (N862)? mem_q[1164] : 
                              (N857)? mem_q[1527] : 
                              (N859)? mem_q[1890] : 
                              (N861)? mem_q[2253] : 
                              (N863)? mem_q[2616] : 1'b0;
  assign commit_instr_o[74] = (N856)? mem_q[74] : 
                              (N858)? mem_q[437] : 
                              (N860)? mem_q[800] : 
                              (N862)? mem_q[1163] : 
                              (N857)? mem_q[1526] : 
                              (N859)? mem_q[1889] : 
                              (N861)? mem_q[2252] : 
                              (N863)? mem_q[2615] : 1'b0;
  assign commit_instr_o[73] = (N856)? mem_q[73] : 
                              (N858)? mem_q[436] : 
                              (N860)? mem_q[799] : 
                              (N862)? mem_q[1162] : 
                              (N857)? mem_q[1525] : 
                              (N859)? mem_q[1888] : 
                              (N861)? mem_q[2251] : 
                              (N863)? mem_q[2614] : 1'b0;
  assign commit_instr_o[72] = (N856)? mem_q[72] : 
                              (N858)? mem_q[435] : 
                              (N860)? mem_q[798] : 
                              (N862)? mem_q[1161] : 
                              (N857)? mem_q[1524] : 
                              (N859)? mem_q[1887] : 
                              (N861)? mem_q[2250] : 
                              (N863)? mem_q[2613] : 1'b0;
  assign commit_instr_o[71] = (N856)? mem_q[71] : 
                              (N858)? mem_q[434] : 
                              (N860)? mem_q[797] : 
                              (N862)? mem_q[1160] : 
                              (N857)? mem_q[1523] : 
                              (N859)? mem_q[1886] : 
                              (N861)? mem_q[2249] : 
                              (N863)? mem_q[2612] : 1'b0;
  assign commit_instr_o[70] = (N856)? mem_q[70] : 
                              (N858)? mem_q[433] : 
                              (N860)? mem_q[796] : 
                              (N862)? mem_q[1159] : 
                              (N857)? mem_q[1522] : 
                              (N859)? mem_q[1885] : 
                              (N861)? mem_q[2248] : 
                              (N863)? mem_q[2611] : 1'b0;
  assign commit_instr_o[69] = (N856)? mem_q[69] : 
                              (N858)? mem_q[432] : 
                              (N860)? mem_q[795] : 
                              (N862)? mem_q[1158] : 
                              (N857)? mem_q[1521] : 
                              (N859)? mem_q[1884] : 
                              (N861)? mem_q[2247] : 
                              (N863)? mem_q[2610] : 1'b0;
  assign commit_instr_o[68] = (N856)? mem_q[68] : 
                              (N858)? mem_q[431] : 
                              (N860)? mem_q[794] : 
                              (N862)? mem_q[1157] : 
                              (N857)? mem_q[1520] : 
                              (N859)? mem_q[1883] : 
                              (N861)? mem_q[2246] : 
                              (N863)? mem_q[2609] : 1'b0;
  assign commit_instr_o[67] = (N856)? mem_q[67] : 
                              (N858)? mem_q[430] : 
                              (N860)? mem_q[793] : 
                              (N862)? mem_q[1156] : 
                              (N857)? mem_q[1519] : 
                              (N859)? mem_q[1882] : 
                              (N861)? mem_q[2245] : 
                              (N863)? mem_q[2608] : 1'b0;
  assign commit_instr_o[66] = (N856)? mem_q[66] : 
                              (N858)? mem_q[429] : 
                              (N860)? mem_q[792] : 
                              (N862)? mem_q[1155] : 
                              (N857)? mem_q[1518] : 
                              (N859)? mem_q[1881] : 
                              (N861)? mem_q[2244] : 
                              (N863)? mem_q[2607] : 1'b0;
  assign commit_instr_o[65] = (N856)? mem_q[65] : 
                              (N858)? mem_q[428] : 
                              (N860)? mem_q[791] : 
                              (N862)? mem_q[1154] : 
                              (N857)? mem_q[1517] : 
                              (N859)? mem_q[1880] : 
                              (N861)? mem_q[2243] : 
                              (N863)? mem_q[2606] : 1'b0;
  assign commit_instr_o[64] = (N856)? mem_q[64] : 
                              (N858)? mem_q[427] : 
                              (N860)? mem_q[790] : 
                              (N862)? mem_q[1153] : 
                              (N857)? mem_q[1516] : 
                              (N859)? mem_q[1879] : 
                              (N861)? mem_q[2242] : 
                              (N863)? mem_q[2605] : 1'b0;
  assign commit_instr_o[63] = (N856)? mem_q[63] : 
                              (N858)? mem_q[426] : 
                              (N860)? mem_q[789] : 
                              (N862)? mem_q[1152] : 
                              (N857)? mem_q[1515] : 
                              (N859)? mem_q[1878] : 
                              (N861)? mem_q[2241] : 
                              (N863)? mem_q[2604] : 1'b0;
  assign commit_instr_o[62] = (N856)? mem_q[62] : 
                              (N858)? mem_q[425] : 
                              (N860)? mem_q[788] : 
                              (N862)? mem_q[1151] : 
                              (N857)? mem_q[1514] : 
                              (N859)? mem_q[1877] : 
                              (N861)? mem_q[2240] : 
                              (N863)? mem_q[2603] : 1'b0;
  assign commit_instr_o[61] = (N856)? mem_q[61] : 
                              (N858)? mem_q[424] : 
                              (N860)? mem_q[787] : 
                              (N862)? mem_q[1150] : 
                              (N857)? mem_q[1513] : 
                              (N859)? mem_q[1876] : 
                              (N861)? mem_q[2239] : 
                              (N863)? mem_q[2602] : 1'b0;
  assign commit_instr_o[60] = (N856)? mem_q[60] : 
                              (N858)? mem_q[423] : 
                              (N860)? mem_q[786] : 
                              (N862)? mem_q[1149] : 
                              (N857)? mem_q[1512] : 
                              (N859)? mem_q[1875] : 
                              (N861)? mem_q[2238] : 
                              (N863)? mem_q[2601] : 1'b0;
  assign commit_instr_o[59] = (N856)? mem_q[59] : 
                              (N858)? mem_q[422] : 
                              (N860)? mem_q[785] : 
                              (N862)? mem_q[1148] : 
                              (N857)? mem_q[1511] : 
                              (N859)? mem_q[1874] : 
                              (N861)? mem_q[2237] : 
                              (N863)? mem_q[2600] : 1'b0;
  assign commit_instr_o[58] = (N856)? mem_q[58] : 
                              (N858)? mem_q[421] : 
                              (N860)? mem_q[784] : 
                              (N862)? mem_q[1147] : 
                              (N857)? mem_q[1510] : 
                              (N859)? mem_q[1873] : 
                              (N861)? mem_q[2236] : 
                              (N863)? mem_q[2599] : 1'b0;
  assign commit_instr_o[57] = (N856)? mem_q[57] : 
                              (N858)? mem_q[420] : 
                              (N860)? mem_q[783] : 
                              (N862)? mem_q[1146] : 
                              (N857)? mem_q[1509] : 
                              (N859)? mem_q[1872] : 
                              (N861)? mem_q[2235] : 
                              (N863)? mem_q[2598] : 1'b0;
  assign commit_instr_o[56] = (N856)? mem_q[56] : 
                              (N858)? mem_q[419] : 
                              (N860)? mem_q[782] : 
                              (N862)? mem_q[1145] : 
                              (N857)? mem_q[1508] : 
                              (N859)? mem_q[1871] : 
                              (N861)? mem_q[2234] : 
                              (N863)? mem_q[2597] : 1'b0;
  assign commit_instr_o[55] = (N856)? mem_q[55] : 
                              (N858)? mem_q[418] : 
                              (N860)? mem_q[781] : 
                              (N862)? mem_q[1144] : 
                              (N857)? mem_q[1507] : 
                              (N859)? mem_q[1870] : 
                              (N861)? mem_q[2233] : 
                              (N863)? mem_q[2596] : 1'b0;
  assign commit_instr_o[54] = (N856)? mem_q[54] : 
                              (N858)? mem_q[417] : 
                              (N860)? mem_q[780] : 
                              (N862)? mem_q[1143] : 
                              (N857)? mem_q[1506] : 
                              (N859)? mem_q[1869] : 
                              (N861)? mem_q[2232] : 
                              (N863)? mem_q[2595] : 1'b0;
  assign commit_instr_o[53] = (N856)? mem_q[53] : 
                              (N858)? mem_q[416] : 
                              (N860)? mem_q[779] : 
                              (N862)? mem_q[1142] : 
                              (N857)? mem_q[1505] : 
                              (N859)? mem_q[1868] : 
                              (N861)? mem_q[2231] : 
                              (N863)? mem_q[2594] : 1'b0;
  assign commit_instr_o[52] = (N856)? mem_q[52] : 
                              (N858)? mem_q[415] : 
                              (N860)? mem_q[778] : 
                              (N862)? mem_q[1141] : 
                              (N857)? mem_q[1504] : 
                              (N859)? mem_q[1867] : 
                              (N861)? mem_q[2230] : 
                              (N863)? mem_q[2593] : 1'b0;
  assign commit_instr_o[51] = (N856)? mem_q[51] : 
                              (N858)? mem_q[414] : 
                              (N860)? mem_q[777] : 
                              (N862)? mem_q[1140] : 
                              (N857)? mem_q[1503] : 
                              (N859)? mem_q[1866] : 
                              (N861)? mem_q[2229] : 
                              (N863)? mem_q[2592] : 1'b0;
  assign commit_instr_o[50] = (N856)? mem_q[50] : 
                              (N858)? mem_q[413] : 
                              (N860)? mem_q[776] : 
                              (N862)? mem_q[1139] : 
                              (N857)? mem_q[1502] : 
                              (N859)? mem_q[1865] : 
                              (N861)? mem_q[2228] : 
                              (N863)? mem_q[2591] : 1'b0;
  assign commit_instr_o[49] = (N856)? mem_q[49] : 
                              (N858)? mem_q[412] : 
                              (N860)? mem_q[775] : 
                              (N862)? mem_q[1138] : 
                              (N857)? mem_q[1501] : 
                              (N859)? mem_q[1864] : 
                              (N861)? mem_q[2227] : 
                              (N863)? mem_q[2590] : 1'b0;
  assign commit_instr_o[48] = (N856)? mem_q[48] : 
                              (N858)? mem_q[411] : 
                              (N860)? mem_q[774] : 
                              (N862)? mem_q[1137] : 
                              (N857)? mem_q[1500] : 
                              (N859)? mem_q[1863] : 
                              (N861)? mem_q[2226] : 
                              (N863)? mem_q[2589] : 1'b0;
  assign commit_instr_o[47] = (N856)? mem_q[47] : 
                              (N858)? mem_q[410] : 
                              (N860)? mem_q[773] : 
                              (N862)? mem_q[1136] : 
                              (N857)? mem_q[1499] : 
                              (N859)? mem_q[1862] : 
                              (N861)? mem_q[2225] : 
                              (N863)? mem_q[2588] : 1'b0;
  assign commit_instr_o[46] = (N856)? mem_q[46] : 
                              (N858)? mem_q[409] : 
                              (N860)? mem_q[772] : 
                              (N862)? mem_q[1135] : 
                              (N857)? mem_q[1498] : 
                              (N859)? mem_q[1861] : 
                              (N861)? mem_q[2224] : 
                              (N863)? mem_q[2587] : 1'b0;
  assign commit_instr_o[45] = (N856)? mem_q[45] : 
                              (N858)? mem_q[408] : 
                              (N860)? mem_q[771] : 
                              (N862)? mem_q[1134] : 
                              (N857)? mem_q[1497] : 
                              (N859)? mem_q[1860] : 
                              (N861)? mem_q[2223] : 
                              (N863)? mem_q[2586] : 1'b0;
  assign commit_instr_o[44] = (N856)? mem_q[44] : 
                              (N858)? mem_q[407] : 
                              (N860)? mem_q[770] : 
                              (N862)? mem_q[1133] : 
                              (N857)? mem_q[1496] : 
                              (N859)? mem_q[1859] : 
                              (N861)? mem_q[2222] : 
                              (N863)? mem_q[2585] : 1'b0;
  assign commit_instr_o[43] = (N856)? mem_q[43] : 
                              (N858)? mem_q[406] : 
                              (N860)? mem_q[769] : 
                              (N862)? mem_q[1132] : 
                              (N857)? mem_q[1495] : 
                              (N859)? mem_q[1858] : 
                              (N861)? mem_q[2221] : 
                              (N863)? mem_q[2584] : 1'b0;
  assign commit_instr_o[42] = (N856)? mem_q[42] : 
                              (N858)? mem_q[405] : 
                              (N860)? mem_q[768] : 
                              (N862)? mem_q[1131] : 
                              (N857)? mem_q[1494] : 
                              (N859)? mem_q[1857] : 
                              (N861)? mem_q[2220] : 
                              (N863)? mem_q[2583] : 1'b0;
  assign commit_instr_o[41] = (N856)? mem_q[41] : 
                              (N858)? mem_q[404] : 
                              (N860)? mem_q[767] : 
                              (N862)? mem_q[1130] : 
                              (N857)? mem_q[1493] : 
                              (N859)? mem_q[1856] : 
                              (N861)? mem_q[2219] : 
                              (N863)? mem_q[2582] : 1'b0;
  assign commit_instr_o[40] = (N856)? mem_q[40] : 
                              (N858)? mem_q[403] : 
                              (N860)? mem_q[766] : 
                              (N862)? mem_q[1129] : 
                              (N857)? mem_q[1492] : 
                              (N859)? mem_q[1855] : 
                              (N861)? mem_q[2218] : 
                              (N863)? mem_q[2581] : 1'b0;
  assign commit_instr_o[39] = (N856)? mem_q[39] : 
                              (N858)? mem_q[402] : 
                              (N860)? mem_q[765] : 
                              (N862)? mem_q[1128] : 
                              (N857)? mem_q[1491] : 
                              (N859)? mem_q[1854] : 
                              (N861)? mem_q[2217] : 
                              (N863)? mem_q[2580] : 1'b0;
  assign commit_instr_o[38] = (N856)? mem_q[38] : 
                              (N858)? mem_q[401] : 
                              (N860)? mem_q[764] : 
                              (N862)? mem_q[1127] : 
                              (N857)? mem_q[1490] : 
                              (N859)? mem_q[1853] : 
                              (N861)? mem_q[2216] : 
                              (N863)? mem_q[2579] : 1'b0;
  assign commit_instr_o[37] = (N856)? mem_q[37] : 
                              (N858)? mem_q[400] : 
                              (N860)? mem_q[763] : 
                              (N862)? mem_q[1126] : 
                              (N857)? mem_q[1489] : 
                              (N859)? mem_q[1852] : 
                              (N861)? mem_q[2215] : 
                              (N863)? mem_q[2578] : 1'b0;
  assign commit_instr_o[36] = (N856)? mem_q[36] : 
                              (N858)? mem_q[399] : 
                              (N860)? mem_q[762] : 
                              (N862)? mem_q[1125] : 
                              (N857)? mem_q[1488] : 
                              (N859)? mem_q[1851] : 
                              (N861)? mem_q[2214] : 
                              (N863)? mem_q[2577] : 1'b0;
  assign commit_instr_o[35] = (N856)? mem_q[35] : 
                              (N858)? mem_q[398] : 
                              (N860)? mem_q[761] : 
                              (N862)? mem_q[1124] : 
                              (N857)? mem_q[1487] : 
                              (N859)? mem_q[1850] : 
                              (N861)? mem_q[2213] : 
                              (N863)? mem_q[2576] : 1'b0;
  assign commit_instr_o[34] = (N856)? mem_q[34] : 
                              (N858)? mem_q[397] : 
                              (N860)? mem_q[760] : 
                              (N862)? mem_q[1123] : 
                              (N857)? mem_q[1486] : 
                              (N859)? mem_q[1849] : 
                              (N861)? mem_q[2212] : 
                              (N863)? mem_q[2575] : 1'b0;
  assign commit_instr_o[33] = (N856)? mem_q[33] : 
                              (N858)? mem_q[396] : 
                              (N860)? mem_q[759] : 
                              (N862)? mem_q[1122] : 
                              (N857)? mem_q[1485] : 
                              (N859)? mem_q[1848] : 
                              (N861)? mem_q[2211] : 
                              (N863)? mem_q[2574] : 1'b0;
  assign commit_instr_o[32] = (N856)? mem_q[32] : 
                              (N858)? mem_q[395] : 
                              (N860)? mem_q[758] : 
                              (N862)? mem_q[1121] : 
                              (N857)? mem_q[1484] : 
                              (N859)? mem_q[1847] : 
                              (N861)? mem_q[2210] : 
                              (N863)? mem_q[2573] : 1'b0;
  assign commit_instr_o[31] = (N856)? mem_q[31] : 
                              (N858)? mem_q[394] : 
                              (N860)? mem_q[757] : 
                              (N862)? mem_q[1120] : 
                              (N857)? mem_q[1483] : 
                              (N859)? mem_q[1846] : 
                              (N861)? mem_q[2209] : 
                              (N863)? mem_q[2572] : 1'b0;
  assign commit_instr_o[30] = (N856)? mem_q[30] : 
                              (N858)? mem_q[393] : 
                              (N860)? mem_q[756] : 
                              (N862)? mem_q[1119] : 
                              (N857)? mem_q[1482] : 
                              (N859)? mem_q[1845] : 
                              (N861)? mem_q[2208] : 
                              (N863)? mem_q[2571] : 1'b0;
  assign commit_instr_o[29] = (N856)? mem_q[29] : 
                              (N858)? mem_q[392] : 
                              (N860)? mem_q[755] : 
                              (N862)? mem_q[1118] : 
                              (N857)? mem_q[1481] : 
                              (N859)? mem_q[1844] : 
                              (N861)? mem_q[2207] : 
                              (N863)? mem_q[2570] : 1'b0;
  assign commit_instr_o[28] = (N856)? mem_q[28] : 
                              (N858)? mem_q[391] : 
                              (N860)? mem_q[754] : 
                              (N862)? mem_q[1117] : 
                              (N857)? mem_q[1480] : 
                              (N859)? mem_q[1843] : 
                              (N861)? mem_q[2206] : 
                              (N863)? mem_q[2569] : 1'b0;
  assign commit_instr_o[27] = (N856)? mem_q[27] : 
                              (N858)? mem_q[390] : 
                              (N860)? mem_q[753] : 
                              (N862)? mem_q[1116] : 
                              (N857)? mem_q[1479] : 
                              (N859)? mem_q[1842] : 
                              (N861)? mem_q[2205] : 
                              (N863)? mem_q[2568] : 1'b0;
  assign commit_instr_o[26] = (N856)? mem_q[26] : 
                              (N858)? mem_q[389] : 
                              (N860)? mem_q[752] : 
                              (N862)? mem_q[1115] : 
                              (N857)? mem_q[1478] : 
                              (N859)? mem_q[1841] : 
                              (N861)? mem_q[2204] : 
                              (N863)? mem_q[2567] : 1'b0;
  assign commit_instr_o[25] = (N856)? mem_q[25] : 
                              (N858)? mem_q[388] : 
                              (N860)? mem_q[751] : 
                              (N862)? mem_q[1114] : 
                              (N857)? mem_q[1477] : 
                              (N859)? mem_q[1840] : 
                              (N861)? mem_q[2203] : 
                              (N863)? mem_q[2566] : 1'b0;
  assign commit_instr_o[24] = (N856)? mem_q[24] : 
                              (N858)? mem_q[387] : 
                              (N860)? mem_q[750] : 
                              (N862)? mem_q[1113] : 
                              (N857)? mem_q[1476] : 
                              (N859)? mem_q[1839] : 
                              (N861)? mem_q[2202] : 
                              (N863)? mem_q[2565] : 1'b0;
  assign commit_instr_o[23] = (N856)? mem_q[23] : 
                              (N858)? mem_q[386] : 
                              (N860)? mem_q[749] : 
                              (N862)? mem_q[1112] : 
                              (N857)? mem_q[1475] : 
                              (N859)? mem_q[1838] : 
                              (N861)? mem_q[2201] : 
                              (N863)? mem_q[2564] : 1'b0;
  assign commit_instr_o[22] = (N856)? mem_q[22] : 
                              (N858)? mem_q[385] : 
                              (N860)? mem_q[748] : 
                              (N862)? mem_q[1111] : 
                              (N857)? mem_q[1474] : 
                              (N859)? mem_q[1837] : 
                              (N861)? mem_q[2200] : 
                              (N863)? mem_q[2563] : 1'b0;
  assign commit_instr_o[21] = (N856)? mem_q[21] : 
                              (N858)? mem_q[384] : 
                              (N860)? mem_q[747] : 
                              (N862)? mem_q[1110] : 
                              (N857)? mem_q[1473] : 
                              (N859)? mem_q[1836] : 
                              (N861)? mem_q[2199] : 
                              (N863)? mem_q[2562] : 1'b0;
  assign commit_instr_o[20] = (N856)? mem_q[20] : 
                              (N858)? mem_q[383] : 
                              (N860)? mem_q[746] : 
                              (N862)? mem_q[1109] : 
                              (N857)? mem_q[1472] : 
                              (N859)? mem_q[1835] : 
                              (N861)? mem_q[2198] : 
                              (N863)? mem_q[2561] : 1'b0;
  assign commit_instr_o[19] = (N856)? mem_q[19] : 
                              (N858)? mem_q[382] : 
                              (N860)? mem_q[745] : 
                              (N862)? mem_q[1108] : 
                              (N857)? mem_q[1471] : 
                              (N859)? mem_q[1834] : 
                              (N861)? mem_q[2197] : 
                              (N863)? mem_q[2560] : 1'b0;
  assign commit_instr_o[18] = (N856)? mem_q[18] : 
                              (N858)? mem_q[381] : 
                              (N860)? mem_q[744] : 
                              (N862)? mem_q[1107] : 
                              (N857)? mem_q[1470] : 
                              (N859)? mem_q[1833] : 
                              (N861)? mem_q[2196] : 
                              (N863)? mem_q[2559] : 1'b0;
  assign commit_instr_o[17] = (N856)? mem_q[17] : 
                              (N858)? mem_q[380] : 
                              (N860)? mem_q[743] : 
                              (N862)? mem_q[1106] : 
                              (N857)? mem_q[1469] : 
                              (N859)? mem_q[1832] : 
                              (N861)? mem_q[2195] : 
                              (N863)? mem_q[2558] : 1'b0;
  assign commit_instr_o[16] = (N856)? mem_q[16] : 
                              (N858)? mem_q[379] : 
                              (N860)? mem_q[742] : 
                              (N862)? mem_q[1105] : 
                              (N857)? mem_q[1468] : 
                              (N859)? mem_q[1831] : 
                              (N861)? mem_q[2194] : 
                              (N863)? mem_q[2557] : 1'b0;
  assign commit_instr_o[15] = (N856)? mem_q[15] : 
                              (N858)? mem_q[378] : 
                              (N860)? mem_q[741] : 
                              (N862)? mem_q[1104] : 
                              (N857)? mem_q[1467] : 
                              (N859)? mem_q[1830] : 
                              (N861)? mem_q[2193] : 
                              (N863)? mem_q[2556] : 1'b0;
  assign commit_instr_o[14] = (N856)? mem_q[14] : 
                              (N858)? mem_q[377] : 
                              (N860)? mem_q[740] : 
                              (N862)? mem_q[1103] : 
                              (N857)? mem_q[1466] : 
                              (N859)? mem_q[1829] : 
                              (N861)? mem_q[2192] : 
                              (N863)? mem_q[2555] : 1'b0;
  assign commit_instr_o[13] = (N856)? mem_q[13] : 
                              (N858)? mem_q[376] : 
                              (N860)? mem_q[739] : 
                              (N862)? mem_q[1102] : 
                              (N857)? mem_q[1465] : 
                              (N859)? mem_q[1828] : 
                              (N861)? mem_q[2191] : 
                              (N863)? mem_q[2554] : 1'b0;
  assign commit_instr_o[12] = (N856)? mem_q[12] : 
                              (N858)? mem_q[375] : 
                              (N860)? mem_q[738] : 
                              (N862)? mem_q[1101] : 
                              (N857)? mem_q[1464] : 
                              (N859)? mem_q[1827] : 
                              (N861)? mem_q[2190] : 
                              (N863)? mem_q[2553] : 1'b0;
  assign commit_instr_o[11] = (N856)? mem_q[11] : 
                              (N858)? mem_q[374] : 
                              (N860)? mem_q[737] : 
                              (N862)? mem_q[1100] : 
                              (N857)? mem_q[1463] : 
                              (N859)? mem_q[1826] : 
                              (N861)? mem_q[2189] : 
                              (N863)? mem_q[2552] : 1'b0;
  assign commit_instr_o[10] = (N856)? mem_q[10] : 
                              (N858)? mem_q[373] : 
                              (N860)? mem_q[736] : 
                              (N862)? mem_q[1099] : 
                              (N857)? mem_q[1462] : 
                              (N859)? mem_q[1825] : 
                              (N861)? mem_q[2188] : 
                              (N863)? mem_q[2551] : 1'b0;
  assign commit_instr_o[9] = (N856)? mem_q[9] : 
                             (N858)? mem_q[372] : 
                             (N860)? mem_q[735] : 
                             (N862)? mem_q[1098] : 
                             (N857)? mem_q[1461] : 
                             (N859)? mem_q[1824] : 
                             (N861)? mem_q[2187] : 
                             (N863)? mem_q[2550] : 1'b0;
  assign commit_instr_o[8] = (N856)? mem_q[8] : 
                             (N858)? mem_q[371] : 
                             (N860)? mem_q[734] : 
                             (N862)? mem_q[1097] : 
                             (N857)? mem_q[1460] : 
                             (N859)? mem_q[1823] : 
                             (N861)? mem_q[2186] : 
                             (N863)? mem_q[2549] : 1'b0;
  assign commit_instr_o[7] = (N856)? mem_q[7] : 
                             (N858)? mem_q[370] : 
                             (N860)? mem_q[733] : 
                             (N862)? mem_q[1096] : 
                             (N857)? mem_q[1459] : 
                             (N859)? mem_q[1822] : 
                             (N861)? mem_q[2185] : 
                             (N863)? mem_q[2548] : 1'b0;
  assign commit_instr_o[6] = (N856)? mem_q[6] : 
                             (N858)? mem_q[369] : 
                             (N860)? mem_q[732] : 
                             (N862)? mem_q[1095] : 
                             (N857)? mem_q[1458] : 
                             (N859)? mem_q[1821] : 
                             (N861)? mem_q[2184] : 
                             (N863)? mem_q[2547] : 1'b0;
  assign commit_instr_o[5] = (N856)? mem_q[5] : 
                             (N858)? mem_q[368] : 
                             (N860)? mem_q[731] : 
                             (N862)? mem_q[1094] : 
                             (N857)? mem_q[1457] : 
                             (N859)? mem_q[1820] : 
                             (N861)? mem_q[2183] : 
                             (N863)? mem_q[2546] : 1'b0;
  assign commit_instr_o[4] = (N856)? mem_q[4] : 
                             (N858)? mem_q[367] : 
                             (N860)? mem_q[730] : 
                             (N862)? mem_q[1093] : 
                             (N857)? mem_q[1456] : 
                             (N859)? mem_q[1819] : 
                             (N861)? mem_q[2182] : 
                             (N863)? mem_q[2545] : 1'b0;
  assign commit_instr_o[3] = (N856)? mem_q[3] : 
                             (N858)? mem_q[366] : 
                             (N860)? mem_q[729] : 
                             (N862)? mem_q[1092] : 
                             (N857)? mem_q[1455] : 
                             (N859)? mem_q[1818] : 
                             (N861)? mem_q[2181] : 
                             (N863)? mem_q[2544] : 1'b0;
  assign commit_instr_o[2] = (N856)? mem_q[2] : 
                             (N858)? mem_q[365] : 
                             (N860)? mem_q[728] : 
                             (N862)? mem_q[1091] : 
                             (N857)? mem_q[1454] : 
                             (N859)? mem_q[1817] : 
                             (N861)? mem_q[2180] : 
                             (N863)? mem_q[2543] : 1'b0;
  assign commit_instr_o[1] = (N856)? mem_q[1] : 
                             (N858)? mem_q[364] : 
                             (N860)? mem_q[727] : 
                             (N862)? mem_q[1090] : 
                             (N857)? mem_q[1453] : 
                             (N859)? mem_q[1816] : 
                             (N861)? mem_q[2179] : 
                             (N863)? mem_q[2542] : 1'b0;
  assign commit_instr_o[0] = (N856)? mem_q[0] : 
                             (N858)? mem_q[363] : 
                             (N860)? mem_q[726] : 
                             (N862)? mem_q[1089] : 
                             (N857)? mem_q[1452] : 
                             (N859)? mem_q[1815] : 
                             (N861)? mem_q[2178] : 
                             (N863)? mem_q[2541] : 1'b0;
  assign commit_instr_o[723] = (N874)? mem_q[361] : 
                               (N876)? mem_q[724] : 
                               (N878)? mem_q[1087] : 
                               (N880)? mem_q[1450] : 
                               (N875)? mem_q[1813] : 
                               (N877)? mem_q[2176] : 
                               (N879)? mem_q[2539] : 
                               (N881)? mem_q[2902] : 1'b0;
  assign commit_instr_o[722] = (N874)? mem_q[360] : 
                               (N876)? mem_q[723] : 
                               (N878)? mem_q[1086] : 
                               (N880)? mem_q[1449] : 
                               (N875)? mem_q[1812] : 
                               (N877)? mem_q[2175] : 
                               (N879)? mem_q[2538] : 
                               (N881)? mem_q[2901] : 1'b0;
  assign commit_instr_o[721] = (N874)? mem_q[359] : 
                               (N876)? mem_q[722] : 
                               (N878)? mem_q[1085] : 
                               (N880)? mem_q[1448] : 
                               (N875)? mem_q[1811] : 
                               (N877)? mem_q[2174] : 
                               (N879)? mem_q[2537] : 
                               (N881)? mem_q[2900] : 1'b0;
  assign commit_instr_o[720] = (N874)? mem_q[358] : 
                               (N876)? mem_q[721] : 
                               (N878)? mem_q[1084] : 
                               (N880)? mem_q[1447] : 
                               (N875)? mem_q[1810] : 
                               (N877)? mem_q[2173] : 
                               (N879)? mem_q[2536] : 
                               (N881)? mem_q[2899] : 1'b0;
  assign commit_instr_o[719] = (N874)? mem_q[357] : 
                               (N876)? mem_q[720] : 
                               (N878)? mem_q[1083] : 
                               (N880)? mem_q[1446] : 
                               (N875)? mem_q[1809] : 
                               (N877)? mem_q[2172] : 
                               (N879)? mem_q[2535] : 
                               (N881)? mem_q[2898] : 1'b0;
  assign commit_instr_o[718] = (N874)? mem_q[356] : 
                               (N876)? mem_q[719] : 
                               (N878)? mem_q[1082] : 
                               (N880)? mem_q[1445] : 
                               (N875)? mem_q[1808] : 
                               (N877)? mem_q[2171] : 
                               (N879)? mem_q[2534] : 
                               (N881)? mem_q[2897] : 1'b0;
  assign commit_instr_o[717] = (N874)? mem_q[355] : 
                               (N876)? mem_q[718] : 
                               (N878)? mem_q[1081] : 
                               (N880)? mem_q[1444] : 
                               (N875)? mem_q[1807] : 
                               (N877)? mem_q[2170] : 
                               (N879)? mem_q[2533] : 
                               (N881)? mem_q[2896] : 1'b0;
  assign commit_instr_o[716] = (N874)? mem_q[354] : 
                               (N876)? mem_q[717] : 
                               (N878)? mem_q[1080] : 
                               (N880)? mem_q[1443] : 
                               (N875)? mem_q[1806] : 
                               (N877)? mem_q[2169] : 
                               (N879)? mem_q[2532] : 
                               (N881)? mem_q[2895] : 1'b0;
  assign commit_instr_o[715] = (N874)? mem_q[353] : 
                               (N876)? mem_q[716] : 
                               (N878)? mem_q[1079] : 
                               (N880)? mem_q[1442] : 
                               (N875)? mem_q[1805] : 
                               (N877)? mem_q[2168] : 
                               (N879)? mem_q[2531] : 
                               (N881)? mem_q[2894] : 1'b0;
  assign commit_instr_o[714] = (N874)? mem_q[352] : 
                               (N876)? mem_q[715] : 
                               (N878)? mem_q[1078] : 
                               (N880)? mem_q[1441] : 
                               (N875)? mem_q[1804] : 
                               (N877)? mem_q[2167] : 
                               (N879)? mem_q[2530] : 
                               (N881)? mem_q[2893] : 1'b0;
  assign commit_instr_o[713] = (N874)? mem_q[351] : 
                               (N876)? mem_q[714] : 
                               (N878)? mem_q[1077] : 
                               (N880)? mem_q[1440] : 
                               (N875)? mem_q[1803] : 
                               (N877)? mem_q[2166] : 
                               (N879)? mem_q[2529] : 
                               (N881)? mem_q[2892] : 1'b0;
  assign commit_instr_o[712] = (N874)? mem_q[350] : 
                               (N876)? mem_q[713] : 
                               (N878)? mem_q[1076] : 
                               (N880)? mem_q[1439] : 
                               (N875)? mem_q[1802] : 
                               (N877)? mem_q[2165] : 
                               (N879)? mem_q[2528] : 
                               (N881)? mem_q[2891] : 1'b0;
  assign commit_instr_o[711] = (N874)? mem_q[349] : 
                               (N876)? mem_q[712] : 
                               (N878)? mem_q[1075] : 
                               (N880)? mem_q[1438] : 
                               (N875)? mem_q[1801] : 
                               (N877)? mem_q[2164] : 
                               (N879)? mem_q[2527] : 
                               (N881)? mem_q[2890] : 1'b0;
  assign commit_instr_o[710] = (N874)? mem_q[348] : 
                               (N876)? mem_q[711] : 
                               (N878)? mem_q[1074] : 
                               (N880)? mem_q[1437] : 
                               (N875)? mem_q[1800] : 
                               (N877)? mem_q[2163] : 
                               (N879)? mem_q[2526] : 
                               (N881)? mem_q[2889] : 1'b0;
  assign commit_instr_o[709] = (N874)? mem_q[347] : 
                               (N876)? mem_q[710] : 
                               (N878)? mem_q[1073] : 
                               (N880)? mem_q[1436] : 
                               (N875)? mem_q[1799] : 
                               (N877)? mem_q[2162] : 
                               (N879)? mem_q[2525] : 
                               (N881)? mem_q[2888] : 1'b0;
  assign commit_instr_o[708] = (N874)? mem_q[346] : 
                               (N876)? mem_q[709] : 
                               (N878)? mem_q[1072] : 
                               (N880)? mem_q[1435] : 
                               (N875)? mem_q[1798] : 
                               (N877)? mem_q[2161] : 
                               (N879)? mem_q[2524] : 
                               (N881)? mem_q[2887] : 1'b0;
  assign commit_instr_o[707] = (N874)? mem_q[345] : 
                               (N876)? mem_q[708] : 
                               (N878)? mem_q[1071] : 
                               (N880)? mem_q[1434] : 
                               (N875)? mem_q[1797] : 
                               (N877)? mem_q[2160] : 
                               (N879)? mem_q[2523] : 
                               (N881)? mem_q[2886] : 1'b0;
  assign commit_instr_o[706] = (N874)? mem_q[344] : 
                               (N876)? mem_q[707] : 
                               (N878)? mem_q[1070] : 
                               (N880)? mem_q[1433] : 
                               (N875)? mem_q[1796] : 
                               (N877)? mem_q[2159] : 
                               (N879)? mem_q[2522] : 
                               (N881)? mem_q[2885] : 1'b0;
  assign commit_instr_o[705] = (N874)? mem_q[343] : 
                               (N876)? mem_q[706] : 
                               (N878)? mem_q[1069] : 
                               (N880)? mem_q[1432] : 
                               (N875)? mem_q[1795] : 
                               (N877)? mem_q[2158] : 
                               (N879)? mem_q[2521] : 
                               (N881)? mem_q[2884] : 1'b0;
  assign commit_instr_o[704] = (N874)? mem_q[342] : 
                               (N876)? mem_q[705] : 
                               (N878)? mem_q[1068] : 
                               (N880)? mem_q[1431] : 
                               (N875)? mem_q[1794] : 
                               (N877)? mem_q[2157] : 
                               (N879)? mem_q[2520] : 
                               (N881)? mem_q[2883] : 1'b0;
  assign commit_instr_o[703] = (N874)? mem_q[341] : 
                               (N876)? mem_q[704] : 
                               (N878)? mem_q[1067] : 
                               (N880)? mem_q[1430] : 
                               (N875)? mem_q[1793] : 
                               (N877)? mem_q[2156] : 
                               (N879)? mem_q[2519] : 
                               (N881)? mem_q[2882] : 1'b0;
  assign commit_instr_o[702] = (N874)? mem_q[340] : 
                               (N876)? mem_q[703] : 
                               (N878)? mem_q[1066] : 
                               (N880)? mem_q[1429] : 
                               (N875)? mem_q[1792] : 
                               (N877)? mem_q[2155] : 
                               (N879)? mem_q[2518] : 
                               (N881)? mem_q[2881] : 1'b0;
  assign commit_instr_o[701] = (N874)? mem_q[339] : 
                               (N876)? mem_q[702] : 
                               (N878)? mem_q[1065] : 
                               (N880)? mem_q[1428] : 
                               (N875)? mem_q[1791] : 
                               (N877)? mem_q[2154] : 
                               (N879)? mem_q[2517] : 
                               (N881)? mem_q[2880] : 1'b0;
  assign commit_instr_o[700] = (N874)? mem_q[338] : 
                               (N876)? mem_q[701] : 
                               (N878)? mem_q[1064] : 
                               (N880)? mem_q[1427] : 
                               (N875)? mem_q[1790] : 
                               (N877)? mem_q[2153] : 
                               (N879)? mem_q[2516] : 
                               (N881)? mem_q[2879] : 1'b0;
  assign commit_instr_o[699] = (N874)? mem_q[337] : 
                               (N876)? mem_q[700] : 
                               (N878)? mem_q[1063] : 
                               (N880)? mem_q[1426] : 
                               (N875)? mem_q[1789] : 
                               (N877)? mem_q[2152] : 
                               (N879)? mem_q[2515] : 
                               (N881)? mem_q[2878] : 1'b0;
  assign commit_instr_o[698] = (N874)? mem_q[336] : 
                               (N876)? mem_q[699] : 
                               (N878)? mem_q[1062] : 
                               (N880)? mem_q[1425] : 
                               (N875)? mem_q[1788] : 
                               (N877)? mem_q[2151] : 
                               (N879)? mem_q[2514] : 
                               (N881)? mem_q[2877] : 1'b0;
  assign commit_instr_o[697] = (N874)? mem_q[335] : 
                               (N876)? mem_q[698] : 
                               (N878)? mem_q[1061] : 
                               (N880)? mem_q[1424] : 
                               (N875)? mem_q[1787] : 
                               (N877)? mem_q[2150] : 
                               (N879)? mem_q[2513] : 
                               (N881)? mem_q[2876] : 1'b0;
  assign commit_instr_o[696] = (N874)? mem_q[334] : 
                               (N876)? mem_q[697] : 
                               (N878)? mem_q[1060] : 
                               (N880)? mem_q[1423] : 
                               (N875)? mem_q[1786] : 
                               (N877)? mem_q[2149] : 
                               (N879)? mem_q[2512] : 
                               (N881)? mem_q[2875] : 1'b0;
  assign commit_instr_o[695] = (N874)? mem_q[333] : 
                               (N876)? mem_q[696] : 
                               (N878)? mem_q[1059] : 
                               (N880)? mem_q[1422] : 
                               (N875)? mem_q[1785] : 
                               (N877)? mem_q[2148] : 
                               (N879)? mem_q[2511] : 
                               (N881)? mem_q[2874] : 1'b0;
  assign commit_instr_o[694] = (N874)? mem_q[332] : 
                               (N876)? mem_q[695] : 
                               (N878)? mem_q[1058] : 
                               (N880)? mem_q[1421] : 
                               (N875)? mem_q[1784] : 
                               (N877)? mem_q[2147] : 
                               (N879)? mem_q[2510] : 
                               (N881)? mem_q[2873] : 1'b0;
  assign commit_instr_o[693] = (N874)? mem_q[331] : 
                               (N876)? mem_q[694] : 
                               (N878)? mem_q[1057] : 
                               (N880)? mem_q[1420] : 
                               (N875)? mem_q[1783] : 
                               (N877)? mem_q[2146] : 
                               (N879)? mem_q[2509] : 
                               (N881)? mem_q[2872] : 1'b0;
  assign commit_instr_o[692] = (N874)? mem_q[330] : 
                               (N876)? mem_q[693] : 
                               (N878)? mem_q[1056] : 
                               (N880)? mem_q[1419] : 
                               (N875)? mem_q[1782] : 
                               (N877)? mem_q[2145] : 
                               (N879)? mem_q[2508] : 
                               (N881)? mem_q[2871] : 1'b0;
  assign commit_instr_o[691] = (N874)? mem_q[329] : 
                               (N876)? mem_q[692] : 
                               (N878)? mem_q[1055] : 
                               (N880)? mem_q[1418] : 
                               (N875)? mem_q[1781] : 
                               (N877)? mem_q[2144] : 
                               (N879)? mem_q[2507] : 
                               (N881)? mem_q[2870] : 1'b0;
  assign commit_instr_o[690] = (N874)? mem_q[328] : 
                               (N876)? mem_q[691] : 
                               (N878)? mem_q[1054] : 
                               (N880)? mem_q[1417] : 
                               (N875)? mem_q[1780] : 
                               (N877)? mem_q[2143] : 
                               (N879)? mem_q[2506] : 
                               (N881)? mem_q[2869] : 1'b0;
  assign commit_instr_o[689] = (N874)? mem_q[327] : 
                               (N876)? mem_q[690] : 
                               (N878)? mem_q[1053] : 
                               (N880)? mem_q[1416] : 
                               (N875)? mem_q[1779] : 
                               (N877)? mem_q[2142] : 
                               (N879)? mem_q[2505] : 
                               (N881)? mem_q[2868] : 1'b0;
  assign commit_instr_o[688] = (N874)? mem_q[326] : 
                               (N876)? mem_q[689] : 
                               (N878)? mem_q[1052] : 
                               (N880)? mem_q[1415] : 
                               (N875)? mem_q[1778] : 
                               (N877)? mem_q[2141] : 
                               (N879)? mem_q[2504] : 
                               (N881)? mem_q[2867] : 1'b0;
  assign commit_instr_o[687] = (N874)? mem_q[325] : 
                               (N876)? mem_q[688] : 
                               (N878)? mem_q[1051] : 
                               (N880)? mem_q[1414] : 
                               (N875)? mem_q[1777] : 
                               (N877)? mem_q[2140] : 
                               (N879)? mem_q[2503] : 
                               (N881)? mem_q[2866] : 1'b0;
  assign commit_instr_o[686] = (N874)? mem_q[324] : 
                               (N876)? mem_q[687] : 
                               (N878)? mem_q[1050] : 
                               (N880)? mem_q[1413] : 
                               (N875)? mem_q[1776] : 
                               (N877)? mem_q[2139] : 
                               (N879)? mem_q[2502] : 
                               (N881)? mem_q[2865] : 1'b0;
  assign commit_instr_o[685] = (N874)? mem_q[323] : 
                               (N876)? mem_q[686] : 
                               (N878)? mem_q[1049] : 
                               (N880)? mem_q[1412] : 
                               (N875)? mem_q[1775] : 
                               (N877)? mem_q[2138] : 
                               (N879)? mem_q[2501] : 
                               (N881)? mem_q[2864] : 1'b0;
  assign commit_instr_o[684] = (N874)? mem_q[322] : 
                               (N876)? mem_q[685] : 
                               (N878)? mem_q[1048] : 
                               (N880)? mem_q[1411] : 
                               (N875)? mem_q[1774] : 
                               (N877)? mem_q[2137] : 
                               (N879)? mem_q[2500] : 
                               (N881)? mem_q[2863] : 1'b0;
  assign commit_instr_o[683] = (N874)? mem_q[321] : 
                               (N876)? mem_q[684] : 
                               (N878)? mem_q[1047] : 
                               (N880)? mem_q[1410] : 
                               (N875)? mem_q[1773] : 
                               (N877)? mem_q[2136] : 
                               (N879)? mem_q[2499] : 
                               (N881)? mem_q[2862] : 1'b0;
  assign commit_instr_o[682] = (N874)? mem_q[320] : 
                               (N876)? mem_q[683] : 
                               (N878)? mem_q[1046] : 
                               (N880)? mem_q[1409] : 
                               (N875)? mem_q[1772] : 
                               (N877)? mem_q[2135] : 
                               (N879)? mem_q[2498] : 
                               (N881)? mem_q[2861] : 1'b0;
  assign commit_instr_o[681] = (N874)? mem_q[319] : 
                               (N876)? mem_q[682] : 
                               (N878)? mem_q[1045] : 
                               (N880)? mem_q[1408] : 
                               (N875)? mem_q[1771] : 
                               (N877)? mem_q[2134] : 
                               (N879)? mem_q[2497] : 
                               (N881)? mem_q[2860] : 1'b0;
  assign commit_instr_o[680] = (N874)? mem_q[318] : 
                               (N876)? mem_q[681] : 
                               (N878)? mem_q[1044] : 
                               (N880)? mem_q[1407] : 
                               (N875)? mem_q[1770] : 
                               (N877)? mem_q[2133] : 
                               (N879)? mem_q[2496] : 
                               (N881)? mem_q[2859] : 1'b0;
  assign commit_instr_o[679] = (N874)? mem_q[317] : 
                               (N876)? mem_q[680] : 
                               (N878)? mem_q[1043] : 
                               (N880)? mem_q[1406] : 
                               (N875)? mem_q[1769] : 
                               (N877)? mem_q[2132] : 
                               (N879)? mem_q[2495] : 
                               (N881)? mem_q[2858] : 1'b0;
  assign commit_instr_o[678] = (N874)? mem_q[316] : 
                               (N876)? mem_q[679] : 
                               (N878)? mem_q[1042] : 
                               (N880)? mem_q[1405] : 
                               (N875)? mem_q[1768] : 
                               (N877)? mem_q[2131] : 
                               (N879)? mem_q[2494] : 
                               (N881)? mem_q[2857] : 1'b0;
  assign commit_instr_o[677] = (N874)? mem_q[315] : 
                               (N876)? mem_q[678] : 
                               (N878)? mem_q[1041] : 
                               (N880)? mem_q[1404] : 
                               (N875)? mem_q[1767] : 
                               (N877)? mem_q[2130] : 
                               (N879)? mem_q[2493] : 
                               (N881)? mem_q[2856] : 1'b0;
  assign commit_instr_o[676] = (N874)? mem_q[314] : 
                               (N876)? mem_q[677] : 
                               (N878)? mem_q[1040] : 
                               (N880)? mem_q[1403] : 
                               (N875)? mem_q[1766] : 
                               (N877)? mem_q[2129] : 
                               (N879)? mem_q[2492] : 
                               (N881)? mem_q[2855] : 1'b0;
  assign commit_instr_o[675] = (N874)? mem_q[313] : 
                               (N876)? mem_q[676] : 
                               (N878)? mem_q[1039] : 
                               (N880)? mem_q[1402] : 
                               (N875)? mem_q[1765] : 
                               (N877)? mem_q[2128] : 
                               (N879)? mem_q[2491] : 
                               (N881)? mem_q[2854] : 1'b0;
  assign commit_instr_o[674] = (N874)? mem_q[312] : 
                               (N876)? mem_q[675] : 
                               (N878)? mem_q[1038] : 
                               (N880)? mem_q[1401] : 
                               (N875)? mem_q[1764] : 
                               (N877)? mem_q[2127] : 
                               (N879)? mem_q[2490] : 
                               (N881)? mem_q[2853] : 1'b0;
  assign commit_instr_o[673] = (N874)? mem_q[311] : 
                               (N876)? mem_q[674] : 
                               (N878)? mem_q[1037] : 
                               (N880)? mem_q[1400] : 
                               (N875)? mem_q[1763] : 
                               (N877)? mem_q[2126] : 
                               (N879)? mem_q[2489] : 
                               (N881)? mem_q[2852] : 1'b0;
  assign commit_instr_o[672] = (N874)? mem_q[310] : 
                               (N876)? mem_q[673] : 
                               (N878)? mem_q[1036] : 
                               (N880)? mem_q[1399] : 
                               (N875)? mem_q[1762] : 
                               (N877)? mem_q[2125] : 
                               (N879)? mem_q[2488] : 
                               (N881)? mem_q[2851] : 1'b0;
  assign commit_instr_o[671] = (N874)? mem_q[309] : 
                               (N876)? mem_q[672] : 
                               (N878)? mem_q[1035] : 
                               (N880)? mem_q[1398] : 
                               (N875)? mem_q[1761] : 
                               (N877)? mem_q[2124] : 
                               (N879)? mem_q[2487] : 
                               (N881)? mem_q[2850] : 1'b0;
  assign commit_instr_o[670] = (N874)? mem_q[308] : 
                               (N876)? mem_q[671] : 
                               (N878)? mem_q[1034] : 
                               (N880)? mem_q[1397] : 
                               (N875)? mem_q[1760] : 
                               (N877)? mem_q[2123] : 
                               (N879)? mem_q[2486] : 
                               (N881)? mem_q[2849] : 1'b0;
  assign commit_instr_o[669] = (N874)? mem_q[307] : 
                               (N876)? mem_q[670] : 
                               (N878)? mem_q[1033] : 
                               (N880)? mem_q[1396] : 
                               (N875)? mem_q[1759] : 
                               (N877)? mem_q[2122] : 
                               (N879)? mem_q[2485] : 
                               (N881)? mem_q[2848] : 1'b0;
  assign commit_instr_o[668] = (N874)? mem_q[306] : 
                               (N876)? mem_q[669] : 
                               (N878)? mem_q[1032] : 
                               (N880)? mem_q[1395] : 
                               (N875)? mem_q[1758] : 
                               (N877)? mem_q[2121] : 
                               (N879)? mem_q[2484] : 
                               (N881)? mem_q[2847] : 1'b0;
  assign commit_instr_o[667] = (N874)? mem_q[305] : 
                               (N876)? mem_q[668] : 
                               (N878)? mem_q[1031] : 
                               (N880)? mem_q[1394] : 
                               (N875)? mem_q[1757] : 
                               (N877)? mem_q[2120] : 
                               (N879)? mem_q[2483] : 
                               (N881)? mem_q[2846] : 1'b0;
  assign commit_instr_o[666] = (N874)? mem_q[304] : 
                               (N876)? mem_q[667] : 
                               (N878)? mem_q[1030] : 
                               (N880)? mem_q[1393] : 
                               (N875)? mem_q[1756] : 
                               (N877)? mem_q[2119] : 
                               (N879)? mem_q[2482] : 
                               (N881)? mem_q[2845] : 1'b0;
  assign commit_instr_o[665] = (N874)? mem_q[303] : 
                               (N876)? mem_q[666] : 
                               (N878)? mem_q[1029] : 
                               (N880)? mem_q[1392] : 
                               (N875)? mem_q[1755] : 
                               (N877)? mem_q[2118] : 
                               (N879)? mem_q[2481] : 
                               (N881)? mem_q[2844] : 1'b0;
  assign commit_instr_o[664] = (N874)? mem_q[302] : 
                               (N876)? mem_q[665] : 
                               (N878)? mem_q[1028] : 
                               (N880)? mem_q[1391] : 
                               (N875)? mem_q[1754] : 
                               (N877)? mem_q[2117] : 
                               (N879)? mem_q[2480] : 
                               (N881)? mem_q[2843] : 1'b0;
  assign commit_instr_o[663] = (N874)? mem_q[301] : 
                               (N876)? mem_q[664] : 
                               (N878)? mem_q[1027] : 
                               (N880)? mem_q[1390] : 
                               (N875)? mem_q[1753] : 
                               (N877)? mem_q[2116] : 
                               (N879)? mem_q[2479] : 
                               (N881)? mem_q[2842] : 1'b0;
  assign commit_instr_o[662] = (N874)? mem_q[300] : 
                               (N876)? mem_q[663] : 
                               (N878)? mem_q[1026] : 
                               (N880)? mem_q[1389] : 
                               (N875)? mem_q[1752] : 
                               (N877)? mem_q[2115] : 
                               (N879)? mem_q[2478] : 
                               (N881)? mem_q[2841] : 1'b0;
  assign commit_instr_o[661] = (N874)? mem_q[299] : 
                               (N876)? mem_q[662] : 
                               (N878)? mem_q[1025] : 
                               (N880)? mem_q[1388] : 
                               (N875)? mem_q[1751] : 
                               (N877)? mem_q[2114] : 
                               (N879)? mem_q[2477] : 
                               (N881)? mem_q[2840] : 1'b0;
  assign commit_instr_o[660] = (N874)? mem_q[298] : 
                               (N876)? mem_q[661] : 
                               (N878)? mem_q[1024] : 
                               (N880)? mem_q[1387] : 
                               (N875)? mem_q[1750] : 
                               (N877)? mem_q[2113] : 
                               (N879)? mem_q[2476] : 
                               (N881)? mem_q[2839] : 1'b0;
  assign commit_instr_o[659] = (N874)? mem_q[297] : 
                               (N876)? mem_q[660] : 
                               (N878)? mem_q[1023] : 
                               (N880)? mem_q[1386] : 
                               (N875)? mem_q[1749] : 
                               (N877)? mem_q[2112] : 
                               (N879)? mem_q[2475] : 
                               (N881)? mem_q[2838] : 1'b0;
  assign commit_instr_o[658] = (N874)? mem_q[296] : 
                               (N876)? mem_q[659] : 
                               (N878)? mem_q[1022] : 
                               (N880)? mem_q[1385] : 
                               (N875)? mem_q[1748] : 
                               (N877)? mem_q[2111] : 
                               (N879)? mem_q[2474] : 
                               (N881)? mem_q[2837] : 1'b0;
  assign commit_instr_o[657] = (N874)? mem_q[295] : 
                               (N876)? mem_q[658] : 
                               (N878)? mem_q[1021] : 
                               (N880)? mem_q[1384] : 
                               (N875)? mem_q[1747] : 
                               (N877)? mem_q[2110] : 
                               (N879)? mem_q[2473] : 
                               (N881)? mem_q[2836] : 1'b0;
  assign commit_instr_o[656] = (N874)? mem_q[294] : 
                               (N876)? mem_q[657] : 
                               (N878)? mem_q[1020] : 
                               (N880)? mem_q[1383] : 
                               (N875)? mem_q[1746] : 
                               (N877)? mem_q[2109] : 
                               (N879)? mem_q[2472] : 
                               (N881)? mem_q[2835] : 1'b0;
  assign commit_instr_o[655] = (N874)? mem_q[293] : 
                               (N876)? mem_q[656] : 
                               (N878)? mem_q[1019] : 
                               (N880)? mem_q[1382] : 
                               (N875)? mem_q[1745] : 
                               (N877)? mem_q[2108] : 
                               (N879)? mem_q[2471] : 
                               (N881)? mem_q[2834] : 1'b0;
  assign commit_instr_o[654] = (N874)? mem_q[292] : 
                               (N876)? mem_q[655] : 
                               (N878)? mem_q[1018] : 
                               (N880)? mem_q[1381] : 
                               (N875)? mem_q[1744] : 
                               (N877)? mem_q[2107] : 
                               (N879)? mem_q[2470] : 
                               (N881)? mem_q[2833] : 1'b0;
  assign commit_instr_o[653] = (N874)? mem_q[291] : 
                               (N876)? mem_q[654] : 
                               (N878)? mem_q[1017] : 
                               (N880)? mem_q[1380] : 
                               (N875)? mem_q[1743] : 
                               (N877)? mem_q[2106] : 
                               (N879)? mem_q[2469] : 
                               (N881)? mem_q[2832] : 1'b0;
  assign commit_instr_o[652] = (N874)? mem_q[290] : 
                               (N876)? mem_q[653] : 
                               (N878)? mem_q[1016] : 
                               (N880)? mem_q[1379] : 
                               (N875)? mem_q[1742] : 
                               (N877)? mem_q[2105] : 
                               (N879)? mem_q[2468] : 
                               (N881)? mem_q[2831] : 1'b0;
  assign commit_instr_o[651] = (N874)? mem_q[289] : 
                               (N876)? mem_q[652] : 
                               (N878)? mem_q[1015] : 
                               (N880)? mem_q[1378] : 
                               (N875)? mem_q[1741] : 
                               (N877)? mem_q[2104] : 
                               (N879)? mem_q[2467] : 
                               (N881)? mem_q[2830] : 1'b0;
  assign commit_instr_o[650] = (N874)? mem_q[288] : 
                               (N876)? mem_q[651] : 
                               (N878)? mem_q[1014] : 
                               (N880)? mem_q[1377] : 
                               (N875)? mem_q[1740] : 
                               (N877)? mem_q[2103] : 
                               (N879)? mem_q[2466] : 
                               (N881)? mem_q[2829] : 1'b0;
  assign commit_instr_o[649] = (N874)? mem_q[287] : 
                               (N876)? mem_q[650] : 
                               (N878)? mem_q[1013] : 
                               (N880)? mem_q[1376] : 
                               (N875)? mem_q[1739] : 
                               (N877)? mem_q[2102] : 
                               (N879)? mem_q[2465] : 
                               (N881)? mem_q[2828] : 1'b0;
  assign commit_instr_o[648] = (N874)? mem_q[286] : 
                               (N876)? mem_q[649] : 
                               (N878)? mem_q[1012] : 
                               (N880)? mem_q[1375] : 
                               (N875)? mem_q[1738] : 
                               (N877)? mem_q[2101] : 
                               (N879)? mem_q[2464] : 
                               (N881)? mem_q[2827] : 1'b0;
  assign commit_instr_o[647] = (N874)? mem_q[285] : 
                               (N876)? mem_q[648] : 
                               (N878)? mem_q[1011] : 
                               (N880)? mem_q[1374] : 
                               (N875)? mem_q[1737] : 
                               (N877)? mem_q[2100] : 
                               (N879)? mem_q[2463] : 
                               (N881)? mem_q[2826] : 1'b0;
  assign commit_instr_o[646] = (N874)? mem_q[284] : 
                               (N876)? mem_q[647] : 
                               (N878)? mem_q[1010] : 
                               (N880)? mem_q[1373] : 
                               (N875)? mem_q[1736] : 
                               (N877)? mem_q[2099] : 
                               (N879)? mem_q[2462] : 
                               (N881)? mem_q[2825] : 1'b0;
  assign commit_instr_o[645] = (N874)? mem_q[283] : 
                               (N876)? mem_q[646] : 
                               (N878)? mem_q[1009] : 
                               (N880)? mem_q[1372] : 
                               (N875)? mem_q[1735] : 
                               (N877)? mem_q[2098] : 
                               (N879)? mem_q[2461] : 
                               (N881)? mem_q[2824] : 1'b0;
  assign commit_instr_o[644] = (N874)? mem_q[282] : 
                               (N876)? mem_q[645] : 
                               (N878)? mem_q[1008] : 
                               (N880)? mem_q[1371] : 
                               (N875)? mem_q[1734] : 
                               (N877)? mem_q[2097] : 
                               (N879)? mem_q[2460] : 
                               (N881)? mem_q[2823] : 1'b0;
  assign commit_instr_o[643] = (N874)? mem_q[281] : 
                               (N876)? mem_q[644] : 
                               (N878)? mem_q[1007] : 
                               (N880)? mem_q[1370] : 
                               (N875)? mem_q[1733] : 
                               (N877)? mem_q[2096] : 
                               (N879)? mem_q[2459] : 
                               (N881)? mem_q[2822] : 1'b0;
  assign commit_instr_o[642] = (N874)? mem_q[280] : 
                               (N876)? mem_q[643] : 
                               (N878)? mem_q[1006] : 
                               (N880)? mem_q[1369] : 
                               (N875)? mem_q[1732] : 
                               (N877)? mem_q[2095] : 
                               (N879)? mem_q[2458] : 
                               (N881)? mem_q[2821] : 1'b0;
  assign commit_instr_o[641] = (N874)? mem_q[279] : 
                               (N876)? mem_q[642] : 
                               (N878)? mem_q[1005] : 
                               (N880)? mem_q[1368] : 
                               (N875)? mem_q[1731] : 
                               (N877)? mem_q[2094] : 
                               (N879)? mem_q[2457] : 
                               (N881)? mem_q[2820] : 1'b0;
  assign commit_instr_o[640] = (N874)? mem_q[278] : 
                               (N876)? mem_q[641] : 
                               (N878)? mem_q[1004] : 
                               (N880)? mem_q[1367] : 
                               (N875)? mem_q[1730] : 
                               (N877)? mem_q[2093] : 
                               (N879)? mem_q[2456] : 
                               (N881)? mem_q[2819] : 1'b0;
  assign commit_instr_o[639] = (N874)? mem_q[277] : 
                               (N876)? mem_q[640] : 
                               (N878)? mem_q[1003] : 
                               (N880)? mem_q[1366] : 
                               (N875)? mem_q[1729] : 
                               (N877)? mem_q[2092] : 
                               (N879)? mem_q[2455] : 
                               (N881)? mem_q[2818] : 1'b0;
  assign commit_instr_o[638] = (N874)? mem_q[276] : 
                               (N876)? mem_q[639] : 
                               (N878)? mem_q[1002] : 
                               (N880)? mem_q[1365] : 
                               (N875)? mem_q[1728] : 
                               (N877)? mem_q[2091] : 
                               (N879)? mem_q[2454] : 
                               (N881)? mem_q[2817] : 1'b0;
  assign commit_instr_o[637] = (N874)? mem_q[275] : 
                               (N876)? mem_q[638] : 
                               (N878)? mem_q[1001] : 
                               (N880)? mem_q[1364] : 
                               (N875)? mem_q[1727] : 
                               (N877)? mem_q[2090] : 
                               (N879)? mem_q[2453] : 
                               (N881)? mem_q[2816] : 1'b0;
  assign commit_instr_o[636] = (N874)? mem_q[274] : 
                               (N876)? mem_q[637] : 
                               (N878)? mem_q[1000] : 
                               (N880)? mem_q[1363] : 
                               (N875)? mem_q[1726] : 
                               (N877)? mem_q[2089] : 
                               (N879)? mem_q[2452] : 
                               (N881)? mem_q[2815] : 1'b0;
  assign commit_instr_o[635] = (N874)? mem_q[273] : 
                               (N876)? mem_q[636] : 
                               (N878)? mem_q[999] : 
                               (N880)? mem_q[1362] : 
                               (N875)? mem_q[1725] : 
                               (N877)? mem_q[2088] : 
                               (N879)? mem_q[2451] : 
                               (N881)? mem_q[2814] : 1'b0;
  assign commit_instr_o[634] = (N874)? mem_q[272] : 
                               (N876)? mem_q[635] : 
                               (N878)? mem_q[998] : 
                               (N880)? mem_q[1361] : 
                               (N875)? mem_q[1724] : 
                               (N877)? mem_q[2087] : 
                               (N879)? mem_q[2450] : 
                               (N881)? mem_q[2813] : 1'b0;
  assign commit_instr_o[633] = (N874)? mem_q[271] : 
                               (N876)? mem_q[634] : 
                               (N878)? mem_q[997] : 
                               (N880)? mem_q[1360] : 
                               (N875)? mem_q[1723] : 
                               (N877)? mem_q[2086] : 
                               (N879)? mem_q[2449] : 
                               (N881)? mem_q[2812] : 1'b0;
  assign commit_instr_o[632] = (N874)? mem_q[270] : 
                               (N876)? mem_q[633] : 
                               (N878)? mem_q[996] : 
                               (N880)? mem_q[1359] : 
                               (N875)? mem_q[1722] : 
                               (N877)? mem_q[2085] : 
                               (N879)? mem_q[2448] : 
                               (N881)? mem_q[2811] : 1'b0;
  assign commit_instr_o[631] = (N874)? mem_q[269] : 
                               (N876)? mem_q[632] : 
                               (N878)? mem_q[995] : 
                               (N880)? mem_q[1358] : 
                               (N875)? mem_q[1721] : 
                               (N877)? mem_q[2084] : 
                               (N879)? mem_q[2447] : 
                               (N881)? mem_q[2810] : 1'b0;
  assign commit_instr_o[630] = (N874)? mem_q[268] : 
                               (N876)? mem_q[631] : 
                               (N878)? mem_q[994] : 
                               (N880)? mem_q[1357] : 
                               (N875)? mem_q[1720] : 
                               (N877)? mem_q[2083] : 
                               (N879)? mem_q[2446] : 
                               (N881)? mem_q[2809] : 1'b0;
  assign commit_instr_o[629] = (N874)? mem_q[267] : 
                               (N876)? mem_q[630] : 
                               (N878)? mem_q[993] : 
                               (N880)? mem_q[1356] : 
                               (N875)? mem_q[1719] : 
                               (N877)? mem_q[2082] : 
                               (N879)? mem_q[2445] : 
                               (N881)? mem_q[2808] : 1'b0;
  assign commit_instr_o[628] = (N874)? mem_q[266] : 
                               (N876)? mem_q[629] : 
                               (N878)? mem_q[992] : 
                               (N880)? mem_q[1355] : 
                               (N875)? mem_q[1718] : 
                               (N877)? mem_q[2081] : 
                               (N879)? mem_q[2444] : 
                               (N881)? mem_q[2807] : 1'b0;
  assign commit_instr_o[627] = (N874)? mem_q[265] : 
                               (N876)? mem_q[628] : 
                               (N878)? mem_q[991] : 
                               (N880)? mem_q[1354] : 
                               (N875)? mem_q[1717] : 
                               (N877)? mem_q[2080] : 
                               (N879)? mem_q[2443] : 
                               (N881)? mem_q[2806] : 1'b0;
  assign commit_instr_o[626] = (N874)? mem_q[264] : 
                               (N876)? mem_q[627] : 
                               (N878)? mem_q[990] : 
                               (N880)? mem_q[1353] : 
                               (N875)? mem_q[1716] : 
                               (N877)? mem_q[2079] : 
                               (N879)? mem_q[2442] : 
                               (N881)? mem_q[2805] : 1'b0;
  assign commit_instr_o[625] = (N874)? mem_q[263] : 
                               (N876)? mem_q[626] : 
                               (N878)? mem_q[989] : 
                               (N880)? mem_q[1352] : 
                               (N875)? mem_q[1715] : 
                               (N877)? mem_q[2078] : 
                               (N879)? mem_q[2441] : 
                               (N881)? mem_q[2804] : 1'b0;
  assign commit_instr_o[624] = (N874)? mem_q[262] : 
                               (N876)? mem_q[625] : 
                               (N878)? mem_q[988] : 
                               (N880)? mem_q[1351] : 
                               (N875)? mem_q[1714] : 
                               (N877)? mem_q[2077] : 
                               (N879)? mem_q[2440] : 
                               (N881)? mem_q[2803] : 1'b0;
  assign commit_instr_o[623] = (N874)? mem_q[261] : 
                               (N876)? mem_q[624] : 
                               (N878)? mem_q[987] : 
                               (N880)? mem_q[1350] : 
                               (N875)? mem_q[1713] : 
                               (N877)? mem_q[2076] : 
                               (N879)? mem_q[2439] : 
                               (N881)? mem_q[2802] : 1'b0;
  assign commit_instr_o[622] = (N874)? mem_q[260] : 
                               (N876)? mem_q[623] : 
                               (N878)? mem_q[986] : 
                               (N880)? mem_q[1349] : 
                               (N875)? mem_q[1712] : 
                               (N877)? mem_q[2075] : 
                               (N879)? mem_q[2438] : 
                               (N881)? mem_q[2801] : 1'b0;
  assign commit_instr_o[621] = (N874)? mem_q[259] : 
                               (N876)? mem_q[622] : 
                               (N878)? mem_q[985] : 
                               (N880)? mem_q[1348] : 
                               (N875)? mem_q[1711] : 
                               (N877)? mem_q[2074] : 
                               (N879)? mem_q[2437] : 
                               (N881)? mem_q[2800] : 1'b0;
  assign commit_instr_o[620] = (N874)? mem_q[258] : 
                               (N876)? mem_q[621] : 
                               (N878)? mem_q[984] : 
                               (N880)? mem_q[1347] : 
                               (N875)? mem_q[1710] : 
                               (N877)? mem_q[2073] : 
                               (N879)? mem_q[2436] : 
                               (N881)? mem_q[2799] : 1'b0;
  assign commit_instr_o[619] = (N874)? mem_q[257] : 
                               (N876)? mem_q[620] : 
                               (N878)? mem_q[983] : 
                               (N880)? mem_q[1346] : 
                               (N875)? mem_q[1709] : 
                               (N877)? mem_q[2072] : 
                               (N879)? mem_q[2435] : 
                               (N881)? mem_q[2798] : 1'b0;
  assign commit_instr_o[618] = (N874)? mem_q[256] : 
                               (N876)? mem_q[619] : 
                               (N878)? mem_q[982] : 
                               (N880)? mem_q[1345] : 
                               (N875)? mem_q[1708] : 
                               (N877)? mem_q[2071] : 
                               (N879)? mem_q[2434] : 
                               (N881)? mem_q[2797] : 1'b0;
  assign commit_instr_o[617] = (N874)? mem_q[255] : 
                               (N876)? mem_q[618] : 
                               (N878)? mem_q[981] : 
                               (N880)? mem_q[1344] : 
                               (N875)? mem_q[1707] : 
                               (N877)? mem_q[2070] : 
                               (N879)? mem_q[2433] : 
                               (N881)? mem_q[2796] : 1'b0;
  assign commit_instr_o[616] = (N874)? mem_q[254] : 
                               (N876)? mem_q[617] : 
                               (N878)? mem_q[980] : 
                               (N880)? mem_q[1343] : 
                               (N875)? mem_q[1706] : 
                               (N877)? mem_q[2069] : 
                               (N879)? mem_q[2432] : 
                               (N881)? mem_q[2795] : 1'b0;
  assign commit_instr_o[615] = (N874)? mem_q[253] : 
                               (N876)? mem_q[616] : 
                               (N878)? mem_q[979] : 
                               (N880)? mem_q[1342] : 
                               (N875)? mem_q[1705] : 
                               (N877)? mem_q[2068] : 
                               (N879)? mem_q[2431] : 
                               (N881)? mem_q[2794] : 1'b0;
  assign commit_instr_o[614] = (N874)? mem_q[252] : 
                               (N876)? mem_q[615] : 
                               (N878)? mem_q[978] : 
                               (N880)? mem_q[1341] : 
                               (N875)? mem_q[1704] : 
                               (N877)? mem_q[2067] : 
                               (N879)? mem_q[2430] : 
                               (N881)? mem_q[2793] : 1'b0;
  assign commit_instr_o[613] = (N874)? mem_q[251] : 
                               (N876)? mem_q[614] : 
                               (N878)? mem_q[977] : 
                               (N880)? mem_q[1340] : 
                               (N875)? mem_q[1703] : 
                               (N877)? mem_q[2066] : 
                               (N879)? mem_q[2429] : 
                               (N881)? mem_q[2792] : 1'b0;
  assign commit_instr_o[612] = (N874)? mem_q[250] : 
                               (N876)? mem_q[613] : 
                               (N878)? mem_q[976] : 
                               (N880)? mem_q[1339] : 
                               (N875)? mem_q[1702] : 
                               (N877)? mem_q[2065] : 
                               (N879)? mem_q[2428] : 
                               (N881)? mem_q[2791] : 1'b0;
  assign commit_instr_o[611] = (N874)? mem_q[249] : 
                               (N876)? mem_q[612] : 
                               (N878)? mem_q[975] : 
                               (N880)? mem_q[1338] : 
                               (N875)? mem_q[1701] : 
                               (N877)? mem_q[2064] : 
                               (N879)? mem_q[2427] : 
                               (N881)? mem_q[2790] : 1'b0;
  assign commit_instr_o[610] = (N874)? mem_q[248] : 
                               (N876)? mem_q[611] : 
                               (N878)? mem_q[974] : 
                               (N880)? mem_q[1337] : 
                               (N875)? mem_q[1700] : 
                               (N877)? mem_q[2063] : 
                               (N879)? mem_q[2426] : 
                               (N881)? mem_q[2789] : 1'b0;
  assign commit_instr_o[609] = (N874)? mem_q[247] : 
                               (N876)? mem_q[610] : 
                               (N878)? mem_q[973] : 
                               (N880)? mem_q[1336] : 
                               (N875)? mem_q[1699] : 
                               (N877)? mem_q[2062] : 
                               (N879)? mem_q[2425] : 
                               (N881)? mem_q[2788] : 1'b0;
  assign commit_instr_o[608] = (N874)? mem_q[246] : 
                               (N876)? mem_q[609] : 
                               (N878)? mem_q[972] : 
                               (N880)? mem_q[1335] : 
                               (N875)? mem_q[1698] : 
                               (N877)? mem_q[2061] : 
                               (N879)? mem_q[2424] : 
                               (N881)? mem_q[2787] : 1'b0;
  assign commit_instr_o[607] = (N874)? mem_q[245] : 
                               (N876)? mem_q[608] : 
                               (N878)? mem_q[971] : 
                               (N880)? mem_q[1334] : 
                               (N875)? mem_q[1697] : 
                               (N877)? mem_q[2060] : 
                               (N879)? mem_q[2423] : 
                               (N881)? mem_q[2786] : 1'b0;
  assign commit_instr_o[606] = (N874)? mem_q[244] : 
                               (N876)? mem_q[607] : 
                               (N878)? mem_q[970] : 
                               (N880)? mem_q[1333] : 
                               (N875)? mem_q[1696] : 
                               (N877)? mem_q[2059] : 
                               (N879)? mem_q[2422] : 
                               (N881)? mem_q[2785] : 1'b0;
  assign commit_instr_o[605] = (N874)? mem_q[243] : 
                               (N876)? mem_q[606] : 
                               (N878)? mem_q[969] : 
                               (N880)? mem_q[1332] : 
                               (N875)? mem_q[1695] : 
                               (N877)? mem_q[2058] : 
                               (N879)? mem_q[2421] : 
                               (N881)? mem_q[2784] : 1'b0;
  assign commit_instr_o[604] = (N874)? mem_q[242] : 
                               (N876)? mem_q[605] : 
                               (N878)? mem_q[968] : 
                               (N880)? mem_q[1331] : 
                               (N875)? mem_q[1694] : 
                               (N877)? mem_q[2057] : 
                               (N879)? mem_q[2420] : 
                               (N881)? mem_q[2783] : 1'b0;
  assign commit_instr_o[603] = (N874)? mem_q[241] : 
                               (N876)? mem_q[604] : 
                               (N878)? mem_q[967] : 
                               (N880)? mem_q[1330] : 
                               (N875)? mem_q[1693] : 
                               (N877)? mem_q[2056] : 
                               (N879)? mem_q[2419] : 
                               (N881)? mem_q[2782] : 1'b0;
  assign commit_instr_o[602] = (N874)? mem_q[240] : 
                               (N876)? mem_q[603] : 
                               (N878)? mem_q[966] : 
                               (N880)? mem_q[1329] : 
                               (N875)? mem_q[1692] : 
                               (N877)? mem_q[2055] : 
                               (N879)? mem_q[2418] : 
                               (N881)? mem_q[2781] : 1'b0;
  assign commit_instr_o[601] = (N874)? mem_q[239] : 
                               (N876)? mem_q[602] : 
                               (N878)? mem_q[965] : 
                               (N880)? mem_q[1328] : 
                               (N875)? mem_q[1691] : 
                               (N877)? mem_q[2054] : 
                               (N879)? mem_q[2417] : 
                               (N881)? mem_q[2780] : 1'b0;
  assign commit_instr_o[600] = (N874)? mem_q[238] : 
                               (N876)? mem_q[601] : 
                               (N878)? mem_q[964] : 
                               (N880)? mem_q[1327] : 
                               (N875)? mem_q[1690] : 
                               (N877)? mem_q[2053] : 
                               (N879)? mem_q[2416] : 
                               (N881)? mem_q[2779] : 1'b0;
  assign commit_instr_o[599] = (N874)? mem_q[237] : 
                               (N876)? mem_q[600] : 
                               (N878)? mem_q[963] : 
                               (N880)? mem_q[1326] : 
                               (N875)? mem_q[1689] : 
                               (N877)? mem_q[2052] : 
                               (N879)? mem_q[2415] : 
                               (N881)? mem_q[2778] : 1'b0;
  assign commit_instr_o[598] = (N874)? mem_q[236] : 
                               (N876)? mem_q[599] : 
                               (N878)? mem_q[962] : 
                               (N880)? mem_q[1325] : 
                               (N875)? mem_q[1688] : 
                               (N877)? mem_q[2051] : 
                               (N879)? mem_q[2414] : 
                               (N881)? mem_q[2777] : 1'b0;
  assign commit_instr_o[597] = (N874)? mem_q[235] : 
                               (N876)? mem_q[598] : 
                               (N878)? mem_q[961] : 
                               (N880)? mem_q[1324] : 
                               (N875)? mem_q[1687] : 
                               (N877)? mem_q[2050] : 
                               (N879)? mem_q[2413] : 
                               (N881)? mem_q[2776] : 1'b0;
  assign commit_instr_o[596] = (N874)? mem_q[234] : 
                               (N876)? mem_q[597] : 
                               (N878)? mem_q[960] : 
                               (N880)? mem_q[1323] : 
                               (N875)? mem_q[1686] : 
                               (N877)? mem_q[2049] : 
                               (N879)? mem_q[2412] : 
                               (N881)? mem_q[2775] : 1'b0;
  assign commit_instr_o[595] = (N874)? mem_q[233] : 
                               (N876)? mem_q[596] : 
                               (N878)? mem_q[959] : 
                               (N880)? mem_q[1322] : 
                               (N875)? mem_q[1685] : 
                               (N877)? mem_q[2048] : 
                               (N879)? mem_q[2411] : 
                               (N881)? mem_q[2774] : 1'b0;
  assign commit_instr_o[594] = (N874)? mem_q[232] : 
                               (N876)? mem_q[595] : 
                               (N878)? mem_q[958] : 
                               (N880)? mem_q[1321] : 
                               (N875)? mem_q[1684] : 
                               (N877)? mem_q[2047] : 
                               (N879)? mem_q[2410] : 
                               (N881)? mem_q[2773] : 1'b0;
  assign commit_instr_o[593] = (N874)? mem_q[231] : 
                               (N876)? mem_q[594] : 
                               (N878)? mem_q[957] : 
                               (N880)? mem_q[1320] : 
                               (N875)? mem_q[1683] : 
                               (N877)? mem_q[2046] : 
                               (N879)? mem_q[2409] : 
                               (N881)? mem_q[2772] : 1'b0;
  assign commit_instr_o[592] = (N874)? mem_q[230] : 
                               (N876)? mem_q[593] : 
                               (N878)? mem_q[956] : 
                               (N880)? mem_q[1319] : 
                               (N875)? mem_q[1682] : 
                               (N877)? mem_q[2045] : 
                               (N879)? mem_q[2408] : 
                               (N881)? mem_q[2771] : 1'b0;
  assign commit_instr_o[591] = (N874)? mem_q[229] : 
                               (N876)? mem_q[592] : 
                               (N878)? mem_q[955] : 
                               (N880)? mem_q[1318] : 
                               (N875)? mem_q[1681] : 
                               (N877)? mem_q[2044] : 
                               (N879)? mem_q[2407] : 
                               (N881)? mem_q[2770] : 1'b0;
  assign commit_instr_o[590] = (N874)? mem_q[228] : 
                               (N876)? mem_q[591] : 
                               (N878)? mem_q[954] : 
                               (N880)? mem_q[1317] : 
                               (N875)? mem_q[1680] : 
                               (N877)? mem_q[2043] : 
                               (N879)? mem_q[2406] : 
                               (N881)? mem_q[2769] : 1'b0;
  assign commit_instr_o[589] = (N874)? mem_q[227] : 
                               (N876)? mem_q[590] : 
                               (N878)? mem_q[953] : 
                               (N880)? mem_q[1316] : 
                               (N875)? mem_q[1679] : 
                               (N877)? mem_q[2042] : 
                               (N879)? mem_q[2405] : 
                               (N881)? mem_q[2768] : 1'b0;
  assign commit_instr_o[588] = (N874)? mem_q[226] : 
                               (N876)? mem_q[589] : 
                               (N878)? mem_q[952] : 
                               (N880)? mem_q[1315] : 
                               (N875)? mem_q[1678] : 
                               (N877)? mem_q[2041] : 
                               (N879)? mem_q[2404] : 
                               (N881)? mem_q[2767] : 1'b0;
  assign commit_instr_o[587] = (N874)? mem_q[225] : 
                               (N876)? mem_q[588] : 
                               (N878)? mem_q[951] : 
                               (N880)? mem_q[1314] : 
                               (N875)? mem_q[1677] : 
                               (N877)? mem_q[2040] : 
                               (N879)? mem_q[2403] : 
                               (N881)? mem_q[2766] : 1'b0;
  assign commit_instr_o[586] = (N874)? mem_q[224] : 
                               (N876)? mem_q[587] : 
                               (N878)? mem_q[950] : 
                               (N880)? mem_q[1313] : 
                               (N875)? mem_q[1676] : 
                               (N877)? mem_q[2039] : 
                               (N879)? mem_q[2402] : 
                               (N881)? mem_q[2765] : 1'b0;
  assign commit_instr_o[585] = (N874)? mem_q[223] : 
                               (N876)? mem_q[586] : 
                               (N878)? mem_q[949] : 
                               (N880)? mem_q[1312] : 
                               (N875)? mem_q[1675] : 
                               (N877)? mem_q[2038] : 
                               (N879)? mem_q[2401] : 
                               (N881)? mem_q[2764] : 1'b0;
  assign commit_instr_o[584] = (N874)? mem_q[222] : 
                               (N876)? mem_q[585] : 
                               (N878)? mem_q[948] : 
                               (N880)? mem_q[1311] : 
                               (N875)? mem_q[1674] : 
                               (N877)? mem_q[2037] : 
                               (N879)? mem_q[2400] : 
                               (N881)? mem_q[2763] : 1'b0;
  assign commit_instr_o[583] = (N874)? mem_q[221] : 
                               (N876)? mem_q[584] : 
                               (N878)? mem_q[947] : 
                               (N880)? mem_q[1310] : 
                               (N875)? mem_q[1673] : 
                               (N877)? mem_q[2036] : 
                               (N879)? mem_q[2399] : 
                               (N881)? mem_q[2762] : 1'b0;
  assign commit_instr_o[582] = (N874)? mem_q[220] : 
                               (N876)? mem_q[583] : 
                               (N878)? mem_q[946] : 
                               (N880)? mem_q[1309] : 
                               (N875)? mem_q[1672] : 
                               (N877)? mem_q[2035] : 
                               (N879)? mem_q[2398] : 
                               (N881)? mem_q[2761] : 1'b0;
  assign commit_instr_o[581] = (N874)? mem_q[219] : 
                               (N876)? mem_q[582] : 
                               (N878)? mem_q[945] : 
                               (N880)? mem_q[1308] : 
                               (N875)? mem_q[1671] : 
                               (N877)? mem_q[2034] : 
                               (N879)? mem_q[2397] : 
                               (N881)? mem_q[2760] : 1'b0;
  assign commit_instr_o[580] = (N874)? mem_q[218] : 
                               (N876)? mem_q[581] : 
                               (N878)? mem_q[944] : 
                               (N880)? mem_q[1307] : 
                               (N875)? mem_q[1670] : 
                               (N877)? mem_q[2033] : 
                               (N879)? mem_q[2396] : 
                               (N881)? mem_q[2759] : 1'b0;
  assign commit_instr_o[579] = (N874)? mem_q[217] : 
                               (N876)? mem_q[580] : 
                               (N878)? mem_q[943] : 
                               (N880)? mem_q[1306] : 
                               (N875)? mem_q[1669] : 
                               (N877)? mem_q[2032] : 
                               (N879)? mem_q[2395] : 
                               (N881)? mem_q[2758] : 1'b0;
  assign commit_instr_o[578] = (N874)? mem_q[216] : 
                               (N876)? mem_q[579] : 
                               (N878)? mem_q[942] : 
                               (N880)? mem_q[1305] : 
                               (N875)? mem_q[1668] : 
                               (N877)? mem_q[2031] : 
                               (N879)? mem_q[2394] : 
                               (N881)? mem_q[2757] : 1'b0;
  assign commit_instr_o[577] = (N874)? mem_q[215] : 
                               (N876)? mem_q[578] : 
                               (N878)? mem_q[941] : 
                               (N880)? mem_q[1304] : 
                               (N875)? mem_q[1667] : 
                               (N877)? mem_q[2030] : 
                               (N879)? mem_q[2393] : 
                               (N881)? mem_q[2756] : 1'b0;
  assign commit_instr_o[576] = (N874)? mem_q[214] : 
                               (N876)? mem_q[577] : 
                               (N878)? mem_q[940] : 
                               (N880)? mem_q[1303] : 
                               (N875)? mem_q[1666] : 
                               (N877)? mem_q[2029] : 
                               (N879)? mem_q[2392] : 
                               (N881)? mem_q[2755] : 1'b0;
  assign commit_instr_o[575] = (N874)? mem_q[213] : 
                               (N876)? mem_q[576] : 
                               (N878)? mem_q[939] : 
                               (N880)? mem_q[1302] : 
                               (N875)? mem_q[1665] : 
                               (N877)? mem_q[2028] : 
                               (N879)? mem_q[2391] : 
                               (N881)? mem_q[2754] : 1'b0;
  assign commit_instr_o[574] = (N874)? mem_q[212] : 
                               (N876)? mem_q[575] : 
                               (N878)? mem_q[938] : 
                               (N880)? mem_q[1301] : 
                               (N875)? mem_q[1664] : 
                               (N877)? mem_q[2027] : 
                               (N879)? mem_q[2390] : 
                               (N881)? mem_q[2753] : 1'b0;
  assign commit_instr_o[573] = (N874)? mem_q[211] : 
                               (N876)? mem_q[574] : 
                               (N878)? mem_q[937] : 
                               (N880)? mem_q[1300] : 
                               (N875)? mem_q[1663] : 
                               (N877)? mem_q[2026] : 
                               (N879)? mem_q[2389] : 
                               (N881)? mem_q[2752] : 1'b0;
  assign commit_instr_o[572] = (N874)? mem_q[210] : 
                               (N876)? mem_q[573] : 
                               (N878)? mem_q[936] : 
                               (N880)? mem_q[1299] : 
                               (N875)? mem_q[1662] : 
                               (N877)? mem_q[2025] : 
                               (N879)? mem_q[2388] : 
                               (N881)? mem_q[2751] : 1'b0;
  assign commit_instr_o[571] = (N874)? mem_q[209] : 
                               (N876)? mem_q[572] : 
                               (N878)? mem_q[935] : 
                               (N880)? mem_q[1298] : 
                               (N875)? mem_q[1661] : 
                               (N877)? mem_q[2024] : 
                               (N879)? mem_q[2387] : 
                               (N881)? mem_q[2750] : 1'b0;
  assign commit_instr_o[570] = (N874)? mem_q[208] : 
                               (N876)? mem_q[571] : 
                               (N878)? mem_q[934] : 
                               (N880)? mem_q[1297] : 
                               (N875)? mem_q[1660] : 
                               (N877)? mem_q[2023] : 
                               (N879)? mem_q[2386] : 
                               (N881)? mem_q[2749] : 1'b0;
  assign commit_instr_o[569] = (N874)? mem_q[207] : 
                               (N876)? mem_q[570] : 
                               (N878)? mem_q[933] : 
                               (N880)? mem_q[1296] : 
                               (N875)? mem_q[1659] : 
                               (N877)? mem_q[2022] : 
                               (N879)? mem_q[2385] : 
                               (N881)? mem_q[2748] : 1'b0;
  assign commit_instr_o[568] = (N874)? mem_q[206] : 
                               (N876)? mem_q[569] : 
                               (N878)? mem_q[932] : 
                               (N880)? mem_q[1295] : 
                               (N875)? mem_q[1658] : 
                               (N877)? mem_q[2021] : 
                               (N879)? mem_q[2384] : 
                               (N881)? mem_q[2747] : 1'b0;
  assign commit_instr_o[567] = (N874)? mem_q[205] : 
                               (N876)? mem_q[568] : 
                               (N878)? mem_q[931] : 
                               (N880)? mem_q[1294] : 
                               (N875)? mem_q[1657] : 
                               (N877)? mem_q[2020] : 
                               (N879)? mem_q[2383] : 
                               (N881)? mem_q[2746] : 1'b0;
  assign commit_instr_o[566] = (N874)? mem_q[204] : 
                               (N876)? mem_q[567] : 
                               (N878)? mem_q[930] : 
                               (N880)? mem_q[1293] : 
                               (N875)? mem_q[1656] : 
                               (N877)? mem_q[2019] : 
                               (N879)? mem_q[2382] : 
                               (N881)? mem_q[2745] : 1'b0;
  assign commit_instr_o[565] = (N874)? mem_q[203] : 
                               (N876)? mem_q[566] : 
                               (N878)? mem_q[929] : 
                               (N880)? mem_q[1292] : 
                               (N875)? mem_q[1655] : 
                               (N877)? mem_q[2018] : 
                               (N879)? mem_q[2381] : 
                               (N881)? mem_q[2744] : 1'b0;
  assign commit_instr_o[564] = (N874)? mem_q[202] : 
                               (N876)? mem_q[565] : 
                               (N878)? mem_q[928] : 
                               (N880)? mem_q[1291] : 
                               (N875)? mem_q[1654] : 
                               (N877)? mem_q[2017] : 
                               (N879)? mem_q[2380] : 
                               (N881)? mem_q[2743] : 1'b0;
  assign commit_instr_o[563] = (N874)? mem_q[201] : 
                               (N876)? mem_q[564] : 
                               (N878)? mem_q[927] : 
                               (N880)? mem_q[1290] : 
                               (N875)? mem_q[1653] : 
                               (N877)? mem_q[2016] : 
                               (N879)? mem_q[2379] : 
                               (N881)? mem_q[2742] : 1'b0;
  assign commit_instr_o[562] = (N874)? mem_q[200] : 
                               (N876)? mem_q[563] : 
                               (N878)? mem_q[926] : 
                               (N880)? mem_q[1289] : 
                               (N875)? mem_q[1652] : 
                               (N877)? mem_q[2015] : 
                               (N879)? mem_q[2378] : 
                               (N881)? mem_q[2741] : 1'b0;
  assign commit_instr_o[561] = (N874)? mem_q[199] : 
                               (N876)? mem_q[562] : 
                               (N878)? mem_q[925] : 
                               (N880)? mem_q[1288] : 
                               (N875)? mem_q[1651] : 
                               (N877)? mem_q[2014] : 
                               (N879)? mem_q[2377] : 
                               (N881)? mem_q[2740] : 1'b0;
  assign commit_instr_o[560] = (N874)? mem_q[198] : 
                               (N876)? mem_q[561] : 
                               (N878)? mem_q[924] : 
                               (N880)? mem_q[1287] : 
                               (N875)? mem_q[1650] : 
                               (N877)? mem_q[2013] : 
                               (N879)? mem_q[2376] : 
                               (N881)? mem_q[2739] : 1'b0;
  assign commit_instr_o[559] = (N874)? mem_q[197] : 
                               (N876)? mem_q[560] : 
                               (N878)? mem_q[923] : 
                               (N880)? mem_q[1286] : 
                               (N875)? mem_q[1649] : 
                               (N877)? mem_q[2012] : 
                               (N879)? mem_q[2375] : 
                               (N881)? mem_q[2738] : 1'b0;
  assign commit_instr_o[558] = (N874)? mem_q[196] : 
                               (N876)? mem_q[559] : 
                               (N878)? mem_q[922] : 
                               (N880)? mem_q[1285] : 
                               (N875)? mem_q[1648] : 
                               (N877)? mem_q[2011] : 
                               (N879)? mem_q[2374] : 
                               (N881)? mem_q[2737] : 1'b0;
  assign commit_instr_o[557] = (N874)? mem_q[195] : 
                               (N876)? mem_q[558] : 
                               (N878)? mem_q[921] : 
                               (N880)? mem_q[1284] : 
                               (N875)? mem_q[1647] : 
                               (N877)? mem_q[2010] : 
                               (N879)? mem_q[2373] : 
                               (N881)? mem_q[2736] : 1'b0;
  assign commit_instr_o[556] = (N874)? mem_q[194] : 
                               (N876)? mem_q[557] : 
                               (N878)? mem_q[920] : 
                               (N880)? mem_q[1283] : 
                               (N875)? mem_q[1646] : 
                               (N877)? mem_q[2009] : 
                               (N879)? mem_q[2372] : 
                               (N881)? mem_q[2735] : 1'b0;
  assign commit_instr_o[555] = (N874)? mem_q[193] : 
                               (N876)? mem_q[556] : 
                               (N878)? mem_q[919] : 
                               (N880)? mem_q[1282] : 
                               (N875)? mem_q[1645] : 
                               (N877)? mem_q[2008] : 
                               (N879)? mem_q[2371] : 
                               (N881)? mem_q[2734] : 1'b0;
  assign commit_instr_o[554] = (N874)? mem_q[192] : 
                               (N876)? mem_q[555] : 
                               (N878)? mem_q[918] : 
                               (N880)? mem_q[1281] : 
                               (N875)? mem_q[1644] : 
                               (N877)? mem_q[2007] : 
                               (N879)? mem_q[2370] : 
                               (N881)? mem_q[2733] : 1'b0;
  assign commit_instr_o[553] = (N874)? mem_q[191] : 
                               (N876)? mem_q[554] : 
                               (N878)? mem_q[917] : 
                               (N880)? mem_q[1280] : 
                               (N875)? mem_q[1643] : 
                               (N877)? mem_q[2006] : 
                               (N879)? mem_q[2369] : 
                               (N881)? mem_q[2732] : 1'b0;
  assign commit_instr_o[552] = (N874)? mem_q[190] : 
                               (N876)? mem_q[553] : 
                               (N878)? mem_q[916] : 
                               (N880)? mem_q[1279] : 
                               (N875)? mem_q[1642] : 
                               (N877)? mem_q[2005] : 
                               (N879)? mem_q[2368] : 
                               (N881)? mem_q[2731] : 1'b0;
  assign commit_instr_o[551] = (N874)? mem_q[189] : 
                               (N876)? mem_q[552] : 
                               (N878)? mem_q[915] : 
                               (N880)? mem_q[1278] : 
                               (N875)? mem_q[1641] : 
                               (N877)? mem_q[2004] : 
                               (N879)? mem_q[2367] : 
                               (N881)? mem_q[2730] : 1'b0;
  assign commit_instr_o[550] = (N874)? mem_q[188] : 
                               (N876)? mem_q[551] : 
                               (N878)? mem_q[914] : 
                               (N880)? mem_q[1277] : 
                               (N875)? mem_q[1640] : 
                               (N877)? mem_q[2003] : 
                               (N879)? mem_q[2366] : 
                               (N881)? mem_q[2729] : 1'b0;
  assign commit_instr_o[549] = (N874)? mem_q[187] : 
                               (N876)? mem_q[550] : 
                               (N878)? mem_q[913] : 
                               (N880)? mem_q[1276] : 
                               (N875)? mem_q[1639] : 
                               (N877)? mem_q[2002] : 
                               (N879)? mem_q[2365] : 
                               (N881)? mem_q[2728] : 1'b0;
  assign commit_instr_o[548] = (N874)? mem_q[186] : 
                               (N876)? mem_q[549] : 
                               (N878)? mem_q[912] : 
                               (N880)? mem_q[1275] : 
                               (N875)? mem_q[1638] : 
                               (N877)? mem_q[2001] : 
                               (N879)? mem_q[2364] : 
                               (N881)? mem_q[2727] : 1'b0;
  assign commit_instr_o[547] = (N874)? mem_q[185] : 
                               (N876)? mem_q[548] : 
                               (N878)? mem_q[911] : 
                               (N880)? mem_q[1274] : 
                               (N875)? mem_q[1637] : 
                               (N877)? mem_q[2000] : 
                               (N879)? mem_q[2363] : 
                               (N881)? mem_q[2726] : 1'b0;
  assign commit_instr_o[546] = (N874)? mem_q[184] : 
                               (N876)? mem_q[547] : 
                               (N878)? mem_q[910] : 
                               (N880)? mem_q[1273] : 
                               (N875)? mem_q[1636] : 
                               (N877)? mem_q[1999] : 
                               (N879)? mem_q[2362] : 
                               (N881)? mem_q[2725] : 1'b0;
  assign commit_instr_o[545] = (N874)? mem_q[183] : 
                               (N876)? mem_q[546] : 
                               (N878)? mem_q[909] : 
                               (N880)? mem_q[1272] : 
                               (N875)? mem_q[1635] : 
                               (N877)? mem_q[1998] : 
                               (N879)? mem_q[2361] : 
                               (N881)? mem_q[2724] : 1'b0;
  assign commit_instr_o[544] = (N874)? mem_q[182] : 
                               (N876)? mem_q[545] : 
                               (N878)? mem_q[908] : 
                               (N880)? mem_q[1271] : 
                               (N875)? mem_q[1634] : 
                               (N877)? mem_q[1997] : 
                               (N879)? mem_q[2360] : 
                               (N881)? mem_q[2723] : 1'b0;
  assign commit_instr_o[543] = (N874)? mem_q[181] : 
                               (N876)? mem_q[544] : 
                               (N878)? mem_q[907] : 
                               (N880)? mem_q[1270] : 
                               (N875)? mem_q[1633] : 
                               (N877)? mem_q[1996] : 
                               (N879)? mem_q[2359] : 
                               (N881)? mem_q[2722] : 1'b0;
  assign commit_instr_o[542] = (N874)? mem_q[180] : 
                               (N876)? mem_q[543] : 
                               (N878)? mem_q[906] : 
                               (N880)? mem_q[1269] : 
                               (N875)? mem_q[1632] : 
                               (N877)? mem_q[1995] : 
                               (N879)? mem_q[2358] : 
                               (N881)? mem_q[2721] : 1'b0;
  assign commit_instr_o[541] = (N874)? mem_q[179] : 
                               (N876)? mem_q[542] : 
                               (N878)? mem_q[905] : 
                               (N880)? mem_q[1268] : 
                               (N875)? mem_q[1631] : 
                               (N877)? mem_q[1994] : 
                               (N879)? mem_q[2357] : 
                               (N881)? mem_q[2720] : 1'b0;
  assign commit_instr_o[540] = (N874)? mem_q[178] : 
                               (N876)? mem_q[541] : 
                               (N878)? mem_q[904] : 
                               (N880)? mem_q[1267] : 
                               (N875)? mem_q[1630] : 
                               (N877)? mem_q[1993] : 
                               (N879)? mem_q[2356] : 
                               (N881)? mem_q[2719] : 1'b0;
  assign commit_instr_o[539] = (N874)? mem_q[177] : 
                               (N876)? mem_q[540] : 
                               (N878)? mem_q[903] : 
                               (N880)? mem_q[1266] : 
                               (N875)? mem_q[1629] : 
                               (N877)? mem_q[1992] : 
                               (N879)? mem_q[2355] : 
                               (N881)? mem_q[2718] : 1'b0;
  assign commit_instr_o[538] = (N874)? mem_q[176] : 
                               (N876)? mem_q[539] : 
                               (N878)? mem_q[902] : 
                               (N880)? mem_q[1265] : 
                               (N875)? mem_q[1628] : 
                               (N877)? mem_q[1991] : 
                               (N879)? mem_q[2354] : 
                               (N881)? mem_q[2717] : 1'b0;
  assign commit_instr_o[537] = (N874)? mem_q[175] : 
                               (N876)? mem_q[538] : 
                               (N878)? mem_q[901] : 
                               (N880)? mem_q[1264] : 
                               (N875)? mem_q[1627] : 
                               (N877)? mem_q[1990] : 
                               (N879)? mem_q[2353] : 
                               (N881)? mem_q[2716] : 1'b0;
  assign commit_instr_o[536] = (N874)? mem_q[174] : 
                               (N876)? mem_q[537] : 
                               (N878)? mem_q[900] : 
                               (N880)? mem_q[1263] : 
                               (N875)? mem_q[1626] : 
                               (N877)? mem_q[1989] : 
                               (N879)? mem_q[2352] : 
                               (N881)? mem_q[2715] : 1'b0;
  assign commit_instr_o[535] = (N874)? mem_q[173] : 
                               (N876)? mem_q[536] : 
                               (N878)? mem_q[899] : 
                               (N880)? mem_q[1262] : 
                               (N875)? mem_q[1625] : 
                               (N877)? mem_q[1988] : 
                               (N879)? mem_q[2351] : 
                               (N881)? mem_q[2714] : 1'b0;
  assign commit_instr_o[534] = (N874)? mem_q[172] : 
                               (N876)? mem_q[535] : 
                               (N878)? mem_q[898] : 
                               (N880)? mem_q[1261] : 
                               (N875)? mem_q[1624] : 
                               (N877)? mem_q[1987] : 
                               (N879)? mem_q[2350] : 
                               (N881)? mem_q[2713] : 1'b0;
  assign commit_instr_o[533] = (N874)? mem_q[171] : 
                               (N876)? mem_q[534] : 
                               (N878)? mem_q[897] : 
                               (N880)? mem_q[1260] : 
                               (N875)? mem_q[1623] : 
                               (N877)? mem_q[1986] : 
                               (N879)? mem_q[2349] : 
                               (N881)? mem_q[2712] : 1'b0;
  assign commit_instr_o[532] = (N874)? mem_q[170] : 
                               (N876)? mem_q[533] : 
                               (N878)? mem_q[896] : 
                               (N880)? mem_q[1259] : 
                               (N875)? mem_q[1622] : 
                               (N877)? mem_q[1985] : 
                               (N879)? mem_q[2348] : 
                               (N881)? mem_q[2711] : 1'b0;
  assign commit_instr_o[531] = (N874)? mem_q[169] : 
                               (N876)? mem_q[532] : 
                               (N878)? mem_q[895] : 
                               (N880)? mem_q[1258] : 
                               (N875)? mem_q[1621] : 
                               (N877)? mem_q[1984] : 
                               (N879)? mem_q[2347] : 
                               (N881)? mem_q[2710] : 1'b0;
  assign commit_instr_o[530] = (N874)? mem_q[168] : 
                               (N876)? mem_q[531] : 
                               (N878)? mem_q[894] : 
                               (N880)? mem_q[1257] : 
                               (N875)? mem_q[1620] : 
                               (N877)? mem_q[1983] : 
                               (N879)? mem_q[2346] : 
                               (N881)? mem_q[2709] : 1'b0;
  assign commit_instr_o[529] = (N874)? mem_q[167] : 
                               (N876)? mem_q[530] : 
                               (N878)? mem_q[893] : 
                               (N880)? mem_q[1256] : 
                               (N875)? mem_q[1619] : 
                               (N877)? mem_q[1982] : 
                               (N879)? mem_q[2345] : 
                               (N881)? mem_q[2708] : 1'b0;
  assign commit_instr_o[528] = (N874)? mem_q[166] : 
                               (N876)? mem_q[529] : 
                               (N878)? mem_q[892] : 
                               (N880)? mem_q[1255] : 
                               (N875)? mem_q[1618] : 
                               (N877)? mem_q[1981] : 
                               (N879)? mem_q[2344] : 
                               (N881)? mem_q[2707] : 1'b0;
  assign commit_instr_o[527] = (N874)? mem_q[165] : 
                               (N876)? mem_q[528] : 
                               (N878)? mem_q[891] : 
                               (N880)? mem_q[1254] : 
                               (N875)? mem_q[1617] : 
                               (N877)? mem_q[1980] : 
                               (N879)? mem_q[2343] : 
                               (N881)? mem_q[2706] : 1'b0;
  assign commit_instr_o[526] = (N874)? mem_q[164] : 
                               (N876)? mem_q[527] : 
                               (N878)? mem_q[890] : 
                               (N880)? mem_q[1253] : 
                               (N875)? mem_q[1616] : 
                               (N877)? mem_q[1979] : 
                               (N879)? mem_q[2342] : 
                               (N881)? mem_q[2705] : 1'b0;
  assign commit_instr_o[525] = (N874)? mem_q[163] : 
                               (N876)? mem_q[526] : 
                               (N878)? mem_q[889] : 
                               (N880)? mem_q[1252] : 
                               (N875)? mem_q[1615] : 
                               (N877)? mem_q[1978] : 
                               (N879)? mem_q[2341] : 
                               (N881)? mem_q[2704] : 1'b0;
  assign commit_instr_o[524] = (N874)? mem_q[162] : 
                               (N876)? mem_q[525] : 
                               (N878)? mem_q[888] : 
                               (N880)? mem_q[1251] : 
                               (N875)? mem_q[1614] : 
                               (N877)? mem_q[1977] : 
                               (N879)? mem_q[2340] : 
                               (N881)? mem_q[2703] : 1'b0;
  assign commit_instr_o[523] = (N874)? mem_q[161] : 
                               (N876)? mem_q[524] : 
                               (N878)? mem_q[887] : 
                               (N880)? mem_q[1250] : 
                               (N875)? mem_q[1613] : 
                               (N877)? mem_q[1976] : 
                               (N879)? mem_q[2339] : 
                               (N881)? mem_q[2702] : 1'b0;
  assign commit_instr_o[522] = (N874)? mem_q[160] : 
                               (N876)? mem_q[523] : 
                               (N878)? mem_q[886] : 
                               (N880)? mem_q[1249] : 
                               (N875)? mem_q[1612] : 
                               (N877)? mem_q[1975] : 
                               (N879)? mem_q[2338] : 
                               (N881)? mem_q[2701] : 1'b0;
  assign commit_instr_o[521] = (N874)? mem_q[159] : 
                               (N876)? mem_q[522] : 
                               (N878)? mem_q[885] : 
                               (N880)? mem_q[1248] : 
                               (N875)? mem_q[1611] : 
                               (N877)? mem_q[1974] : 
                               (N879)? mem_q[2337] : 
                               (N881)? mem_q[2700] : 1'b0;
  assign commit_instr_o[520] = (N874)? mem_q[158] : 
                               (N876)? mem_q[521] : 
                               (N878)? mem_q[884] : 
                               (N880)? mem_q[1247] : 
                               (N875)? mem_q[1610] : 
                               (N877)? mem_q[1973] : 
                               (N879)? mem_q[2336] : 
                               (N881)? mem_q[2699] : 1'b0;
  assign commit_instr_o[519] = (N874)? mem_q[157] : 
                               (N876)? mem_q[520] : 
                               (N878)? mem_q[883] : 
                               (N880)? mem_q[1246] : 
                               (N875)? mem_q[1609] : 
                               (N877)? mem_q[1972] : 
                               (N879)? mem_q[2335] : 
                               (N881)? mem_q[2698] : 1'b0;
  assign commit_instr_o[518] = (N874)? mem_q[156] : 
                               (N876)? mem_q[519] : 
                               (N878)? mem_q[882] : 
                               (N880)? mem_q[1245] : 
                               (N875)? mem_q[1608] : 
                               (N877)? mem_q[1971] : 
                               (N879)? mem_q[2334] : 
                               (N881)? mem_q[2697] : 1'b0;
  assign commit_instr_o[517] = (N874)? mem_q[155] : 
                               (N876)? mem_q[518] : 
                               (N878)? mem_q[881] : 
                               (N880)? mem_q[1244] : 
                               (N875)? mem_q[1607] : 
                               (N877)? mem_q[1970] : 
                               (N879)? mem_q[2333] : 
                               (N881)? mem_q[2696] : 1'b0;
  assign commit_instr_o[516] = (N874)? mem_q[154] : 
                               (N876)? mem_q[517] : 
                               (N878)? mem_q[880] : 
                               (N880)? mem_q[1243] : 
                               (N875)? mem_q[1606] : 
                               (N877)? mem_q[1969] : 
                               (N879)? mem_q[2332] : 
                               (N881)? mem_q[2695] : 1'b0;
  assign commit_instr_o[515] = (N874)? mem_q[153] : 
                               (N876)? mem_q[516] : 
                               (N878)? mem_q[879] : 
                               (N880)? mem_q[1242] : 
                               (N875)? mem_q[1605] : 
                               (N877)? mem_q[1968] : 
                               (N879)? mem_q[2331] : 
                               (N881)? mem_q[2694] : 1'b0;
  assign commit_instr_o[514] = (N874)? mem_q[152] : 
                               (N876)? mem_q[515] : 
                               (N878)? mem_q[878] : 
                               (N880)? mem_q[1241] : 
                               (N875)? mem_q[1604] : 
                               (N877)? mem_q[1967] : 
                               (N879)? mem_q[2330] : 
                               (N881)? mem_q[2693] : 1'b0;
  assign commit_instr_o[513] = (N874)? mem_q[151] : 
                               (N876)? mem_q[514] : 
                               (N878)? mem_q[877] : 
                               (N880)? mem_q[1240] : 
                               (N875)? mem_q[1603] : 
                               (N877)? mem_q[1966] : 
                               (N879)? mem_q[2329] : 
                               (N881)? mem_q[2692] : 1'b0;
  assign commit_instr_o[512] = (N874)? mem_q[150] : 
                               (N876)? mem_q[513] : 
                               (N878)? mem_q[876] : 
                               (N880)? mem_q[1239] : 
                               (N875)? mem_q[1602] : 
                               (N877)? mem_q[1965] : 
                               (N879)? mem_q[2328] : 
                               (N881)? mem_q[2691] : 1'b0;
  assign commit_instr_o[511] = (N874)? mem_q[149] : 
                               (N876)? mem_q[512] : 
                               (N878)? mem_q[875] : 
                               (N880)? mem_q[1238] : 
                               (N875)? mem_q[1601] : 
                               (N877)? mem_q[1964] : 
                               (N879)? mem_q[2327] : 
                               (N881)? mem_q[2690] : 1'b0;
  assign commit_instr_o[510] = (N874)? mem_q[148] : 
                               (N876)? mem_q[511] : 
                               (N878)? mem_q[874] : 
                               (N880)? mem_q[1237] : 
                               (N875)? mem_q[1600] : 
                               (N877)? mem_q[1963] : 
                               (N879)? mem_q[2326] : 
                               (N881)? mem_q[2689] : 1'b0;
  assign commit_instr_o[509] = (N874)? mem_q[147] : 
                               (N876)? mem_q[510] : 
                               (N878)? mem_q[873] : 
                               (N880)? mem_q[1236] : 
                               (N875)? mem_q[1599] : 
                               (N877)? mem_q[1962] : 
                               (N879)? mem_q[2325] : 
                               (N881)? mem_q[2688] : 1'b0;
  assign commit_instr_o[508] = (N874)? mem_q[146] : 
                               (N876)? mem_q[509] : 
                               (N878)? mem_q[872] : 
                               (N880)? mem_q[1235] : 
                               (N875)? mem_q[1598] : 
                               (N877)? mem_q[1961] : 
                               (N879)? mem_q[2324] : 
                               (N881)? mem_q[2687] : 1'b0;
  assign commit_instr_o[507] = (N874)? mem_q[145] : 
                               (N876)? mem_q[508] : 
                               (N878)? mem_q[871] : 
                               (N880)? mem_q[1234] : 
                               (N875)? mem_q[1597] : 
                               (N877)? mem_q[1960] : 
                               (N879)? mem_q[2323] : 
                               (N881)? mem_q[2686] : 1'b0;
  assign commit_instr_o[506] = (N874)? mem_q[144] : 
                               (N876)? mem_q[507] : 
                               (N878)? mem_q[870] : 
                               (N880)? mem_q[1233] : 
                               (N875)? mem_q[1596] : 
                               (N877)? mem_q[1959] : 
                               (N879)? mem_q[2322] : 
                               (N881)? mem_q[2685] : 1'b0;
  assign commit_instr_o[505] = (N874)? mem_q[143] : 
                               (N876)? mem_q[506] : 
                               (N878)? mem_q[869] : 
                               (N880)? mem_q[1232] : 
                               (N875)? mem_q[1595] : 
                               (N877)? mem_q[1958] : 
                               (N879)? mem_q[2321] : 
                               (N881)? mem_q[2684] : 1'b0;
  assign commit_instr_o[504] = (N874)? mem_q[142] : 
                               (N876)? mem_q[505] : 
                               (N878)? mem_q[868] : 
                               (N880)? mem_q[1231] : 
                               (N875)? mem_q[1594] : 
                               (N877)? mem_q[1957] : 
                               (N879)? mem_q[2320] : 
                               (N881)? mem_q[2683] : 1'b0;
  assign commit_instr_o[503] = (N874)? mem_q[141] : 
                               (N876)? mem_q[504] : 
                               (N878)? mem_q[867] : 
                               (N880)? mem_q[1230] : 
                               (N875)? mem_q[1593] : 
                               (N877)? mem_q[1956] : 
                               (N879)? mem_q[2319] : 
                               (N881)? mem_q[2682] : 1'b0;
  assign commit_instr_o[502] = (N874)? mem_q[140] : 
                               (N876)? mem_q[503] : 
                               (N878)? mem_q[866] : 
                               (N880)? mem_q[1229] : 
                               (N875)? mem_q[1592] : 
                               (N877)? mem_q[1955] : 
                               (N879)? mem_q[2318] : 
                               (N881)? mem_q[2681] : 1'b0;
  assign commit_instr_o[501] = (N874)? mem_q[139] : 
                               (N876)? mem_q[502] : 
                               (N878)? mem_q[865] : 
                               (N880)? mem_q[1228] : 
                               (N875)? mem_q[1591] : 
                               (N877)? mem_q[1954] : 
                               (N879)? mem_q[2317] : 
                               (N881)? mem_q[2680] : 1'b0;
  assign commit_instr_o[500] = (N874)? mem_q[138] : 
                               (N876)? mem_q[501] : 
                               (N878)? mem_q[864] : 
                               (N880)? mem_q[1227] : 
                               (N875)? mem_q[1590] : 
                               (N877)? mem_q[1953] : 
                               (N879)? mem_q[2316] : 
                               (N881)? mem_q[2679] : 1'b0;
  assign commit_instr_o[499] = (N874)? mem_q[137] : 
                               (N876)? mem_q[500] : 
                               (N878)? mem_q[863] : 
                               (N880)? mem_q[1226] : 
                               (N875)? mem_q[1589] : 
                               (N877)? mem_q[1952] : 
                               (N879)? mem_q[2315] : 
                               (N881)? mem_q[2678] : 1'b0;
  assign commit_instr_o[498] = (N874)? mem_q[136] : 
                               (N876)? mem_q[499] : 
                               (N878)? mem_q[862] : 
                               (N880)? mem_q[1225] : 
                               (N875)? mem_q[1588] : 
                               (N877)? mem_q[1951] : 
                               (N879)? mem_q[2314] : 
                               (N881)? mem_q[2677] : 1'b0;
  assign commit_instr_o[497] = (N874)? mem_q[135] : 
                               (N876)? mem_q[498] : 
                               (N878)? mem_q[861] : 
                               (N880)? mem_q[1224] : 
                               (N875)? mem_q[1587] : 
                               (N877)? mem_q[1950] : 
                               (N879)? mem_q[2313] : 
                               (N881)? mem_q[2676] : 1'b0;
  assign commit_instr_o[496] = (N874)? mem_q[134] : 
                               (N876)? mem_q[497] : 
                               (N878)? mem_q[860] : 
                               (N880)? mem_q[1223] : 
                               (N875)? mem_q[1586] : 
                               (N877)? mem_q[1949] : 
                               (N879)? mem_q[2312] : 
                               (N881)? mem_q[2675] : 1'b0;
  assign commit_instr_o[495] = (N874)? mem_q[133] : 
                               (N876)? mem_q[496] : 
                               (N878)? mem_q[859] : 
                               (N880)? mem_q[1222] : 
                               (N875)? mem_q[1585] : 
                               (N877)? mem_q[1948] : 
                               (N879)? mem_q[2311] : 
                               (N881)? mem_q[2674] : 1'b0;
  assign commit_instr_o[494] = (N874)? mem_q[132] : 
                               (N876)? mem_q[495] : 
                               (N878)? mem_q[858] : 
                               (N880)? mem_q[1221] : 
                               (N875)? mem_q[1584] : 
                               (N877)? mem_q[1947] : 
                               (N879)? mem_q[2310] : 
                               (N881)? mem_q[2673] : 1'b0;
  assign commit_instr_o[493] = (N874)? mem_q[131] : 
                               (N876)? mem_q[494] : 
                               (N878)? mem_q[857] : 
                               (N880)? mem_q[1220] : 
                               (N875)? mem_q[1583] : 
                               (N877)? mem_q[1946] : 
                               (N879)? mem_q[2309] : 
                               (N881)? mem_q[2672] : 1'b0;
  assign commit_instr_o[492] = (N874)? mem_q[130] : 
                               (N876)? mem_q[493] : 
                               (N878)? mem_q[856] : 
                               (N880)? mem_q[1219] : 
                               (N875)? mem_q[1582] : 
                               (N877)? mem_q[1945] : 
                               (N879)? mem_q[2308] : 
                               (N881)? mem_q[2671] : 1'b0;
  assign commit_instr_o[491] = (N874)? mem_q[129] : 
                               (N876)? mem_q[492] : 
                               (N878)? mem_q[855] : 
                               (N880)? mem_q[1218] : 
                               (N875)? mem_q[1581] : 
                               (N877)? mem_q[1944] : 
                               (N879)? mem_q[2307] : 
                               (N881)? mem_q[2670] : 1'b0;
  assign commit_instr_o[490] = (N874)? mem_q[128] : 
                               (N876)? mem_q[491] : 
                               (N878)? mem_q[854] : 
                               (N880)? mem_q[1217] : 
                               (N875)? mem_q[1580] : 
                               (N877)? mem_q[1943] : 
                               (N879)? mem_q[2306] : 
                               (N881)? mem_q[2669] : 1'b0;
  assign commit_instr_o[489] = (N874)? mem_q[127] : 
                               (N876)? mem_q[490] : 
                               (N878)? mem_q[853] : 
                               (N880)? mem_q[1216] : 
                               (N875)? mem_q[1579] : 
                               (N877)? mem_q[1942] : 
                               (N879)? mem_q[2305] : 
                               (N881)? mem_q[2668] : 1'b0;
  assign commit_instr_o[488] = (N874)? mem_q[126] : 
                               (N876)? mem_q[489] : 
                               (N878)? mem_q[852] : 
                               (N880)? mem_q[1215] : 
                               (N875)? mem_q[1578] : 
                               (N877)? mem_q[1941] : 
                               (N879)? mem_q[2304] : 
                               (N881)? mem_q[2667] : 1'b0;
  assign commit_instr_o[487] = (N874)? mem_q[125] : 
                               (N876)? mem_q[488] : 
                               (N878)? mem_q[851] : 
                               (N880)? mem_q[1214] : 
                               (N875)? mem_q[1577] : 
                               (N877)? mem_q[1940] : 
                               (N879)? mem_q[2303] : 
                               (N881)? mem_q[2666] : 1'b0;
  assign commit_instr_o[486] = (N874)? mem_q[124] : 
                               (N876)? mem_q[487] : 
                               (N878)? mem_q[850] : 
                               (N880)? mem_q[1213] : 
                               (N875)? mem_q[1576] : 
                               (N877)? mem_q[1939] : 
                               (N879)? mem_q[2302] : 
                               (N881)? mem_q[2665] : 1'b0;
  assign commit_instr_o[485] = (N874)? mem_q[123] : 
                               (N876)? mem_q[486] : 
                               (N878)? mem_q[849] : 
                               (N880)? mem_q[1212] : 
                               (N875)? mem_q[1575] : 
                               (N877)? mem_q[1938] : 
                               (N879)? mem_q[2301] : 
                               (N881)? mem_q[2664] : 1'b0;
  assign commit_instr_o[484] = (N874)? mem_q[122] : 
                               (N876)? mem_q[485] : 
                               (N878)? mem_q[848] : 
                               (N880)? mem_q[1211] : 
                               (N875)? mem_q[1574] : 
                               (N877)? mem_q[1937] : 
                               (N879)? mem_q[2300] : 
                               (N881)? mem_q[2663] : 1'b0;
  assign commit_instr_o[483] = (N874)? mem_q[121] : 
                               (N876)? mem_q[484] : 
                               (N878)? mem_q[847] : 
                               (N880)? mem_q[1210] : 
                               (N875)? mem_q[1573] : 
                               (N877)? mem_q[1936] : 
                               (N879)? mem_q[2299] : 
                               (N881)? mem_q[2662] : 1'b0;
  assign commit_instr_o[482] = (N874)? mem_q[120] : 
                               (N876)? mem_q[483] : 
                               (N878)? mem_q[846] : 
                               (N880)? mem_q[1209] : 
                               (N875)? mem_q[1572] : 
                               (N877)? mem_q[1935] : 
                               (N879)? mem_q[2298] : 
                               (N881)? mem_q[2661] : 1'b0;
  assign commit_instr_o[481] = (N874)? mem_q[119] : 
                               (N876)? mem_q[482] : 
                               (N878)? mem_q[845] : 
                               (N880)? mem_q[1208] : 
                               (N875)? mem_q[1571] : 
                               (N877)? mem_q[1934] : 
                               (N879)? mem_q[2297] : 
                               (N881)? mem_q[2660] : 1'b0;
  assign commit_instr_o[480] = (N874)? mem_q[118] : 
                               (N876)? mem_q[481] : 
                               (N878)? mem_q[844] : 
                               (N880)? mem_q[1207] : 
                               (N875)? mem_q[1570] : 
                               (N877)? mem_q[1933] : 
                               (N879)? mem_q[2296] : 
                               (N881)? mem_q[2659] : 1'b0;
  assign commit_instr_o[479] = (N874)? mem_q[117] : 
                               (N876)? mem_q[480] : 
                               (N878)? mem_q[843] : 
                               (N880)? mem_q[1206] : 
                               (N875)? mem_q[1569] : 
                               (N877)? mem_q[1932] : 
                               (N879)? mem_q[2295] : 
                               (N881)? mem_q[2658] : 1'b0;
  assign commit_instr_o[478] = (N874)? mem_q[116] : 
                               (N876)? mem_q[479] : 
                               (N878)? mem_q[842] : 
                               (N880)? mem_q[1205] : 
                               (N875)? mem_q[1568] : 
                               (N877)? mem_q[1931] : 
                               (N879)? mem_q[2294] : 
                               (N881)? mem_q[2657] : 1'b0;
  assign commit_instr_o[477] = (N874)? mem_q[115] : 
                               (N876)? mem_q[478] : 
                               (N878)? mem_q[841] : 
                               (N880)? mem_q[1204] : 
                               (N875)? mem_q[1567] : 
                               (N877)? mem_q[1930] : 
                               (N879)? mem_q[2293] : 
                               (N881)? mem_q[2656] : 1'b0;
  assign commit_instr_o[476] = (N874)? mem_q[114] : 
                               (N876)? mem_q[477] : 
                               (N878)? mem_q[840] : 
                               (N880)? mem_q[1203] : 
                               (N875)? mem_q[1566] : 
                               (N877)? mem_q[1929] : 
                               (N879)? mem_q[2292] : 
                               (N881)? mem_q[2655] : 1'b0;
  assign commit_instr_o[475] = (N874)? mem_q[113] : 
                               (N876)? mem_q[476] : 
                               (N878)? mem_q[839] : 
                               (N880)? mem_q[1202] : 
                               (N875)? mem_q[1565] : 
                               (N877)? mem_q[1928] : 
                               (N879)? mem_q[2291] : 
                               (N881)? mem_q[2654] : 1'b0;
  assign commit_instr_o[474] = (N874)? mem_q[112] : 
                               (N876)? mem_q[475] : 
                               (N878)? mem_q[838] : 
                               (N880)? mem_q[1201] : 
                               (N875)? mem_q[1564] : 
                               (N877)? mem_q[1927] : 
                               (N879)? mem_q[2290] : 
                               (N881)? mem_q[2653] : 1'b0;
  assign commit_instr_o[473] = (N874)? mem_q[111] : 
                               (N876)? mem_q[474] : 
                               (N878)? mem_q[837] : 
                               (N880)? mem_q[1200] : 
                               (N875)? mem_q[1563] : 
                               (N877)? mem_q[1926] : 
                               (N879)? mem_q[2289] : 
                               (N881)? mem_q[2652] : 1'b0;
  assign commit_instr_o[472] = (N874)? mem_q[110] : 
                               (N876)? mem_q[473] : 
                               (N878)? mem_q[836] : 
                               (N880)? mem_q[1199] : 
                               (N875)? mem_q[1562] : 
                               (N877)? mem_q[1925] : 
                               (N879)? mem_q[2288] : 
                               (N881)? mem_q[2651] : 1'b0;
  assign commit_instr_o[471] = (N874)? mem_q[109] : 
                               (N876)? mem_q[472] : 
                               (N878)? mem_q[835] : 
                               (N880)? mem_q[1198] : 
                               (N875)? mem_q[1561] : 
                               (N877)? mem_q[1924] : 
                               (N879)? mem_q[2287] : 
                               (N881)? mem_q[2650] : 1'b0;
  assign commit_instr_o[470] = (N874)? mem_q[108] : 
                               (N876)? mem_q[471] : 
                               (N878)? mem_q[834] : 
                               (N880)? mem_q[1197] : 
                               (N875)? mem_q[1560] : 
                               (N877)? mem_q[1923] : 
                               (N879)? mem_q[2286] : 
                               (N881)? mem_q[2649] : 1'b0;
  assign commit_instr_o[469] = (N874)? mem_q[107] : 
                               (N876)? mem_q[470] : 
                               (N878)? mem_q[833] : 
                               (N880)? mem_q[1196] : 
                               (N875)? mem_q[1559] : 
                               (N877)? mem_q[1922] : 
                               (N879)? mem_q[2285] : 
                               (N881)? mem_q[2648] : 1'b0;
  assign commit_instr_o[468] = (N874)? mem_q[106] : 
                               (N876)? mem_q[469] : 
                               (N878)? mem_q[832] : 
                               (N880)? mem_q[1195] : 
                               (N875)? mem_q[1558] : 
                               (N877)? mem_q[1921] : 
                               (N879)? mem_q[2284] : 
                               (N881)? mem_q[2647] : 1'b0;
  assign commit_instr_o[467] = (N874)? mem_q[105] : 
                               (N876)? mem_q[468] : 
                               (N878)? mem_q[831] : 
                               (N880)? mem_q[1194] : 
                               (N875)? mem_q[1557] : 
                               (N877)? mem_q[1920] : 
                               (N879)? mem_q[2283] : 
                               (N881)? mem_q[2646] : 1'b0;
  assign commit_instr_o[466] = (N874)? mem_q[104] : 
                               (N876)? mem_q[467] : 
                               (N878)? mem_q[830] : 
                               (N880)? mem_q[1193] : 
                               (N875)? mem_q[1556] : 
                               (N877)? mem_q[1919] : 
                               (N879)? mem_q[2282] : 
                               (N881)? mem_q[2645] : 1'b0;
  assign commit_instr_o[465] = (N874)? mem_q[103] : 
                               (N876)? mem_q[466] : 
                               (N878)? mem_q[829] : 
                               (N880)? mem_q[1192] : 
                               (N875)? mem_q[1555] : 
                               (N877)? mem_q[1918] : 
                               (N879)? mem_q[2281] : 
                               (N881)? mem_q[2644] : 1'b0;
  assign commit_instr_o[464] = (N874)? mem_q[102] : 
                               (N876)? mem_q[465] : 
                               (N878)? mem_q[828] : 
                               (N880)? mem_q[1191] : 
                               (N875)? mem_q[1554] : 
                               (N877)? mem_q[1917] : 
                               (N879)? mem_q[2280] : 
                               (N881)? mem_q[2643] : 1'b0;
  assign commit_instr_o[463] = (N874)? mem_q[101] : 
                               (N876)? mem_q[464] : 
                               (N878)? mem_q[827] : 
                               (N880)? mem_q[1190] : 
                               (N875)? mem_q[1553] : 
                               (N877)? mem_q[1916] : 
                               (N879)? mem_q[2279] : 
                               (N881)? mem_q[2642] : 1'b0;
  assign commit_instr_o[462] = (N874)? mem_q[100] : 
                               (N876)? mem_q[463] : 
                               (N878)? mem_q[826] : 
                               (N880)? mem_q[1189] : 
                               (N875)? mem_q[1552] : 
                               (N877)? mem_q[1915] : 
                               (N879)? mem_q[2278] : 
                               (N881)? mem_q[2641] : 1'b0;
  assign commit_instr_o[461] = (N874)? mem_q[99] : 
                               (N876)? mem_q[462] : 
                               (N878)? mem_q[825] : 
                               (N880)? mem_q[1188] : 
                               (N875)? mem_q[1551] : 
                               (N877)? mem_q[1914] : 
                               (N879)? mem_q[2277] : 
                               (N881)? mem_q[2640] : 1'b0;
  assign commit_instr_o[460] = (N874)? mem_q[98] : 
                               (N876)? mem_q[461] : 
                               (N878)? mem_q[824] : 
                               (N880)? mem_q[1187] : 
                               (N875)? mem_q[1550] : 
                               (N877)? mem_q[1913] : 
                               (N879)? mem_q[2276] : 
                               (N881)? mem_q[2639] : 1'b0;
  assign commit_instr_o[459] = (N874)? mem_q[97] : 
                               (N876)? mem_q[460] : 
                               (N878)? mem_q[823] : 
                               (N880)? mem_q[1186] : 
                               (N875)? mem_q[1549] : 
                               (N877)? mem_q[1912] : 
                               (N879)? mem_q[2275] : 
                               (N881)? mem_q[2638] : 1'b0;
  assign commit_instr_o[458] = (N874)? mem_q[96] : 
                               (N876)? mem_q[459] : 
                               (N878)? mem_q[822] : 
                               (N880)? mem_q[1185] : 
                               (N875)? mem_q[1548] : 
                               (N877)? mem_q[1911] : 
                               (N879)? mem_q[2274] : 
                               (N881)? mem_q[2637] : 1'b0;
  assign commit_instr_o[457] = (N874)? mem_q[95] : 
                               (N876)? mem_q[458] : 
                               (N878)? mem_q[821] : 
                               (N880)? mem_q[1184] : 
                               (N875)? mem_q[1547] : 
                               (N877)? mem_q[1910] : 
                               (N879)? mem_q[2273] : 
                               (N881)? mem_q[2636] : 1'b0;
  assign commit_instr_o[456] = (N874)? mem_q[94] : 
                               (N876)? mem_q[457] : 
                               (N878)? mem_q[820] : 
                               (N880)? mem_q[1183] : 
                               (N875)? mem_q[1546] : 
                               (N877)? mem_q[1909] : 
                               (N879)? mem_q[2272] : 
                               (N881)? mem_q[2635] : 1'b0;
  assign commit_instr_o[455] = (N874)? mem_q[93] : 
                               (N876)? mem_q[456] : 
                               (N878)? mem_q[819] : 
                               (N880)? mem_q[1182] : 
                               (N875)? mem_q[1545] : 
                               (N877)? mem_q[1908] : 
                               (N879)? mem_q[2271] : 
                               (N881)? mem_q[2634] : 1'b0;
  assign commit_instr_o[454] = (N874)? mem_q[92] : 
                               (N876)? mem_q[455] : 
                               (N878)? mem_q[818] : 
                               (N880)? mem_q[1181] : 
                               (N875)? mem_q[1544] : 
                               (N877)? mem_q[1907] : 
                               (N879)? mem_q[2270] : 
                               (N881)? mem_q[2633] : 1'b0;
  assign commit_instr_o[453] = (N874)? mem_q[91] : 
                               (N876)? mem_q[454] : 
                               (N878)? mem_q[817] : 
                               (N880)? mem_q[1180] : 
                               (N875)? mem_q[1543] : 
                               (N877)? mem_q[1906] : 
                               (N879)? mem_q[2269] : 
                               (N881)? mem_q[2632] : 1'b0;
  assign commit_instr_o[452] = (N874)? mem_q[90] : 
                               (N876)? mem_q[453] : 
                               (N878)? mem_q[816] : 
                               (N880)? mem_q[1179] : 
                               (N875)? mem_q[1542] : 
                               (N877)? mem_q[1905] : 
                               (N879)? mem_q[2268] : 
                               (N881)? mem_q[2631] : 1'b0;
  assign commit_instr_o[451] = (N874)? mem_q[89] : 
                               (N876)? mem_q[452] : 
                               (N878)? mem_q[815] : 
                               (N880)? mem_q[1178] : 
                               (N875)? mem_q[1541] : 
                               (N877)? mem_q[1904] : 
                               (N879)? mem_q[2267] : 
                               (N881)? mem_q[2630] : 1'b0;
  assign commit_instr_o[450] = (N874)? mem_q[88] : 
                               (N876)? mem_q[451] : 
                               (N878)? mem_q[814] : 
                               (N880)? mem_q[1177] : 
                               (N875)? mem_q[1540] : 
                               (N877)? mem_q[1903] : 
                               (N879)? mem_q[2266] : 
                               (N881)? mem_q[2629] : 1'b0;
  assign commit_instr_o[449] = (N874)? mem_q[87] : 
                               (N876)? mem_q[450] : 
                               (N878)? mem_q[813] : 
                               (N880)? mem_q[1176] : 
                               (N875)? mem_q[1539] : 
                               (N877)? mem_q[1902] : 
                               (N879)? mem_q[2265] : 
                               (N881)? mem_q[2628] : 1'b0;
  assign commit_instr_o[448] = (N874)? mem_q[86] : 
                               (N876)? mem_q[449] : 
                               (N878)? mem_q[812] : 
                               (N880)? mem_q[1175] : 
                               (N875)? mem_q[1538] : 
                               (N877)? mem_q[1901] : 
                               (N879)? mem_q[2264] : 
                               (N881)? mem_q[2627] : 1'b0;
  assign commit_instr_o[447] = (N874)? mem_q[85] : 
                               (N876)? mem_q[448] : 
                               (N878)? mem_q[811] : 
                               (N880)? mem_q[1174] : 
                               (N875)? mem_q[1537] : 
                               (N877)? mem_q[1900] : 
                               (N879)? mem_q[2263] : 
                               (N881)? mem_q[2626] : 1'b0;
  assign commit_instr_o[446] = (N874)? mem_q[84] : 
                               (N876)? mem_q[447] : 
                               (N878)? mem_q[810] : 
                               (N880)? mem_q[1173] : 
                               (N875)? mem_q[1536] : 
                               (N877)? mem_q[1899] : 
                               (N879)? mem_q[2262] : 
                               (N881)? mem_q[2625] : 1'b0;
  assign commit_instr_o[445] = (N874)? mem_q[83] : 
                               (N876)? mem_q[446] : 
                               (N878)? mem_q[809] : 
                               (N880)? mem_q[1172] : 
                               (N875)? mem_q[1535] : 
                               (N877)? mem_q[1898] : 
                               (N879)? mem_q[2261] : 
                               (N881)? mem_q[2624] : 1'b0;
  assign commit_instr_o[444] = (N874)? mem_q[82] : 
                               (N876)? mem_q[445] : 
                               (N878)? mem_q[808] : 
                               (N880)? mem_q[1171] : 
                               (N875)? mem_q[1534] : 
                               (N877)? mem_q[1897] : 
                               (N879)? mem_q[2260] : 
                               (N881)? mem_q[2623] : 1'b0;
  assign commit_instr_o[443] = (N874)? mem_q[81] : 
                               (N876)? mem_q[444] : 
                               (N878)? mem_q[807] : 
                               (N880)? mem_q[1170] : 
                               (N875)? mem_q[1533] : 
                               (N877)? mem_q[1896] : 
                               (N879)? mem_q[2259] : 
                               (N881)? mem_q[2622] : 1'b0;
  assign commit_instr_o[442] = (N874)? mem_q[80] : 
                               (N876)? mem_q[443] : 
                               (N878)? mem_q[806] : 
                               (N880)? mem_q[1169] : 
                               (N875)? mem_q[1532] : 
                               (N877)? mem_q[1895] : 
                               (N879)? mem_q[2258] : 
                               (N881)? mem_q[2621] : 1'b0;
  assign commit_instr_o[441] = (N874)? mem_q[79] : 
                               (N876)? mem_q[442] : 
                               (N878)? mem_q[805] : 
                               (N880)? mem_q[1168] : 
                               (N875)? mem_q[1531] : 
                               (N877)? mem_q[1894] : 
                               (N879)? mem_q[2257] : 
                               (N881)? mem_q[2620] : 1'b0;
  assign commit_instr_o[440] = (N874)? mem_q[78] : 
                               (N876)? mem_q[441] : 
                               (N878)? mem_q[804] : 
                               (N880)? mem_q[1167] : 
                               (N875)? mem_q[1530] : 
                               (N877)? mem_q[1893] : 
                               (N879)? mem_q[2256] : 
                               (N881)? mem_q[2619] : 1'b0;
  assign commit_instr_o[439] = (N874)? mem_q[77] : 
                               (N876)? mem_q[440] : 
                               (N878)? mem_q[803] : 
                               (N880)? mem_q[1166] : 
                               (N875)? mem_q[1529] : 
                               (N877)? mem_q[1892] : 
                               (N879)? mem_q[2255] : 
                               (N881)? mem_q[2618] : 1'b0;
  assign commit_instr_o[438] = (N874)? mem_q[76] : 
                               (N876)? mem_q[439] : 
                               (N878)? mem_q[802] : 
                               (N880)? mem_q[1165] : 
                               (N875)? mem_q[1528] : 
                               (N877)? mem_q[1891] : 
                               (N879)? mem_q[2254] : 
                               (N881)? mem_q[2617] : 1'b0;
  assign commit_instr_o[437] = (N874)? mem_q[75] : 
                               (N876)? mem_q[438] : 
                               (N878)? mem_q[801] : 
                               (N880)? mem_q[1164] : 
                               (N875)? mem_q[1527] : 
                               (N877)? mem_q[1890] : 
                               (N879)? mem_q[2253] : 
                               (N881)? mem_q[2616] : 1'b0;
  assign commit_instr_o[436] = (N874)? mem_q[74] : 
                               (N876)? mem_q[437] : 
                               (N878)? mem_q[800] : 
                               (N880)? mem_q[1163] : 
                               (N875)? mem_q[1526] : 
                               (N877)? mem_q[1889] : 
                               (N879)? mem_q[2252] : 
                               (N881)? mem_q[2615] : 1'b0;
  assign commit_instr_o[435] = (N874)? mem_q[73] : 
                               (N876)? mem_q[436] : 
                               (N878)? mem_q[799] : 
                               (N880)? mem_q[1162] : 
                               (N875)? mem_q[1525] : 
                               (N877)? mem_q[1888] : 
                               (N879)? mem_q[2251] : 
                               (N881)? mem_q[2614] : 1'b0;
  assign commit_instr_o[434] = (N874)? mem_q[72] : 
                               (N876)? mem_q[435] : 
                               (N878)? mem_q[798] : 
                               (N880)? mem_q[1161] : 
                               (N875)? mem_q[1524] : 
                               (N877)? mem_q[1887] : 
                               (N879)? mem_q[2250] : 
                               (N881)? mem_q[2613] : 1'b0;
  assign commit_instr_o[433] = (N874)? mem_q[71] : 
                               (N876)? mem_q[434] : 
                               (N878)? mem_q[797] : 
                               (N880)? mem_q[1160] : 
                               (N875)? mem_q[1523] : 
                               (N877)? mem_q[1886] : 
                               (N879)? mem_q[2249] : 
                               (N881)? mem_q[2612] : 1'b0;
  assign commit_instr_o[432] = (N874)? mem_q[70] : 
                               (N876)? mem_q[433] : 
                               (N878)? mem_q[796] : 
                               (N880)? mem_q[1159] : 
                               (N875)? mem_q[1522] : 
                               (N877)? mem_q[1885] : 
                               (N879)? mem_q[2248] : 
                               (N881)? mem_q[2611] : 1'b0;
  assign commit_instr_o[431] = (N874)? mem_q[69] : 
                               (N876)? mem_q[432] : 
                               (N878)? mem_q[795] : 
                               (N880)? mem_q[1158] : 
                               (N875)? mem_q[1521] : 
                               (N877)? mem_q[1884] : 
                               (N879)? mem_q[2247] : 
                               (N881)? mem_q[2610] : 1'b0;
  assign commit_instr_o[430] = (N874)? mem_q[68] : 
                               (N876)? mem_q[431] : 
                               (N878)? mem_q[794] : 
                               (N880)? mem_q[1157] : 
                               (N875)? mem_q[1520] : 
                               (N877)? mem_q[1883] : 
                               (N879)? mem_q[2246] : 
                               (N881)? mem_q[2609] : 1'b0;
  assign commit_instr_o[429] = (N874)? mem_q[67] : 
                               (N876)? mem_q[430] : 
                               (N878)? mem_q[793] : 
                               (N880)? mem_q[1156] : 
                               (N875)? mem_q[1519] : 
                               (N877)? mem_q[1882] : 
                               (N879)? mem_q[2245] : 
                               (N881)? mem_q[2608] : 1'b0;
  assign commit_instr_o[428] = (N874)? mem_q[66] : 
                               (N876)? mem_q[429] : 
                               (N878)? mem_q[792] : 
                               (N880)? mem_q[1155] : 
                               (N875)? mem_q[1518] : 
                               (N877)? mem_q[1881] : 
                               (N879)? mem_q[2244] : 
                               (N881)? mem_q[2607] : 1'b0;
  assign commit_instr_o[427] = (N874)? mem_q[65] : 
                               (N876)? mem_q[428] : 
                               (N878)? mem_q[791] : 
                               (N880)? mem_q[1154] : 
                               (N875)? mem_q[1517] : 
                               (N877)? mem_q[1880] : 
                               (N879)? mem_q[2243] : 
                               (N881)? mem_q[2606] : 1'b0;
  assign commit_instr_o[426] = (N874)? mem_q[64] : 
                               (N876)? mem_q[427] : 
                               (N878)? mem_q[790] : 
                               (N880)? mem_q[1153] : 
                               (N875)? mem_q[1516] : 
                               (N877)? mem_q[1879] : 
                               (N879)? mem_q[2242] : 
                               (N881)? mem_q[2605] : 1'b0;
  assign commit_instr_o[425] = (N874)? mem_q[63] : 
                               (N876)? mem_q[426] : 
                               (N878)? mem_q[789] : 
                               (N880)? mem_q[1152] : 
                               (N875)? mem_q[1515] : 
                               (N877)? mem_q[1878] : 
                               (N879)? mem_q[2241] : 
                               (N881)? mem_q[2604] : 1'b0;
  assign commit_instr_o[424] = (N874)? mem_q[62] : 
                               (N876)? mem_q[425] : 
                               (N878)? mem_q[788] : 
                               (N880)? mem_q[1151] : 
                               (N875)? mem_q[1514] : 
                               (N877)? mem_q[1877] : 
                               (N879)? mem_q[2240] : 
                               (N881)? mem_q[2603] : 1'b0;
  assign commit_instr_o[423] = (N874)? mem_q[61] : 
                               (N876)? mem_q[424] : 
                               (N878)? mem_q[787] : 
                               (N880)? mem_q[1150] : 
                               (N875)? mem_q[1513] : 
                               (N877)? mem_q[1876] : 
                               (N879)? mem_q[2239] : 
                               (N881)? mem_q[2602] : 1'b0;
  assign commit_instr_o[422] = (N874)? mem_q[60] : 
                               (N876)? mem_q[423] : 
                               (N878)? mem_q[786] : 
                               (N880)? mem_q[1149] : 
                               (N875)? mem_q[1512] : 
                               (N877)? mem_q[1875] : 
                               (N879)? mem_q[2238] : 
                               (N881)? mem_q[2601] : 1'b0;
  assign commit_instr_o[421] = (N874)? mem_q[59] : 
                               (N876)? mem_q[422] : 
                               (N878)? mem_q[785] : 
                               (N880)? mem_q[1148] : 
                               (N875)? mem_q[1511] : 
                               (N877)? mem_q[1874] : 
                               (N879)? mem_q[2237] : 
                               (N881)? mem_q[2600] : 1'b0;
  assign commit_instr_o[420] = (N874)? mem_q[58] : 
                               (N876)? mem_q[421] : 
                               (N878)? mem_q[784] : 
                               (N880)? mem_q[1147] : 
                               (N875)? mem_q[1510] : 
                               (N877)? mem_q[1873] : 
                               (N879)? mem_q[2236] : 
                               (N881)? mem_q[2599] : 1'b0;
  assign commit_instr_o[419] = (N874)? mem_q[57] : 
                               (N876)? mem_q[420] : 
                               (N878)? mem_q[783] : 
                               (N880)? mem_q[1146] : 
                               (N875)? mem_q[1509] : 
                               (N877)? mem_q[1872] : 
                               (N879)? mem_q[2235] : 
                               (N881)? mem_q[2598] : 1'b0;
  assign commit_instr_o[418] = (N874)? mem_q[56] : 
                               (N876)? mem_q[419] : 
                               (N878)? mem_q[782] : 
                               (N880)? mem_q[1145] : 
                               (N875)? mem_q[1508] : 
                               (N877)? mem_q[1871] : 
                               (N879)? mem_q[2234] : 
                               (N881)? mem_q[2597] : 1'b0;
  assign commit_instr_o[417] = (N874)? mem_q[55] : 
                               (N876)? mem_q[418] : 
                               (N878)? mem_q[781] : 
                               (N880)? mem_q[1144] : 
                               (N875)? mem_q[1507] : 
                               (N877)? mem_q[1870] : 
                               (N879)? mem_q[2233] : 
                               (N881)? mem_q[2596] : 1'b0;
  assign commit_instr_o[416] = (N874)? mem_q[54] : 
                               (N876)? mem_q[417] : 
                               (N878)? mem_q[780] : 
                               (N880)? mem_q[1143] : 
                               (N875)? mem_q[1506] : 
                               (N877)? mem_q[1869] : 
                               (N879)? mem_q[2232] : 
                               (N881)? mem_q[2595] : 1'b0;
  assign commit_instr_o[415] = (N874)? mem_q[53] : 
                               (N876)? mem_q[416] : 
                               (N878)? mem_q[779] : 
                               (N880)? mem_q[1142] : 
                               (N875)? mem_q[1505] : 
                               (N877)? mem_q[1868] : 
                               (N879)? mem_q[2231] : 
                               (N881)? mem_q[2594] : 1'b0;
  assign commit_instr_o[414] = (N874)? mem_q[52] : 
                               (N876)? mem_q[415] : 
                               (N878)? mem_q[778] : 
                               (N880)? mem_q[1141] : 
                               (N875)? mem_q[1504] : 
                               (N877)? mem_q[1867] : 
                               (N879)? mem_q[2230] : 
                               (N881)? mem_q[2593] : 1'b0;
  assign commit_instr_o[413] = (N874)? mem_q[51] : 
                               (N876)? mem_q[414] : 
                               (N878)? mem_q[777] : 
                               (N880)? mem_q[1140] : 
                               (N875)? mem_q[1503] : 
                               (N877)? mem_q[1866] : 
                               (N879)? mem_q[2229] : 
                               (N881)? mem_q[2592] : 1'b0;
  assign commit_instr_o[412] = (N874)? mem_q[50] : 
                               (N876)? mem_q[413] : 
                               (N878)? mem_q[776] : 
                               (N880)? mem_q[1139] : 
                               (N875)? mem_q[1502] : 
                               (N877)? mem_q[1865] : 
                               (N879)? mem_q[2228] : 
                               (N881)? mem_q[2591] : 1'b0;
  assign commit_instr_o[411] = (N874)? mem_q[49] : 
                               (N876)? mem_q[412] : 
                               (N878)? mem_q[775] : 
                               (N880)? mem_q[1138] : 
                               (N875)? mem_q[1501] : 
                               (N877)? mem_q[1864] : 
                               (N879)? mem_q[2227] : 
                               (N881)? mem_q[2590] : 1'b0;
  assign commit_instr_o[410] = (N874)? mem_q[48] : 
                               (N876)? mem_q[411] : 
                               (N878)? mem_q[774] : 
                               (N880)? mem_q[1137] : 
                               (N875)? mem_q[1500] : 
                               (N877)? mem_q[1863] : 
                               (N879)? mem_q[2226] : 
                               (N881)? mem_q[2589] : 1'b0;
  assign commit_instr_o[409] = (N874)? mem_q[47] : 
                               (N876)? mem_q[410] : 
                               (N878)? mem_q[773] : 
                               (N880)? mem_q[1136] : 
                               (N875)? mem_q[1499] : 
                               (N877)? mem_q[1862] : 
                               (N879)? mem_q[2225] : 
                               (N881)? mem_q[2588] : 1'b0;
  assign commit_instr_o[408] = (N874)? mem_q[46] : 
                               (N876)? mem_q[409] : 
                               (N878)? mem_q[772] : 
                               (N880)? mem_q[1135] : 
                               (N875)? mem_q[1498] : 
                               (N877)? mem_q[1861] : 
                               (N879)? mem_q[2224] : 
                               (N881)? mem_q[2587] : 1'b0;
  assign commit_instr_o[407] = (N874)? mem_q[45] : 
                               (N876)? mem_q[408] : 
                               (N878)? mem_q[771] : 
                               (N880)? mem_q[1134] : 
                               (N875)? mem_q[1497] : 
                               (N877)? mem_q[1860] : 
                               (N879)? mem_q[2223] : 
                               (N881)? mem_q[2586] : 1'b0;
  assign commit_instr_o[406] = (N874)? mem_q[44] : 
                               (N876)? mem_q[407] : 
                               (N878)? mem_q[770] : 
                               (N880)? mem_q[1133] : 
                               (N875)? mem_q[1496] : 
                               (N877)? mem_q[1859] : 
                               (N879)? mem_q[2222] : 
                               (N881)? mem_q[2585] : 1'b0;
  assign commit_instr_o[405] = (N874)? mem_q[43] : 
                               (N876)? mem_q[406] : 
                               (N878)? mem_q[769] : 
                               (N880)? mem_q[1132] : 
                               (N875)? mem_q[1495] : 
                               (N877)? mem_q[1858] : 
                               (N879)? mem_q[2221] : 
                               (N881)? mem_q[2584] : 1'b0;
  assign commit_instr_o[404] = (N874)? mem_q[42] : 
                               (N876)? mem_q[405] : 
                               (N878)? mem_q[768] : 
                               (N880)? mem_q[1131] : 
                               (N875)? mem_q[1494] : 
                               (N877)? mem_q[1857] : 
                               (N879)? mem_q[2220] : 
                               (N881)? mem_q[2583] : 1'b0;
  assign commit_instr_o[403] = (N874)? mem_q[41] : 
                               (N876)? mem_q[404] : 
                               (N878)? mem_q[767] : 
                               (N880)? mem_q[1130] : 
                               (N875)? mem_q[1493] : 
                               (N877)? mem_q[1856] : 
                               (N879)? mem_q[2219] : 
                               (N881)? mem_q[2582] : 1'b0;
  assign commit_instr_o[402] = (N874)? mem_q[40] : 
                               (N876)? mem_q[403] : 
                               (N878)? mem_q[766] : 
                               (N880)? mem_q[1129] : 
                               (N875)? mem_q[1492] : 
                               (N877)? mem_q[1855] : 
                               (N879)? mem_q[2218] : 
                               (N881)? mem_q[2581] : 1'b0;
  assign commit_instr_o[401] = (N874)? mem_q[39] : 
                               (N876)? mem_q[402] : 
                               (N878)? mem_q[765] : 
                               (N880)? mem_q[1128] : 
                               (N875)? mem_q[1491] : 
                               (N877)? mem_q[1854] : 
                               (N879)? mem_q[2217] : 
                               (N881)? mem_q[2580] : 1'b0;
  assign commit_instr_o[400] = (N874)? mem_q[38] : 
                               (N876)? mem_q[401] : 
                               (N878)? mem_q[764] : 
                               (N880)? mem_q[1127] : 
                               (N875)? mem_q[1490] : 
                               (N877)? mem_q[1853] : 
                               (N879)? mem_q[2216] : 
                               (N881)? mem_q[2579] : 1'b0;
  assign commit_instr_o[399] = (N874)? mem_q[37] : 
                               (N876)? mem_q[400] : 
                               (N878)? mem_q[763] : 
                               (N880)? mem_q[1126] : 
                               (N875)? mem_q[1489] : 
                               (N877)? mem_q[1852] : 
                               (N879)? mem_q[2215] : 
                               (N881)? mem_q[2578] : 1'b0;
  assign commit_instr_o[398] = (N874)? mem_q[36] : 
                               (N876)? mem_q[399] : 
                               (N878)? mem_q[762] : 
                               (N880)? mem_q[1125] : 
                               (N875)? mem_q[1488] : 
                               (N877)? mem_q[1851] : 
                               (N879)? mem_q[2214] : 
                               (N881)? mem_q[2577] : 1'b0;
  assign commit_instr_o[397] = (N874)? mem_q[35] : 
                               (N876)? mem_q[398] : 
                               (N878)? mem_q[761] : 
                               (N880)? mem_q[1124] : 
                               (N875)? mem_q[1487] : 
                               (N877)? mem_q[1850] : 
                               (N879)? mem_q[2213] : 
                               (N881)? mem_q[2576] : 1'b0;
  assign commit_instr_o[396] = (N874)? mem_q[34] : 
                               (N876)? mem_q[397] : 
                               (N878)? mem_q[760] : 
                               (N880)? mem_q[1123] : 
                               (N875)? mem_q[1486] : 
                               (N877)? mem_q[1849] : 
                               (N879)? mem_q[2212] : 
                               (N881)? mem_q[2575] : 1'b0;
  assign commit_instr_o[395] = (N874)? mem_q[33] : 
                               (N876)? mem_q[396] : 
                               (N878)? mem_q[759] : 
                               (N880)? mem_q[1122] : 
                               (N875)? mem_q[1485] : 
                               (N877)? mem_q[1848] : 
                               (N879)? mem_q[2211] : 
                               (N881)? mem_q[2574] : 1'b0;
  assign commit_instr_o[394] = (N874)? mem_q[32] : 
                               (N876)? mem_q[395] : 
                               (N878)? mem_q[758] : 
                               (N880)? mem_q[1121] : 
                               (N875)? mem_q[1484] : 
                               (N877)? mem_q[1847] : 
                               (N879)? mem_q[2210] : 
                               (N881)? mem_q[2573] : 1'b0;
  assign commit_instr_o[393] = (N874)? mem_q[31] : 
                               (N876)? mem_q[394] : 
                               (N878)? mem_q[757] : 
                               (N880)? mem_q[1120] : 
                               (N875)? mem_q[1483] : 
                               (N877)? mem_q[1846] : 
                               (N879)? mem_q[2209] : 
                               (N881)? mem_q[2572] : 1'b0;
  assign commit_instr_o[392] = (N874)? mem_q[30] : 
                               (N876)? mem_q[393] : 
                               (N878)? mem_q[756] : 
                               (N880)? mem_q[1119] : 
                               (N875)? mem_q[1482] : 
                               (N877)? mem_q[1845] : 
                               (N879)? mem_q[2208] : 
                               (N881)? mem_q[2571] : 1'b0;
  assign commit_instr_o[391] = (N874)? mem_q[29] : 
                               (N876)? mem_q[392] : 
                               (N878)? mem_q[755] : 
                               (N880)? mem_q[1118] : 
                               (N875)? mem_q[1481] : 
                               (N877)? mem_q[1844] : 
                               (N879)? mem_q[2207] : 
                               (N881)? mem_q[2570] : 1'b0;
  assign commit_instr_o[390] = (N874)? mem_q[28] : 
                               (N876)? mem_q[391] : 
                               (N878)? mem_q[754] : 
                               (N880)? mem_q[1117] : 
                               (N875)? mem_q[1480] : 
                               (N877)? mem_q[1843] : 
                               (N879)? mem_q[2206] : 
                               (N881)? mem_q[2569] : 1'b0;
  assign commit_instr_o[389] = (N874)? mem_q[27] : 
                               (N876)? mem_q[390] : 
                               (N878)? mem_q[753] : 
                               (N880)? mem_q[1116] : 
                               (N875)? mem_q[1479] : 
                               (N877)? mem_q[1842] : 
                               (N879)? mem_q[2205] : 
                               (N881)? mem_q[2568] : 1'b0;
  assign commit_instr_o[388] = (N874)? mem_q[26] : 
                               (N876)? mem_q[389] : 
                               (N878)? mem_q[752] : 
                               (N880)? mem_q[1115] : 
                               (N875)? mem_q[1478] : 
                               (N877)? mem_q[1841] : 
                               (N879)? mem_q[2204] : 
                               (N881)? mem_q[2567] : 1'b0;
  assign commit_instr_o[387] = (N874)? mem_q[25] : 
                               (N876)? mem_q[388] : 
                               (N878)? mem_q[751] : 
                               (N880)? mem_q[1114] : 
                               (N875)? mem_q[1477] : 
                               (N877)? mem_q[1840] : 
                               (N879)? mem_q[2203] : 
                               (N881)? mem_q[2566] : 1'b0;
  assign commit_instr_o[386] = (N874)? mem_q[24] : 
                               (N876)? mem_q[387] : 
                               (N878)? mem_q[750] : 
                               (N880)? mem_q[1113] : 
                               (N875)? mem_q[1476] : 
                               (N877)? mem_q[1839] : 
                               (N879)? mem_q[2202] : 
                               (N881)? mem_q[2565] : 1'b0;
  assign commit_instr_o[385] = (N874)? mem_q[23] : 
                               (N876)? mem_q[386] : 
                               (N878)? mem_q[749] : 
                               (N880)? mem_q[1112] : 
                               (N875)? mem_q[1475] : 
                               (N877)? mem_q[1838] : 
                               (N879)? mem_q[2201] : 
                               (N881)? mem_q[2564] : 1'b0;
  assign commit_instr_o[384] = (N874)? mem_q[22] : 
                               (N876)? mem_q[385] : 
                               (N878)? mem_q[748] : 
                               (N880)? mem_q[1111] : 
                               (N875)? mem_q[1474] : 
                               (N877)? mem_q[1837] : 
                               (N879)? mem_q[2200] : 
                               (N881)? mem_q[2563] : 1'b0;
  assign commit_instr_o[383] = (N874)? mem_q[21] : 
                               (N876)? mem_q[384] : 
                               (N878)? mem_q[747] : 
                               (N880)? mem_q[1110] : 
                               (N875)? mem_q[1473] : 
                               (N877)? mem_q[1836] : 
                               (N879)? mem_q[2199] : 
                               (N881)? mem_q[2562] : 1'b0;
  assign commit_instr_o[382] = (N874)? mem_q[20] : 
                               (N876)? mem_q[383] : 
                               (N878)? mem_q[746] : 
                               (N880)? mem_q[1109] : 
                               (N875)? mem_q[1472] : 
                               (N877)? mem_q[1835] : 
                               (N879)? mem_q[2198] : 
                               (N881)? mem_q[2561] : 1'b0;
  assign commit_instr_o[381] = (N874)? mem_q[19] : 
                               (N876)? mem_q[382] : 
                               (N878)? mem_q[745] : 
                               (N880)? mem_q[1108] : 
                               (N875)? mem_q[1471] : 
                               (N877)? mem_q[1834] : 
                               (N879)? mem_q[2197] : 
                               (N881)? mem_q[2560] : 1'b0;
  assign commit_instr_o[380] = (N874)? mem_q[18] : 
                               (N876)? mem_q[381] : 
                               (N878)? mem_q[744] : 
                               (N880)? mem_q[1107] : 
                               (N875)? mem_q[1470] : 
                               (N877)? mem_q[1833] : 
                               (N879)? mem_q[2196] : 
                               (N881)? mem_q[2559] : 1'b0;
  assign commit_instr_o[379] = (N874)? mem_q[17] : 
                               (N876)? mem_q[380] : 
                               (N878)? mem_q[743] : 
                               (N880)? mem_q[1106] : 
                               (N875)? mem_q[1469] : 
                               (N877)? mem_q[1832] : 
                               (N879)? mem_q[2195] : 
                               (N881)? mem_q[2558] : 1'b0;
  assign commit_instr_o[378] = (N874)? mem_q[16] : 
                               (N876)? mem_q[379] : 
                               (N878)? mem_q[742] : 
                               (N880)? mem_q[1105] : 
                               (N875)? mem_q[1468] : 
                               (N877)? mem_q[1831] : 
                               (N879)? mem_q[2194] : 
                               (N881)? mem_q[2557] : 1'b0;
  assign commit_instr_o[377] = (N874)? mem_q[15] : 
                               (N876)? mem_q[378] : 
                               (N878)? mem_q[741] : 
                               (N880)? mem_q[1104] : 
                               (N875)? mem_q[1467] : 
                               (N877)? mem_q[1830] : 
                               (N879)? mem_q[2193] : 
                               (N881)? mem_q[2556] : 1'b0;
  assign commit_instr_o[376] = (N874)? mem_q[14] : 
                               (N876)? mem_q[377] : 
                               (N878)? mem_q[740] : 
                               (N880)? mem_q[1103] : 
                               (N875)? mem_q[1466] : 
                               (N877)? mem_q[1829] : 
                               (N879)? mem_q[2192] : 
                               (N881)? mem_q[2555] : 1'b0;
  assign commit_instr_o[375] = (N874)? mem_q[13] : 
                               (N876)? mem_q[376] : 
                               (N878)? mem_q[739] : 
                               (N880)? mem_q[1102] : 
                               (N875)? mem_q[1465] : 
                               (N877)? mem_q[1828] : 
                               (N879)? mem_q[2191] : 
                               (N881)? mem_q[2554] : 1'b0;
  assign commit_instr_o[374] = (N874)? mem_q[12] : 
                               (N876)? mem_q[375] : 
                               (N878)? mem_q[738] : 
                               (N880)? mem_q[1101] : 
                               (N875)? mem_q[1464] : 
                               (N877)? mem_q[1827] : 
                               (N879)? mem_q[2190] : 
                               (N881)? mem_q[2553] : 1'b0;
  assign commit_instr_o[373] = (N874)? mem_q[11] : 
                               (N876)? mem_q[374] : 
                               (N878)? mem_q[737] : 
                               (N880)? mem_q[1100] : 
                               (N875)? mem_q[1463] : 
                               (N877)? mem_q[1826] : 
                               (N879)? mem_q[2189] : 
                               (N881)? mem_q[2552] : 1'b0;
  assign commit_instr_o[372] = (N874)? mem_q[10] : 
                               (N876)? mem_q[373] : 
                               (N878)? mem_q[736] : 
                               (N880)? mem_q[1099] : 
                               (N875)? mem_q[1462] : 
                               (N877)? mem_q[1825] : 
                               (N879)? mem_q[2188] : 
                               (N881)? mem_q[2551] : 1'b0;
  assign commit_instr_o[371] = (N874)? mem_q[9] : 
                               (N876)? mem_q[372] : 
                               (N878)? mem_q[735] : 
                               (N880)? mem_q[1098] : 
                               (N875)? mem_q[1461] : 
                               (N877)? mem_q[1824] : 
                               (N879)? mem_q[2187] : 
                               (N881)? mem_q[2550] : 1'b0;
  assign commit_instr_o[370] = (N874)? mem_q[8] : 
                               (N876)? mem_q[371] : 
                               (N878)? mem_q[734] : 
                               (N880)? mem_q[1097] : 
                               (N875)? mem_q[1460] : 
                               (N877)? mem_q[1823] : 
                               (N879)? mem_q[2186] : 
                               (N881)? mem_q[2549] : 1'b0;
  assign commit_instr_o[369] = (N874)? mem_q[7] : 
                               (N876)? mem_q[370] : 
                               (N878)? mem_q[733] : 
                               (N880)? mem_q[1096] : 
                               (N875)? mem_q[1459] : 
                               (N877)? mem_q[1822] : 
                               (N879)? mem_q[2185] : 
                               (N881)? mem_q[2548] : 1'b0;
  assign commit_instr_o[368] = (N874)? mem_q[6] : 
                               (N876)? mem_q[369] : 
                               (N878)? mem_q[732] : 
                               (N880)? mem_q[1095] : 
                               (N875)? mem_q[1458] : 
                               (N877)? mem_q[1821] : 
                               (N879)? mem_q[2184] : 
                               (N881)? mem_q[2547] : 1'b0;
  assign commit_instr_o[367] = (N874)? mem_q[5] : 
                               (N876)? mem_q[368] : 
                               (N878)? mem_q[731] : 
                               (N880)? mem_q[1094] : 
                               (N875)? mem_q[1457] : 
                               (N877)? mem_q[1820] : 
                               (N879)? mem_q[2183] : 
                               (N881)? mem_q[2546] : 1'b0;
  assign commit_instr_o[366] = (N874)? mem_q[4] : 
                               (N876)? mem_q[367] : 
                               (N878)? mem_q[730] : 
                               (N880)? mem_q[1093] : 
                               (N875)? mem_q[1456] : 
                               (N877)? mem_q[1819] : 
                               (N879)? mem_q[2182] : 
                               (N881)? mem_q[2545] : 1'b0;
  assign commit_instr_o[365] = (N874)? mem_q[3] : 
                               (N876)? mem_q[366] : 
                               (N878)? mem_q[729] : 
                               (N880)? mem_q[1092] : 
                               (N875)? mem_q[1455] : 
                               (N877)? mem_q[1818] : 
                               (N879)? mem_q[2181] : 
                               (N881)? mem_q[2544] : 1'b0;
  assign commit_instr_o[364] = (N874)? mem_q[2] : 
                               (N876)? mem_q[365] : 
                               (N878)? mem_q[728] : 
                               (N880)? mem_q[1091] : 
                               (N875)? mem_q[1454] : 
                               (N877)? mem_q[1817] : 
                               (N879)? mem_q[2180] : 
                               (N881)? mem_q[2543] : 1'b0;
  assign commit_instr_o[363] = (N874)? mem_q[1] : 
                               (N876)? mem_q[364] : 
                               (N878)? mem_q[727] : 
                               (N880)? mem_q[1090] : 
                               (N875)? mem_q[1453] : 
                               (N877)? mem_q[1816] : 
                               (N879)? mem_q[2179] : 
                               (N881)? mem_q[2542] : 1'b0;
  assign commit_instr_o[362] = (N874)? mem_q[0] : 
                               (N876)? mem_q[363] : 
                               (N878)? mem_q[726] : 
                               (N880)? mem_q[1089] : 
                               (N875)? mem_q[1452] : 
                               (N877)? mem_q[1815] : 
                               (N879)? mem_q[2178] : 
                               (N881)? mem_q[2541] : 1'b0;
  assign N5901 = (N5893)? N4072 : 
                 (N5895)? N4331 : 
                 (N5897)? N4590 : 
                 (N5899)? N4849 : 
                 (N5894)? N5108 : 
                 (N5896)? N5367 : 
                 (N5898)? N5626 : 
                 (N5900)? N5885 : 1'b0;
  assign N6952 = (N5893)? mem_n[294] : 
                 (N5895)? mem_n[657] : 
                 (N5897)? mem_n[1020] : 
                 (N5899)? mem_n[1383] : 
                 (N5894)? mem_n[1746] : 
                 (N5896)? mem_n[2109] : 
                 (N5898)? mem_n[2472] : 
                 (N5900)? mem_n[2835] : 1'b0;
  assign N6953 = (N5893)? mem_n[293] : 
                 (N5895)? mem_n[656] : 
                 (N5897)? mem_n[1019] : 
                 (N5899)? mem_n[1382] : 
                 (N5894)? mem_n[1745] : 
                 (N5896)? mem_n[2108] : 
                 (N5898)? mem_n[2471] : 
                 (N5900)? mem_n[2834] : 1'b0;
  assign N6954 = (N5893)? mem_n[292] : 
                 (N5895)? mem_n[655] : 
                 (N5897)? mem_n[1018] : 
                 (N5899)? mem_n[1381] : 
                 (N5894)? mem_n[1744] : 
                 (N5896)? mem_n[2107] : 
                 (N5898)? mem_n[2470] : 
                 (N5900)? mem_n[2833] : 1'b0;
  assign N6955 = (N5893)? mem_n[291] : 
                 (N5895)? mem_n[654] : 
                 (N5897)? mem_n[1017] : 
                 (N5899)? mem_n[1380] : 
                 (N5894)? mem_n[1743] : 
                 (N5896)? mem_n[2106] : 
                 (N5898)? mem_n[2469] : 
                 (N5900)? mem_n[2832] : 1'b0;
  assign N7992 = N6952 | N7989;
  assign N7993 = N7990 | N7991;
  assign N7994 = N7992 | N7993;
  assign N7996 = N7995 | N6953;
  assign N7997 = N6954 | N6955;
  assign N7998 = N7996 | N7997;
  assign N12136 = (N12128)? N4072 : 
                  (N12130)? N4331 : 
                  (N12132)? N4590 : 
                  (N12134)? N4849 : 
                  (N12129)? N5108 : 
                  (N12131)? N5367 : 
                  (N12133)? N5626 : 
                  (N12135)? N5885 : 1'b0;
  assign N13187 = (N12128)? mem_n[294] : 
                  (N12130)? mem_n[657] : 
                  (N12132)? mem_n[1020] : 
                  (N12134)? mem_n[1383] : 
                  (N12129)? mem_n[1746] : 
                  (N12131)? mem_n[2109] : 
                  (N12133)? mem_n[2472] : 
                  (N12135)? mem_n[2835] : 1'b0;
  assign N13188 = (N12128)? mem_n[293] : 
                  (N12130)? mem_n[656] : 
                  (N12132)? mem_n[1019] : 
                  (N12134)? mem_n[1382] : 
                  (N12129)? mem_n[1745] : 
                  (N12131)? mem_n[2108] : 
                  (N12133)? mem_n[2471] : 
                  (N12135)? mem_n[2834] : 1'b0;
  assign N13189 = (N12128)? mem_n[292] : 
                  (N12130)? mem_n[655] : 
                  (N12132)? mem_n[1018] : 
                  (N12134)? mem_n[1381] : 
                  (N12129)? mem_n[1744] : 
                  (N12131)? mem_n[2107] : 
                  (N12133)? mem_n[2470] : 
                  (N12135)? mem_n[2833] : 1'b0;
  assign N13190 = (N12128)? mem_n[291] : 
                  (N12130)? mem_n[654] : 
                  (N12132)? mem_n[1017] : 
                  (N12134)? mem_n[1380] : 
                  (N12129)? mem_n[1743] : 
                  (N12131)? mem_n[2106] : 
                  (N12133)? mem_n[2469] : 
                  (N12135)? mem_n[2832] : 1'b0;
  assign N14227 = N13187 | N14224;
  assign N14228 = N14225 | N14226;
  assign N14229 = N14227 | N14228;
  assign N14231 = N14230 | N13188;
  assign N14232 = N13189 | N13190;
  assign N14233 = N14231 | N14232;
  assign N18371 = (N18363)? N4072 : 
                  (N18365)? N4331 : 
                  (N18367)? N4590 : 
                  (N18369)? N4849 : 
                  (N18364)? N5108 : 
                  (N18366)? N5367 : 
                  (N18368)? N5626 : 
                  (N18370)? N5885 : 1'b0;
  assign N19422 = (N18363)? mem_n[294] : 
                  (N18365)? mem_n[657] : 
                  (N18367)? mem_n[1020] : 
                  (N18369)? mem_n[1383] : 
                  (N18364)? mem_n[1746] : 
                  (N18366)? mem_n[2109] : 
                  (N18368)? mem_n[2472] : 
                  (N18370)? mem_n[2835] : 1'b0;
  assign N19423 = (N18363)? mem_n[293] : 
                  (N18365)? mem_n[656] : 
                  (N18367)? mem_n[1019] : 
                  (N18369)? mem_n[1382] : 
                  (N18364)? mem_n[1745] : 
                  (N18366)? mem_n[2108] : 
                  (N18368)? mem_n[2471] : 
                  (N18370)? mem_n[2834] : 1'b0;
  assign N19424 = (N18363)? mem_n[292] : 
                  (N18365)? mem_n[655] : 
                  (N18367)? mem_n[1018] : 
                  (N18369)? mem_n[1381] : 
                  (N18364)? mem_n[1744] : 
                  (N18366)? mem_n[2107] : 
                  (N18368)? mem_n[2470] : 
                  (N18370)? mem_n[2833] : 1'b0;
  assign N19425 = (N18363)? mem_n[291] : 
                  (N18365)? mem_n[654] : 
                  (N18367)? mem_n[1017] : 
                  (N18369)? mem_n[1380] : 
                  (N18364)? mem_n[1743] : 
                  (N18366)? mem_n[2106] : 
                  (N18368)? mem_n[2469] : 
                  (N18370)? mem_n[2832] : 1'b0;
  assign N20462 = N19422 | N20459;
  assign N20463 = N20460 | N20461;
  assign N20464 = N20462 | N20463;
  assign N20466 = N20465 | N19423;
  assign N20467 = N19424 | N19425;
  assign N20468 = N20466 | N20467;
  assign N24606 = (N24598)? N4072 : 
                  (N24600)? N4331 : 
                  (N24602)? N4590 : 
                  (N24604)? N4849 : 
                  (N24599)? N5108 : 
                  (N24601)? N5367 : 
                  (N24603)? N5626 : 
                  (N24605)? N5885 : 1'b0;
  assign N25657 = (N24598)? mem_n[294] : 
                  (N24600)? mem_n[657] : 
                  (N24602)? mem_n[1020] : 
                  (N24604)? mem_n[1383] : 
                  (N24599)? mem_n[1746] : 
                  (N24601)? mem_n[2109] : 
                  (N24603)? mem_n[2472] : 
                  (N24605)? mem_n[2835] : 1'b0;
  assign N25658 = (N24598)? mem_n[293] : 
                  (N24600)? mem_n[656] : 
                  (N24602)? mem_n[1019] : 
                  (N24604)? mem_n[1382] : 
                  (N24599)? mem_n[1745] : 
                  (N24601)? mem_n[2108] : 
                  (N24603)? mem_n[2471] : 
                  (N24605)? mem_n[2834] : 1'b0;
  assign N25659 = (N24598)? mem_n[292] : 
                  (N24600)? mem_n[655] : 
                  (N24602)? mem_n[1018] : 
                  (N24604)? mem_n[1381] : 
                  (N24599)? mem_n[1744] : 
                  (N24601)? mem_n[2107] : 
                  (N24603)? mem_n[2470] : 
                  (N24605)? mem_n[2833] : 1'b0;
  assign N25660 = (N24598)? mem_n[291] : 
                  (N24600)? mem_n[654] : 
                  (N24602)? mem_n[1017] : 
                  (N24604)? mem_n[1380] : 
                  (N24599)? mem_n[1743] : 
                  (N24601)? mem_n[2106] : 
                  (N24603)? mem_n[2469] : 
                  (N24605)? mem_n[2832] : 1'b0;
  assign N26697 = N25657 | N26694;
  assign N26698 = N26695 | N26696;
  assign N26699 = N26697 | N26698;
  assign N26701 = N26700 | N25658;
  assign N26702 = N25659 | N25660;
  assign N26703 = N26701 | N26702;
  assign N33732 = mem_q[271:266] == rs1_i;
  assign N33735 = mem_q[271:266] == rs2_i;
  assign N33737 = mem_q[271:266] == rs3_i;
  assign N34077 = mem_q[634:629] == rs1_i;
  assign N34080 = mem_q[634:629] == rs2_i;
  assign N34082 = mem_q[634:629] == rs3_i;
  assign N34422 = mem_q[997:992] == rs1_i;
  assign N34425 = mem_q[997:992] == rs2_i;
  assign N34427 = mem_q[997:992] == rs3_i;
  assign N34767 = mem_q[1360:1355] == rs1_i;
  assign N34770 = mem_q[1360:1355] == rs2_i;
  assign N34772 = mem_q[1360:1355] == rs3_i;
  assign N35112 = mem_q[1723:1718] == rs1_i;
  assign N35115 = mem_q[1723:1718] == rs2_i;
  assign N35117 = mem_q[1723:1718] == rs3_i;
  assign N35457 = mem_q[2086:2081] == rs1_i;
  assign N35460 = mem_q[2086:2081] == rs2_i;
  assign N35462 = mem_q[2086:2081] == rs3_i;
  assign N35802 = mem_q[2449:2444] == rs1_i;
  assign N35805 = mem_q[2449:2444] == rs2_i;
  assign N35807 = mem_q[2449:2444] == rs3_i;
  assign N36147 = mem_q[2812:2807] == rs1_i;
  assign N36150 = mem_q[2812:2807] == rs2_i;
  assign N36152 = mem_q[2812:2807] == rs3_i;
  assign N36491 = (N5893)? mem_q[271] : 
                  (N5895)? mem_q[634] : 
                  (N5897)? mem_q[997] : 
                  (N5899)? mem_q[1360] : 
                  (N5894)? mem_q[1723] : 
                  (N5896)? mem_q[2086] : 
                  (N5898)? mem_q[2449] : 
                  (N5900)? mem_q[2812] : 1'b0;
  assign N36492 = (N5893)? mem_q[270] : 
                  (N5895)? mem_q[633] : 
                  (N5897)? mem_q[996] : 
                  (N5899)? mem_q[1359] : 
                  (N5894)? mem_q[1722] : 
                  (N5896)? mem_q[2085] : 
                  (N5898)? mem_q[2448] : 
                  (N5900)? mem_q[2811] : 1'b0;
  assign N36493 = (N5893)? mem_q[269] : 
                  (N5895)? mem_q[632] : 
                  (N5897)? mem_q[995] : 
                  (N5899)? mem_q[1358] : 
                  (N5894)? mem_q[1721] : 
                  (N5896)? mem_q[2084] : 
                  (N5898)? mem_q[2447] : 
                  (N5900)? mem_q[2810] : 1'b0;
  assign N36494 = (N5893)? mem_q[268] : 
                  (N5895)? mem_q[631] : 
                  (N5897)? mem_q[994] : 
                  (N5899)? mem_q[1357] : 
                  (N5894)? mem_q[1720] : 
                  (N5896)? mem_q[2083] : 
                  (N5898)? mem_q[2446] : 
                  (N5900)? mem_q[2809] : 1'b0;
  assign N36495 = (N5893)? mem_q[267] : 
                  (N5895)? mem_q[630] : 
                  (N5897)? mem_q[993] : 
                  (N5899)? mem_q[1356] : 
                  (N5894)? mem_q[1719] : 
                  (N5896)? mem_q[2082] : 
                  (N5898)? mem_q[2445] : 
                  (N5900)? mem_q[2808] : 1'b0;
  assign N36496 = (N5893)? mem_q[266] : 
                  (N5895)? mem_q[629] : 
                  (N5897)? mem_q[992] : 
                  (N5899)? mem_q[1355] : 
                  (N5894)? mem_q[1718] : 
                  (N5896)? mem_q[2081] : 
                  (N5898)? mem_q[2444] : 
                  (N5900)? mem_q[2807] : 1'b0;
  assign N36498 = { N36491, N36492, N36493, N36494, N36495, N36496 } == rs1_i;
  assign N36567 = { N36491, N36492, N36493, N36494, N36495, N36496 } == rs2_i;
  assign N36638 = { N36491, N36492, N36493, N36494, N36495, N36496 } == rs3_i;
  assign N36648 = (N12128)? mem_q[271] : 
                  (N12130)? mem_q[634] : 
                  (N12132)? mem_q[997] : 
                  (N12134)? mem_q[1360] : 
                  (N12129)? mem_q[1723] : 
                  (N12131)? mem_q[2086] : 
                  (N12133)? mem_q[2449] : 
                  (N12135)? mem_q[2812] : 1'b0;
  assign N36649 = (N12128)? mem_q[270] : 
                  (N12130)? mem_q[633] : 
                  (N12132)? mem_q[996] : 
                  (N12134)? mem_q[1359] : 
                  (N12129)? mem_q[1722] : 
                  (N12131)? mem_q[2085] : 
                  (N12133)? mem_q[2448] : 
                  (N12135)? mem_q[2811] : 1'b0;
  assign N36650 = (N12128)? mem_q[269] : 
                  (N12130)? mem_q[632] : 
                  (N12132)? mem_q[995] : 
                  (N12134)? mem_q[1358] : 
                  (N12129)? mem_q[1721] : 
                  (N12131)? mem_q[2084] : 
                  (N12133)? mem_q[2447] : 
                  (N12135)? mem_q[2810] : 1'b0;
  assign N36651 = (N12128)? mem_q[268] : 
                  (N12130)? mem_q[631] : 
                  (N12132)? mem_q[994] : 
                  (N12134)? mem_q[1357] : 
                  (N12129)? mem_q[1720] : 
                  (N12131)? mem_q[2083] : 
                  (N12133)? mem_q[2446] : 
                  (N12135)? mem_q[2809] : 1'b0;
  assign N36652 = (N12128)? mem_q[267] : 
                  (N12130)? mem_q[630] : 
                  (N12132)? mem_q[993] : 
                  (N12134)? mem_q[1356] : 
                  (N12129)? mem_q[1719] : 
                  (N12131)? mem_q[2082] : 
                  (N12133)? mem_q[2445] : 
                  (N12135)? mem_q[2808] : 1'b0;
  assign N36653 = (N12128)? mem_q[266] : 
                  (N12130)? mem_q[629] : 
                  (N12132)? mem_q[992] : 
                  (N12134)? mem_q[1355] : 
                  (N12129)? mem_q[1718] : 
                  (N12131)? mem_q[2081] : 
                  (N12133)? mem_q[2444] : 
                  (N12135)? mem_q[2807] : 1'b0;
  assign N36655 = { N36648, N36649, N36650, N36651, N36652, N36653 } == rs1_i;
  assign N36726 = { N36648, N36649, N36650, N36651, N36652, N36653 } == rs2_i;
  assign N36797 = { N36648, N36649, N36650, N36651, N36652, N36653 } == rs3_i;
  assign N36807 = (N18363)? mem_q[271] : 
                  (N18365)? mem_q[634] : 
                  (N18367)? mem_q[997] : 
                  (N18369)? mem_q[1360] : 
                  (N18364)? mem_q[1723] : 
                  (N18366)? mem_q[2086] : 
                  (N18368)? mem_q[2449] : 
                  (N18370)? mem_q[2812] : 1'b0;
  assign N36808 = (N18363)? mem_q[270] : 
                  (N18365)? mem_q[633] : 
                  (N18367)? mem_q[996] : 
                  (N18369)? mem_q[1359] : 
                  (N18364)? mem_q[1722] : 
                  (N18366)? mem_q[2085] : 
                  (N18368)? mem_q[2448] : 
                  (N18370)? mem_q[2811] : 1'b0;
  assign N36809 = (N18363)? mem_q[269] : 
                  (N18365)? mem_q[632] : 
                  (N18367)? mem_q[995] : 
                  (N18369)? mem_q[1358] : 
                  (N18364)? mem_q[1721] : 
                  (N18366)? mem_q[2084] : 
                  (N18368)? mem_q[2447] : 
                  (N18370)? mem_q[2810] : 1'b0;
  assign N36810 = (N18363)? mem_q[268] : 
                  (N18365)? mem_q[631] : 
                  (N18367)? mem_q[994] : 
                  (N18369)? mem_q[1357] : 
                  (N18364)? mem_q[1720] : 
                  (N18366)? mem_q[2083] : 
                  (N18368)? mem_q[2446] : 
                  (N18370)? mem_q[2809] : 1'b0;
  assign N36811 = (N18363)? mem_q[267] : 
                  (N18365)? mem_q[630] : 
                  (N18367)? mem_q[993] : 
                  (N18369)? mem_q[1356] : 
                  (N18364)? mem_q[1719] : 
                  (N18366)? mem_q[2082] : 
                  (N18368)? mem_q[2445] : 
                  (N18370)? mem_q[2808] : 1'b0;
  assign N36812 = (N18363)? mem_q[266] : 
                  (N18365)? mem_q[629] : 
                  (N18367)? mem_q[992] : 
                  (N18369)? mem_q[1355] : 
                  (N18364)? mem_q[1718] : 
                  (N18366)? mem_q[2081] : 
                  (N18368)? mem_q[2444] : 
                  (N18370)? mem_q[2807] : 1'b0;
  assign N36814 = { N36807, N36808, N36809, N36810, N36811, N36812 } == rs1_i;
  assign N36885 = { N36807, N36808, N36809, N36810, N36811, N36812 } == rs2_i;
  assign N36956 = { N36807, N36808, N36809, N36810, N36811, N36812 } == rs3_i;
  assign N36966 = (N24598)? mem_q[271] : 
                  (N24600)? mem_q[634] : 
                  (N24602)? mem_q[997] : 
                  (N24604)? mem_q[1360] : 
                  (N24599)? mem_q[1723] : 
                  (N24601)? mem_q[2086] : 
                  (N24603)? mem_q[2449] : 
                  (N24605)? mem_q[2812] : 1'b0;
  assign N36967 = (N24598)? mem_q[270] : 
                  (N24600)? mem_q[633] : 
                  (N24602)? mem_q[996] : 
                  (N24604)? mem_q[1359] : 
                  (N24599)? mem_q[1722] : 
                  (N24601)? mem_q[2085] : 
                  (N24603)? mem_q[2448] : 
                  (N24605)? mem_q[2811] : 1'b0;
  assign N36968 = (N24598)? mem_q[269] : 
                  (N24600)? mem_q[632] : 
                  (N24602)? mem_q[995] : 
                  (N24604)? mem_q[1358] : 
                  (N24599)? mem_q[1721] : 
                  (N24601)? mem_q[2084] : 
                  (N24603)? mem_q[2447] : 
                  (N24605)? mem_q[2810] : 1'b0;
  assign N36969 = (N24598)? mem_q[268] : 
                  (N24600)? mem_q[631] : 
                  (N24602)? mem_q[994] : 
                  (N24604)? mem_q[1357] : 
                  (N24599)? mem_q[1720] : 
                  (N24601)? mem_q[2083] : 
                  (N24603)? mem_q[2446] : 
                  (N24605)? mem_q[2809] : 1'b0;
  assign N36970 = (N24598)? mem_q[267] : 
                  (N24600)? mem_q[630] : 
                  (N24602)? mem_q[993] : 
                  (N24604)? mem_q[1356] : 
                  (N24599)? mem_q[1719] : 
                  (N24601)? mem_q[2082] : 
                  (N24603)? mem_q[2445] : 
                  (N24605)? mem_q[2808] : 1'b0;
  assign N36971 = (N24598)? mem_q[266] : 
                  (N24600)? mem_q[629] : 
                  (N24602)? mem_q[992] : 
                  (N24604)? mem_q[1355] : 
                  (N24599)? mem_q[1718] : 
                  (N24601)? mem_q[2081] : 
                  (N24603)? mem_q[2444] : 
                  (N24605)? mem_q[2807] : 1'b0;
  assign N36973 = { N36966, N36967, N36968, N36969, N36970, N36971 } == rs1_i;
  assign N37044 = { N36966, N36967, N36968, N36969, N36970, N36971 } == rs2_i;
  assign N37114 = { N36966, N36967, N36968, N36969, N36970, N36971 } == rs3_i;

  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      issue_instr_o[297] <= 1'b0;
    end else if(N38661) begin
      issue_instr_o[297] <= issue_pointer_n[2];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      issue_instr_o[296] <= 1'b0;
    end else if(N38661) begin
      issue_instr_o[296] <= issue_pointer_n[1];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      issue_instr_o[295] <= 1'b0;
    end else if(N38661) begin
      issue_instr_o[295] <= issue_pointer_n[0];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2903] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2903] <= mem_n[2903];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2902] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2902] <= mem_n[2902];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2901] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2901] <= mem_n[2901];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2900] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2900] <= mem_n[2900];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2899] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2899] <= mem_n[2899];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2898] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2898] <= mem_n[2898];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2897] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2897] <= mem_n[2897];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2896] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2896] <= mem_n[2896];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2895] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2895] <= mem_n[2895];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2894] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2894] <= mem_n[2894];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2893] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2893] <= mem_n[2893];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2892] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2892] <= mem_n[2892];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2891] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2891] <= mem_n[2891];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2890] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2890] <= mem_n[2890];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2889] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2889] <= mem_n[2889];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2888] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2888] <= mem_n[2888];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2887] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2887] <= mem_n[2887];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2886] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2886] <= mem_n[2886];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2885] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2885] <= mem_n[2885];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2884] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2884] <= mem_n[2884];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2883] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2883] <= mem_n[2883];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2882] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2882] <= mem_n[2882];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2881] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2881] <= mem_n[2881];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2880] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2880] <= mem_n[2880];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2879] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2879] <= mem_n[2879];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2878] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2878] <= mem_n[2878];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2877] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2877] <= mem_n[2877];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2876] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2876] <= mem_n[2876];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2875] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2875] <= mem_n[2875];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2874] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2874] <= mem_n[2874];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2873] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2873] <= mem_n[2873];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2872] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2872] <= mem_n[2872];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2871] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2871] <= mem_n[2871];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2870] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2870] <= mem_n[2870];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2869] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2869] <= mem_n[2869];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2868] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2868] <= mem_n[2868];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2867] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2867] <= mem_n[2867];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2866] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2866] <= mem_n[2866];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2865] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2865] <= mem_n[2865];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2864] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2864] <= mem_n[2864];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2863] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2863] <= mem_n[2863];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2862] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2862] <= mem_n[2862];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2861] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2861] <= mem_n[2861];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2860] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2860] <= mem_n[2860];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2859] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2859] <= mem_n[2859];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2858] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2858] <= mem_n[2858];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2857] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2857] <= mem_n[2857];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2856] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2856] <= mem_n[2856];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2855] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2855] <= mem_n[2855];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2854] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2854] <= mem_n[2854];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2853] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2853] <= mem_n[2853];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2852] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2852] <= mem_n[2852];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2851] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2851] <= mem_n[2851];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2850] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2850] <= mem_n[2850];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2849] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2849] <= mem_n[2849];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2848] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2848] <= mem_n[2848];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2847] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2847] <= mem_n[2847];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2846] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2846] <= mem_n[2846];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2845] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2845] <= mem_n[2845];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2844] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2844] <= mem_n[2844];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2843] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2843] <= mem_n[2843];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2842] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2842] <= mem_n[2842];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2841] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2841] <= mem_n[2841];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2840] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2840] <= mem_n[2840];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2839] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2839] <= mem_n[2839];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2838] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2838] <= mem_n[2838];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2837] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2837] <= mem_n[2837];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2836] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2836] <= mem_n[2836];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2835] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2835] <= mem_n[2835];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2834] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2834] <= mem_n[2834];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2833] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2833] <= mem_n[2833];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2832] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2832] <= mem_n[2832];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2831] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2831] <= mem_n[2831];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2830] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2830] <= mem_n[2830];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2829] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2829] <= mem_n[2829];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2828] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2828] <= mem_n[2828];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2827] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2827] <= mem_n[2827];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2826] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2826] <= mem_n[2826];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2825] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2825] <= mem_n[2825];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2824] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2824] <= mem_n[2824];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2823] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2823] <= mem_n[2823];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2822] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2822] <= mem_n[2822];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2821] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2821] <= mem_n[2821];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2820] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2820] <= mem_n[2820];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2819] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2819] <= mem_n[2819];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2818] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2818] <= mem_n[2818];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2817] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2817] <= mem_n[2817];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2816] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2816] <= mem_n[2816];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2815] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2815] <= mem_n[2815];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2814] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2814] <= mem_n[2814];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2813] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2813] <= mem_n[2813];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2812] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2812] <= mem_n[2812];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2811] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2811] <= mem_n[2811];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2810] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2810] <= mem_n[2810];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2809] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2809] <= mem_n[2809];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2808] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2808] <= mem_n[2808];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2807] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2807] <= mem_n[2807];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2806] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2806] <= mem_n[2806];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2805] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2805] <= mem_n[2805];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2804] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2804] <= mem_n[2804];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2803] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2803] <= mem_n[2803];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2802] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2802] <= mem_n[2802];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2801] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2801] <= mem_n[2801];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2800] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2800] <= mem_n[2800];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2799] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2799] <= mem_n[2799];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2798] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2798] <= mem_n[2798];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2797] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2797] <= mem_n[2797];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2796] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2796] <= mem_n[2796];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2795] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2795] <= mem_n[2795];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2794] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2794] <= mem_n[2794];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2793] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2793] <= mem_n[2793];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2792] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2792] <= mem_n[2792];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2791] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2791] <= mem_n[2791];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2790] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2790] <= mem_n[2790];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2789] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2789] <= mem_n[2789];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2788] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2788] <= mem_n[2788];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2787] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2787] <= mem_n[2787];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2786] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2786] <= mem_n[2786];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2785] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2785] <= mem_n[2785];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2784] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2784] <= mem_n[2784];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2783] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2783] <= mem_n[2783];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2782] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2782] <= mem_n[2782];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2781] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2781] <= mem_n[2781];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2780] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2780] <= mem_n[2780];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2779] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2779] <= mem_n[2779];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2778] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2778] <= mem_n[2778];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2777] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2777] <= mem_n[2777];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2776] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2776] <= mem_n[2776];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2775] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2775] <= mem_n[2775];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2774] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2774] <= mem_n[2774];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2773] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2773] <= mem_n[2773];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2772] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2772] <= mem_n[2772];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2771] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2771] <= mem_n[2771];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2770] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2770] <= mem_n[2770];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2769] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2769] <= mem_n[2769];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2768] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2768] <= mem_n[2768];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2767] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2767] <= mem_n[2767];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2766] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2766] <= mem_n[2766];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2765] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2765] <= mem_n[2765];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2764] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2764] <= mem_n[2764];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2763] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2763] <= mem_n[2763];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2762] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2762] <= mem_n[2762];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2761] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2761] <= mem_n[2761];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2760] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2760] <= mem_n[2760];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2759] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2759] <= mem_n[2759];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2758] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2758] <= mem_n[2758];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2757] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2757] <= mem_n[2757];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2756] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2756] <= mem_n[2756];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2755] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2755] <= mem_n[2755];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2754] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2754] <= mem_n[2754];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2753] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2753] <= mem_n[2753];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2752] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2752] <= mem_n[2752];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2751] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2751] <= mem_n[2751];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2750] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2750] <= mem_n[2750];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2749] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2749] <= mem_n[2749];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2748] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2748] <= mem_n[2748];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2747] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2747] <= mem_n[2747];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2746] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2746] <= mem_n[2746];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2745] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2745] <= mem_n[2745];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2744] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2744] <= mem_n[2744];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2743] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2743] <= mem_n[2743];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2742] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2742] <= mem_n[2742];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2741] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2741] <= mem_n[2741];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2740] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2740] <= mem_n[2740];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2739] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2739] <= mem_n[2739];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2738] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2738] <= mem_n[2738];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2737] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2737] <= mem_n[2737];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2736] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2736] <= mem_n[2736];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2735] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2735] <= mem_n[2735];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2734] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2734] <= mem_n[2734];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2733] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2733] <= mem_n[2733];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2732] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2732] <= mem_n[2732];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2731] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2731] <= mem_n[2731];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2730] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2730] <= mem_n[2730];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2729] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2729] <= mem_n[2729];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2728] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2728] <= mem_n[2728];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2727] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2727] <= mem_n[2727];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2726] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2726] <= mem_n[2726];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2725] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2725] <= mem_n[2725];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2724] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2724] <= mem_n[2724];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2723] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2723] <= mem_n[2723];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2722] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2722] <= mem_n[2722];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2721] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2721] <= mem_n[2721];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2720] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2720] <= mem_n[2720];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2719] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2719] <= mem_n[2719];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2718] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2718] <= mem_n[2718];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2717] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2717] <= mem_n[2717];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2716] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2716] <= mem_n[2716];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2715] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2715] <= mem_n[2715];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2714] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2714] <= mem_n[2714];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2713] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2713] <= mem_n[2713];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2712] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2712] <= mem_n[2712];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2711] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2711] <= mem_n[2711];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2710] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2710] <= mem_n[2710];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2709] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2709] <= mem_n[2709];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2708] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2708] <= mem_n[2708];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2707] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2707] <= mem_n[2707];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2706] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2706] <= mem_n[2706];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2705] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2705] <= mem_n[2705];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2704] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2704] <= mem_n[2704];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2703] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2703] <= mem_n[2703];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2702] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2702] <= mem_n[2702];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2701] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2701] <= mem_n[2701];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2700] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2700] <= mem_n[2700];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2699] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2699] <= mem_n[2699];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2698] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2698] <= mem_n[2698];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2697] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2697] <= mem_n[2697];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2696] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2696] <= mem_n[2696];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2695] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2695] <= mem_n[2695];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2694] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2694] <= mem_n[2694];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2693] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2693] <= mem_n[2693];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2692] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2692] <= mem_n[2692];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2691] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2691] <= mem_n[2691];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2690] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2690] <= mem_n[2690];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2689] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2689] <= mem_n[2689];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2688] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2688] <= mem_n[2688];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2687] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2687] <= mem_n[2687];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2686] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2686] <= mem_n[2686];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2685] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2685] <= mem_n[2685];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2684] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2684] <= mem_n[2684];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2683] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2683] <= mem_n[2683];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2682] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2682] <= mem_n[2682];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2681] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2681] <= mem_n[2681];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2680] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2680] <= mem_n[2680];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2679] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2679] <= mem_n[2679];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2678] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2678] <= mem_n[2678];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2677] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2677] <= mem_n[2677];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2676] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2676] <= mem_n[2676];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2675] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2675] <= mem_n[2675];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2674] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2674] <= mem_n[2674];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2673] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2673] <= mem_n[2673];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2672] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2672] <= mem_n[2672];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2671] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2671] <= mem_n[2671];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2670] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2670] <= mem_n[2670];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2669] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2669] <= mem_n[2669];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2668] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2668] <= mem_n[2668];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2667] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2667] <= mem_n[2667];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2666] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2666] <= mem_n[2666];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2665] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2665] <= mem_n[2665];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2664] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2664] <= mem_n[2664];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2663] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2663] <= mem_n[2663];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2662] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2662] <= mem_n[2662];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2661] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2661] <= mem_n[2661];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2660] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2660] <= mem_n[2660];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2659] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2659] <= mem_n[2659];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2658] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2658] <= mem_n[2658];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2657] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2657] <= mem_n[2657];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2656] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2656] <= mem_n[2656];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2655] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2655] <= mem_n[2655];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2654] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2654] <= mem_n[2654];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2653] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2653] <= mem_n[2653];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2652] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2652] <= mem_n[2652];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2651] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2651] <= mem_n[2651];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2650] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2650] <= mem_n[2650];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2649] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2649] <= mem_n[2649];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2648] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2648] <= mem_n[2648];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2647] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2647] <= mem_n[2647];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2646] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2646] <= mem_n[2646];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2645] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2645] <= mem_n[2645];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2644] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2644] <= mem_n[2644];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2643] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2643] <= mem_n[2643];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2642] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2642] <= mem_n[2642];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2641] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2641] <= mem_n[2641];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2640] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2640] <= mem_n[2640];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2639] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2639] <= mem_n[2639];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2638] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2638] <= mem_n[2638];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2637] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2637] <= mem_n[2637];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2636] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2636] <= mem_n[2636];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2635] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2635] <= mem_n[2635];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2634] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2634] <= mem_n[2634];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2633] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2633] <= mem_n[2633];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2632] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2632] <= mem_n[2632];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2631] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2631] <= mem_n[2631];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2630] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2630] <= mem_n[2630];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2629] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2629] <= mem_n[2629];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2628] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2628] <= mem_n[2628];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2627] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2627] <= mem_n[2627];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2626] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2626] <= mem_n[2626];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2625] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2625] <= mem_n[2625];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2624] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2624] <= mem_n[2624];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2623] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2623] <= mem_n[2623];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2622] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2622] <= mem_n[2622];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2621] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2621] <= mem_n[2621];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2620] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2620] <= mem_n[2620];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2619] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2619] <= mem_n[2619];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2618] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2618] <= mem_n[2618];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2617] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2617] <= mem_n[2617];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2616] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2616] <= mem_n[2616];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2615] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2615] <= mem_n[2615];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2614] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2614] <= mem_n[2614];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2613] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2613] <= mem_n[2613];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2612] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2612] <= mem_n[2612];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2611] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2611] <= mem_n[2611];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2610] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2610] <= mem_n[2610];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2609] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2609] <= mem_n[2609];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2608] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2608] <= mem_n[2608];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2607] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2607] <= mem_n[2607];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2606] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2606] <= mem_n[2606];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2605] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2605] <= mem_n[2605];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2604] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2604] <= mem_n[2604];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2603] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2603] <= mem_n[2603];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2602] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2602] <= mem_n[2602];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2601] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2601] <= mem_n[2601];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2600] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2600] <= mem_n[2600];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2599] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2599] <= mem_n[2599];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2598] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2598] <= mem_n[2598];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2597] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2597] <= mem_n[2597];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2596] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2596] <= mem_n[2596];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2595] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2595] <= mem_n[2595];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2594] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2594] <= mem_n[2594];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2593] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2593] <= mem_n[2593];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2592] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2592] <= mem_n[2592];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2591] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2591] <= mem_n[2591];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2590] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2590] <= mem_n[2590];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2589] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2589] <= mem_n[2589];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2588] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2588] <= mem_n[2588];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2587] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2587] <= mem_n[2587];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2586] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2586] <= mem_n[2586];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2585] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2585] <= mem_n[2585];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2584] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2584] <= mem_n[2584];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2583] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2583] <= mem_n[2583];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2582] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2582] <= mem_n[2582];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2581] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2581] <= mem_n[2581];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2580] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2580] <= mem_n[2580];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2579] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2579] <= mem_n[2579];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2578] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2578] <= mem_n[2578];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2577] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2577] <= mem_n[2577];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2576] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2576] <= mem_n[2576];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2575] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2575] <= mem_n[2575];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2574] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2574] <= mem_n[2574];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2573] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2573] <= mem_n[2573];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2572] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2572] <= mem_n[2572];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2571] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2571] <= mem_n[2571];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2570] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2570] <= mem_n[2570];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2569] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2569] <= mem_n[2569];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2568] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2568] <= mem_n[2568];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2567] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2567] <= mem_n[2567];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2566] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2566] <= mem_n[2566];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2565] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2565] <= mem_n[2565];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2564] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2564] <= mem_n[2564];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2563] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2563] <= mem_n[2563];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2562] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2562] <= mem_n[2562];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2561] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2561] <= mem_n[2561];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2560] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2560] <= mem_n[2560];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2559] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2559] <= mem_n[2559];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2558] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2558] <= mem_n[2558];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2557] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2557] <= mem_n[2557];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2556] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2556] <= mem_n[2556];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2555] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2555] <= mem_n[2555];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2554] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2554] <= mem_n[2554];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2553] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2553] <= mem_n[2553];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2552] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2552] <= mem_n[2552];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2551] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2551] <= mem_n[2551];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2550] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2550] <= mem_n[2550];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2549] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2549] <= mem_n[2549];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2548] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2548] <= mem_n[2548];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2547] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2547] <= mem_n[2547];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2546] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2546] <= mem_n[2546];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2545] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2545] <= mem_n[2545];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2544] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2544] <= mem_n[2544];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2543] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2543] <= mem_n[2543];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2542] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2542] <= mem_n[2542];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2541] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2541] <= mem_n[2541];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2540] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2540] <= mem_n[2540];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2539] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2539] <= mem_n[2539];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2538] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2538] <= mem_n[2538];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2537] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2537] <= mem_n[2537];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2536] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2536] <= mem_n[2536];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2535] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2535] <= mem_n[2535];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2534] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2534] <= mem_n[2534];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2533] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2533] <= mem_n[2533];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2532] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2532] <= mem_n[2532];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2531] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2531] <= mem_n[2531];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2530] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2530] <= mem_n[2530];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2529] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2529] <= mem_n[2529];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2528] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2528] <= mem_n[2528];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2527] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2527] <= mem_n[2527];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2526] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2526] <= mem_n[2526];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2525] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2525] <= mem_n[2525];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2524] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2524] <= mem_n[2524];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2523] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2523] <= mem_n[2523];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2522] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2522] <= mem_n[2522];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2521] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2521] <= mem_n[2521];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2520] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2520] <= mem_n[2520];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2519] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2519] <= mem_n[2519];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2518] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2518] <= mem_n[2518];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2517] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2517] <= mem_n[2517];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2516] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2516] <= mem_n[2516];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2515] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2515] <= mem_n[2515];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2514] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2514] <= mem_n[2514];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2513] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2513] <= mem_n[2513];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2512] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2512] <= mem_n[2512];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2511] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2511] <= mem_n[2511];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2510] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2510] <= mem_n[2510];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2509] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2509] <= mem_n[2509];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2508] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2508] <= mem_n[2508];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2507] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2507] <= mem_n[2507];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2506] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2506] <= mem_n[2506];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2505] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2505] <= mem_n[2505];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2504] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2504] <= mem_n[2504];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2503] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2503] <= mem_n[2503];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2502] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2502] <= mem_n[2502];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2501] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2501] <= mem_n[2501];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2500] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2500] <= mem_n[2500];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2499] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2499] <= mem_n[2499];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2498] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2498] <= mem_n[2498];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2497] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2497] <= mem_n[2497];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2496] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2496] <= mem_n[2496];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2495] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2495] <= mem_n[2495];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2494] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2494] <= mem_n[2494];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2493] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2493] <= mem_n[2493];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2492] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2492] <= mem_n[2492];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2491] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2491] <= mem_n[2491];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2490] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2490] <= mem_n[2490];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2489] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2489] <= mem_n[2489];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2488] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2488] <= mem_n[2488];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2487] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2487] <= mem_n[2487];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2486] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2486] <= mem_n[2486];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2485] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2485] <= mem_n[2485];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2484] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2484] <= mem_n[2484];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2483] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2483] <= mem_n[2483];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2482] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2482] <= mem_n[2482];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2481] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2481] <= mem_n[2481];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2480] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2480] <= mem_n[2480];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2479] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2479] <= mem_n[2479];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2478] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2478] <= mem_n[2478];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2477] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2477] <= mem_n[2477];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2476] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2476] <= mem_n[2476];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2475] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2475] <= mem_n[2475];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2474] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2474] <= mem_n[2474];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2473] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2473] <= mem_n[2473];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2472] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2472] <= mem_n[2472];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2471] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2471] <= mem_n[2471];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2470] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2470] <= mem_n[2470];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2469] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2469] <= mem_n[2469];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2468] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2468] <= mem_n[2468];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2467] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2467] <= mem_n[2467];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2466] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2466] <= mem_n[2466];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2465] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2465] <= mem_n[2465];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2464] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2464] <= mem_n[2464];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2463] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2463] <= mem_n[2463];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2462] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2462] <= mem_n[2462];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2461] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2461] <= mem_n[2461];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2460] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2460] <= mem_n[2460];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2459] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2459] <= mem_n[2459];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2458] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2458] <= mem_n[2458];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2457] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2457] <= mem_n[2457];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2456] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2456] <= mem_n[2456];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2455] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2455] <= mem_n[2455];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2454] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2454] <= mem_n[2454];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2453] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2453] <= mem_n[2453];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2452] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2452] <= mem_n[2452];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2451] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2451] <= mem_n[2451];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2450] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2450] <= mem_n[2450];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2449] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2449] <= mem_n[2449];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2448] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2448] <= mem_n[2448];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2447] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2447] <= mem_n[2447];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2446] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2446] <= mem_n[2446];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2445] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2445] <= mem_n[2445];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2444] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2444] <= mem_n[2444];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2443] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2443] <= mem_n[2443];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2442] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2442] <= mem_n[2442];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2441] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2441] <= mem_n[2441];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2440] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2440] <= mem_n[2440];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2439] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2439] <= mem_n[2439];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2438] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2438] <= mem_n[2438];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2437] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2437] <= mem_n[2437];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2436] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2436] <= mem_n[2436];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2435] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2435] <= mem_n[2435];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2434] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2434] <= mem_n[2434];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2433] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2433] <= mem_n[2433];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2432] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2432] <= mem_n[2432];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2431] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2431] <= mem_n[2431];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2430] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2430] <= mem_n[2430];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2429] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2429] <= mem_n[2429];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2428] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2428] <= mem_n[2428];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2427] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2427] <= mem_n[2427];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2426] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2426] <= mem_n[2426];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2425] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2425] <= mem_n[2425];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2424] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2424] <= mem_n[2424];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2423] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2423] <= mem_n[2423];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2422] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2422] <= mem_n[2422];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2421] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2421] <= mem_n[2421];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2420] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2420] <= mem_n[2420];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2419] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2419] <= mem_n[2419];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2418] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2418] <= mem_n[2418];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2417] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2417] <= mem_n[2417];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2416] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2416] <= mem_n[2416];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2415] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2415] <= mem_n[2415];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2414] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2414] <= mem_n[2414];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2413] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2413] <= mem_n[2413];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2412] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2412] <= mem_n[2412];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2411] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2411] <= mem_n[2411];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2410] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2410] <= mem_n[2410];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2409] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2409] <= mem_n[2409];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2408] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2408] <= mem_n[2408];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2407] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2407] <= mem_n[2407];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2406] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2406] <= mem_n[2406];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2405] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2405] <= mem_n[2405];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2404] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2404] <= mem_n[2404];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2403] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2403] <= mem_n[2403];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2402] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2402] <= mem_n[2402];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2401] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2401] <= mem_n[2401];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2400] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2400] <= mem_n[2400];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2399] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2399] <= mem_n[2399];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2398] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2398] <= mem_n[2398];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2397] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2397] <= mem_n[2397];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2396] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2396] <= mem_n[2396];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2395] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2395] <= mem_n[2395];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2394] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2394] <= mem_n[2394];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2393] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2393] <= mem_n[2393];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2392] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2392] <= mem_n[2392];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2391] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2391] <= mem_n[2391];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2390] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2390] <= mem_n[2390];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2389] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2389] <= mem_n[2389];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2388] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2388] <= mem_n[2388];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2387] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2387] <= mem_n[2387];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2386] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2386] <= mem_n[2386];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2385] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2385] <= mem_n[2385];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2384] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2384] <= mem_n[2384];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2383] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2383] <= mem_n[2383];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2382] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2382] <= mem_n[2382];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2381] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2381] <= mem_n[2381];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2380] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2380] <= mem_n[2380];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2379] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2379] <= mem_n[2379];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2378] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2378] <= mem_n[2378];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2377] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2377] <= mem_n[2377];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2376] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2376] <= mem_n[2376];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2375] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2375] <= mem_n[2375];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2374] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2374] <= mem_n[2374];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2373] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2373] <= mem_n[2373];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2372] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2372] <= mem_n[2372];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2371] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2371] <= mem_n[2371];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2370] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2370] <= mem_n[2370];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2369] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2369] <= mem_n[2369];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2368] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2368] <= mem_n[2368];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2367] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2367] <= mem_n[2367];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2366] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2366] <= mem_n[2366];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2365] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2365] <= mem_n[2365];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2364] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2364] <= mem_n[2364];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2363] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2363] <= mem_n[2363];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2362] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2362] <= mem_n[2362];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2361] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2361] <= mem_n[2361];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2360] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2360] <= mem_n[2360];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2359] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2359] <= mem_n[2359];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2358] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2358] <= mem_n[2358];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2357] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2357] <= mem_n[2357];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2356] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2356] <= mem_n[2356];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2355] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2355] <= mem_n[2355];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2354] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2354] <= mem_n[2354];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2353] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2353] <= mem_n[2353];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2352] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2352] <= mem_n[2352];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2351] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2351] <= mem_n[2351];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2350] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2350] <= mem_n[2350];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2349] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2349] <= mem_n[2349];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2348] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2348] <= mem_n[2348];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2347] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2347] <= mem_n[2347];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2346] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2346] <= mem_n[2346];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2345] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2345] <= mem_n[2345];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2344] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2344] <= mem_n[2344];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2343] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2343] <= mem_n[2343];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2342] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2342] <= mem_n[2342];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2341] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2341] <= mem_n[2341];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2340] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2340] <= mem_n[2340];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2339] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2339] <= mem_n[2339];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2338] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2338] <= mem_n[2338];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2337] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2337] <= mem_n[2337];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2336] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2336] <= mem_n[2336];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2335] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2335] <= mem_n[2335];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2334] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2334] <= mem_n[2334];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2333] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2333] <= mem_n[2333];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2332] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2332] <= mem_n[2332];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2331] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2331] <= mem_n[2331];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2330] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2330] <= mem_n[2330];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2329] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2329] <= mem_n[2329];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2328] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2328] <= mem_n[2328];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2327] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2327] <= mem_n[2327];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2326] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2326] <= mem_n[2326];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2325] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2325] <= mem_n[2325];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2324] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2324] <= mem_n[2324];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2323] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2323] <= mem_n[2323];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2322] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2322] <= mem_n[2322];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2321] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2321] <= mem_n[2321];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2320] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2320] <= mem_n[2320];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2319] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2319] <= mem_n[2319];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2318] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2318] <= mem_n[2318];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2317] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2317] <= mem_n[2317];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2316] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2316] <= mem_n[2316];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2315] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2315] <= mem_n[2315];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2314] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2314] <= mem_n[2314];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2313] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2313] <= mem_n[2313];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2312] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2312] <= mem_n[2312];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2311] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2311] <= mem_n[2311];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2310] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2310] <= mem_n[2310];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2309] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2309] <= mem_n[2309];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2308] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2308] <= mem_n[2308];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2307] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2307] <= mem_n[2307];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2306] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2306] <= mem_n[2306];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2305] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2305] <= mem_n[2305];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2304] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2304] <= mem_n[2304];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2303] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2303] <= mem_n[2303];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2302] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2302] <= mem_n[2302];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2301] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2301] <= mem_n[2301];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2300] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2300] <= mem_n[2300];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2299] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2299] <= mem_n[2299];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2298] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2298] <= mem_n[2298];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2297] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2297] <= mem_n[2297];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2296] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2296] <= mem_n[2296];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2295] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2295] <= mem_n[2295];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2294] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2294] <= mem_n[2294];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2293] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2293] <= mem_n[2293];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2292] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2292] <= mem_n[2292];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2291] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2291] <= mem_n[2291];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2290] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2290] <= mem_n[2290];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2289] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2289] <= mem_n[2289];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2288] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2288] <= mem_n[2288];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2287] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2287] <= mem_n[2287];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2286] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2286] <= mem_n[2286];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2285] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2285] <= mem_n[2285];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2284] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2284] <= mem_n[2284];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2283] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2283] <= mem_n[2283];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2282] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2282] <= mem_n[2282];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2281] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2281] <= mem_n[2281];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2280] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2280] <= mem_n[2280];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2279] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2279] <= mem_n[2279];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2278] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2278] <= mem_n[2278];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2277] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2277] <= mem_n[2277];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2276] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2276] <= mem_n[2276];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2275] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2275] <= mem_n[2275];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2274] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2274] <= mem_n[2274];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2273] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2273] <= mem_n[2273];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2272] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2272] <= mem_n[2272];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2271] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2271] <= mem_n[2271];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2270] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2270] <= mem_n[2270];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2269] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2269] <= mem_n[2269];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2268] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2268] <= mem_n[2268];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2267] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2267] <= mem_n[2267];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2266] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2266] <= mem_n[2266];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2265] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2265] <= mem_n[2265];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2264] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2264] <= mem_n[2264];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2263] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2263] <= mem_n[2263];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2262] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2262] <= mem_n[2262];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2261] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2261] <= mem_n[2261];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2260] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2260] <= mem_n[2260];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2259] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2259] <= mem_n[2259];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2258] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2258] <= mem_n[2258];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2257] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2257] <= mem_n[2257];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2256] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2256] <= mem_n[2256];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2255] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2255] <= mem_n[2255];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2254] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2254] <= mem_n[2254];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2253] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2253] <= mem_n[2253];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2252] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2252] <= mem_n[2252];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2251] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2251] <= mem_n[2251];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2250] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2250] <= mem_n[2250];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2249] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2249] <= mem_n[2249];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2248] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2248] <= mem_n[2248];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2247] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2247] <= mem_n[2247];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2246] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2246] <= mem_n[2246];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2245] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2245] <= mem_n[2245];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2244] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2244] <= mem_n[2244];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2243] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2243] <= mem_n[2243];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2242] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2242] <= mem_n[2242];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2241] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2241] <= mem_n[2241];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2240] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2240] <= mem_n[2240];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2239] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2239] <= mem_n[2239];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2238] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2238] <= mem_n[2238];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2237] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2237] <= mem_n[2237];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2236] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2236] <= mem_n[2236];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2235] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2235] <= mem_n[2235];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2234] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2234] <= mem_n[2234];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2233] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2233] <= mem_n[2233];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2232] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2232] <= mem_n[2232];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2231] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2231] <= mem_n[2231];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2230] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2230] <= mem_n[2230];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2229] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2229] <= mem_n[2229];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2228] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2228] <= mem_n[2228];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2227] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2227] <= mem_n[2227];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2226] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2226] <= mem_n[2226];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2225] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2225] <= mem_n[2225];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2224] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2224] <= mem_n[2224];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2223] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2223] <= mem_n[2223];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2222] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2222] <= mem_n[2222];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2221] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2221] <= mem_n[2221];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2220] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2220] <= mem_n[2220];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2219] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2219] <= mem_n[2219];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2218] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2218] <= mem_n[2218];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2217] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2217] <= mem_n[2217];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2216] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2216] <= mem_n[2216];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2215] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2215] <= mem_n[2215];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2214] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2214] <= mem_n[2214];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2213] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2213] <= mem_n[2213];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2212] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2212] <= mem_n[2212];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2211] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2211] <= mem_n[2211];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2210] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2210] <= mem_n[2210];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2209] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2209] <= mem_n[2209];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2208] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2208] <= mem_n[2208];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2207] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2207] <= mem_n[2207];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2206] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2206] <= mem_n[2206];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2205] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2205] <= mem_n[2205];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2204] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2204] <= mem_n[2204];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2203] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2203] <= mem_n[2203];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2202] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2202] <= mem_n[2202];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2201] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2201] <= mem_n[2201];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2200] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2200] <= mem_n[2200];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2199] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2199] <= mem_n[2199];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2198] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2198] <= mem_n[2198];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2197] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2197] <= mem_n[2197];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2196] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2196] <= mem_n[2196];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2195] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2195] <= mem_n[2195];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2194] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2194] <= mem_n[2194];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2193] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2193] <= mem_n[2193];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2192] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2192] <= mem_n[2192];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2191] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2191] <= mem_n[2191];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2190] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2190] <= mem_n[2190];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2189] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2189] <= mem_n[2189];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2188] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2188] <= mem_n[2188];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2187] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2187] <= mem_n[2187];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2186] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2186] <= mem_n[2186];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2185] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2185] <= mem_n[2185];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2184] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2184] <= mem_n[2184];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2183] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2183] <= mem_n[2183];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2182] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2182] <= mem_n[2182];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2181] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2181] <= mem_n[2181];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2180] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2180] <= mem_n[2180];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2179] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2179] <= mem_n[2179];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2178] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2178] <= mem_n[2178];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2177] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2177] <= mem_n[2177];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2176] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2176] <= mem_n[2176];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2175] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2175] <= mem_n[2175];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2174] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2174] <= mem_n[2174];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2173] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2173] <= mem_n[2173];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2172] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2172] <= mem_n[2172];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2171] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2171] <= mem_n[2171];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2170] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2170] <= mem_n[2170];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2169] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2169] <= mem_n[2169];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2168] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2168] <= mem_n[2168];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2167] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2167] <= mem_n[2167];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2166] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2166] <= mem_n[2166];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2165] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2165] <= mem_n[2165];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2164] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2164] <= mem_n[2164];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2163] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2163] <= mem_n[2163];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2162] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2162] <= mem_n[2162];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2161] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2161] <= mem_n[2161];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2160] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2160] <= mem_n[2160];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2159] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2159] <= mem_n[2159];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2158] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2158] <= mem_n[2158];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2157] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2157] <= mem_n[2157];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2156] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2156] <= mem_n[2156];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2155] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2155] <= mem_n[2155];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2154] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2154] <= mem_n[2154];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2153] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2153] <= mem_n[2153];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2152] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2152] <= mem_n[2152];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2151] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2151] <= mem_n[2151];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2150] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2150] <= mem_n[2150];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2149] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2149] <= mem_n[2149];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2148] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2148] <= mem_n[2148];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2147] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2147] <= mem_n[2147];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2146] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2146] <= mem_n[2146];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2145] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2145] <= mem_n[2145];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2144] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2144] <= mem_n[2144];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2143] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2143] <= mem_n[2143];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2142] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2142] <= mem_n[2142];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2141] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2141] <= mem_n[2141];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2140] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2140] <= mem_n[2140];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2139] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2139] <= mem_n[2139];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2138] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2138] <= mem_n[2138];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2137] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2137] <= mem_n[2137];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2136] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2136] <= mem_n[2136];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2135] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2135] <= mem_n[2135];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2134] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2134] <= mem_n[2134];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2133] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2133] <= mem_n[2133];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2132] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2132] <= mem_n[2132];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2131] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2131] <= mem_n[2131];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2130] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2130] <= mem_n[2130];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2129] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2129] <= mem_n[2129];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2128] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2128] <= mem_n[2128];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2127] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2127] <= mem_n[2127];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2126] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2126] <= mem_n[2126];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2125] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2125] <= mem_n[2125];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2124] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2124] <= mem_n[2124];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2123] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2123] <= mem_n[2123];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2122] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2122] <= mem_n[2122];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2121] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2121] <= mem_n[2121];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2120] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2120] <= mem_n[2120];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2119] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2119] <= mem_n[2119];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2118] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2118] <= mem_n[2118];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2117] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2117] <= mem_n[2117];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2116] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2116] <= mem_n[2116];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2115] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2115] <= mem_n[2115];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2114] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2114] <= mem_n[2114];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2113] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2113] <= mem_n[2113];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2112] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2112] <= mem_n[2112];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2111] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2111] <= mem_n[2111];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2110] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2110] <= mem_n[2110];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2109] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2109] <= mem_n[2109];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2108] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2108] <= mem_n[2108];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2107] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2107] <= mem_n[2107];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2106] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2106] <= mem_n[2106];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2105] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2105] <= mem_n[2105];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2104] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2104] <= mem_n[2104];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2103] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2103] <= mem_n[2103];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2102] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2102] <= mem_n[2102];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2101] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2101] <= mem_n[2101];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2100] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2100] <= mem_n[2100];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2099] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2099] <= mem_n[2099];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2098] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2098] <= mem_n[2098];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2097] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2097] <= mem_n[2097];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2096] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2096] <= mem_n[2096];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2095] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2095] <= mem_n[2095];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2094] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2094] <= mem_n[2094];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2093] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2093] <= mem_n[2093];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2092] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2092] <= mem_n[2092];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2091] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2091] <= mem_n[2091];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2090] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2090] <= mem_n[2090];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2089] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2089] <= mem_n[2089];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2088] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2088] <= mem_n[2088];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2087] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2087] <= mem_n[2087];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2086] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2086] <= mem_n[2086];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2085] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2085] <= mem_n[2085];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2084] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2084] <= mem_n[2084];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2083] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2083] <= mem_n[2083];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2082] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2082] <= mem_n[2082];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2081] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2081] <= mem_n[2081];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2080] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2080] <= mem_n[2080];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2079] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2079] <= mem_n[2079];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2078] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2078] <= mem_n[2078];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2077] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2077] <= mem_n[2077];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2076] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2076] <= mem_n[2076];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2075] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2075] <= mem_n[2075];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2074] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2074] <= mem_n[2074];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2073] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2073] <= mem_n[2073];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2072] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2072] <= mem_n[2072];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2071] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2071] <= mem_n[2071];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2070] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2070] <= mem_n[2070];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2069] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2069] <= mem_n[2069];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2068] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2068] <= mem_n[2068];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2067] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2067] <= mem_n[2067];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2066] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2066] <= mem_n[2066];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2065] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2065] <= mem_n[2065];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2064] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2064] <= mem_n[2064];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2063] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2063] <= mem_n[2063];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2062] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2062] <= mem_n[2062];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2061] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2061] <= mem_n[2061];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2060] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2060] <= mem_n[2060];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2059] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2059] <= mem_n[2059];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2058] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2058] <= mem_n[2058];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2057] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2057] <= mem_n[2057];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2056] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2056] <= mem_n[2056];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2055] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2055] <= mem_n[2055];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2054] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2054] <= mem_n[2054];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2053] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2053] <= mem_n[2053];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2052] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2052] <= mem_n[2052];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2051] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2051] <= mem_n[2051];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2050] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2050] <= mem_n[2050];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2049] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2049] <= mem_n[2049];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2048] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2048] <= mem_n[2048];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2047] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2047] <= mem_n[2047];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2046] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2046] <= mem_n[2046];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2045] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2045] <= mem_n[2045];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2044] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2044] <= mem_n[2044];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2043] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2043] <= mem_n[2043];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2042] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2042] <= mem_n[2042];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2041] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2041] <= mem_n[2041];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2040] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2040] <= mem_n[2040];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2039] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2039] <= mem_n[2039];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2038] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2038] <= mem_n[2038];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2037] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2037] <= mem_n[2037];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2036] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2036] <= mem_n[2036];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2035] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2035] <= mem_n[2035];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2034] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2034] <= mem_n[2034];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2033] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2033] <= mem_n[2033];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2032] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2032] <= mem_n[2032];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2031] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2031] <= mem_n[2031];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2030] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2030] <= mem_n[2030];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2029] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2029] <= mem_n[2029];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2028] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2028] <= mem_n[2028];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2027] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2027] <= mem_n[2027];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2026] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2026] <= mem_n[2026];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2025] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2025] <= mem_n[2025];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2024] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2024] <= mem_n[2024];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2023] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2023] <= mem_n[2023];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2022] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2022] <= mem_n[2022];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2021] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2021] <= mem_n[2021];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2020] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2020] <= mem_n[2020];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2019] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2019] <= mem_n[2019];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2018] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2018] <= mem_n[2018];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2017] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2017] <= mem_n[2017];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2016] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2016] <= mem_n[2016];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2015] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2015] <= mem_n[2015];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2014] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2014] <= mem_n[2014];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2013] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2013] <= mem_n[2013];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2012] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2012] <= mem_n[2012];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2011] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2011] <= mem_n[2011];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2010] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2010] <= mem_n[2010];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2009] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2009] <= mem_n[2009];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2008] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2008] <= mem_n[2008];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2007] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2007] <= mem_n[2007];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2006] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2006] <= mem_n[2006];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2005] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2005] <= mem_n[2005];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2004] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2004] <= mem_n[2004];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2003] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2003] <= mem_n[2003];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2002] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2002] <= mem_n[2002];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2001] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2001] <= mem_n[2001];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2000] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2000] <= mem_n[2000];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1999] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1999] <= mem_n[1999];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1998] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1998] <= mem_n[1998];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1997] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1997] <= mem_n[1997];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1996] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1996] <= mem_n[1996];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1995] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1995] <= mem_n[1995];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1994] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1994] <= mem_n[1994];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1993] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1993] <= mem_n[1993];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1992] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1992] <= mem_n[1992];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1991] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1991] <= mem_n[1991];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1990] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1990] <= mem_n[1990];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1989] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1989] <= mem_n[1989];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1988] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1988] <= mem_n[1988];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1987] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1987] <= mem_n[1987];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1986] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1986] <= mem_n[1986];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1985] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1985] <= mem_n[1985];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1984] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1984] <= mem_n[1984];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1983] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1983] <= mem_n[1983];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1982] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1982] <= mem_n[1982];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1981] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1981] <= mem_n[1981];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1980] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1980] <= mem_n[1980];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1979] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1979] <= mem_n[1979];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1978] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1978] <= mem_n[1978];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1977] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1977] <= mem_n[1977];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1976] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1976] <= mem_n[1976];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1975] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1975] <= mem_n[1975];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1974] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1974] <= mem_n[1974];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1973] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1973] <= mem_n[1973];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1972] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1972] <= mem_n[1972];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1971] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1971] <= mem_n[1971];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1970] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1970] <= mem_n[1970];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1969] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1969] <= mem_n[1969];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1968] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1968] <= mem_n[1968];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1967] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1967] <= mem_n[1967];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1966] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1966] <= mem_n[1966];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1965] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1965] <= mem_n[1965];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1964] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1964] <= mem_n[1964];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1963] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1963] <= mem_n[1963];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1962] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1962] <= mem_n[1962];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1961] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1961] <= mem_n[1961];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1960] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1960] <= mem_n[1960];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1959] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1959] <= mem_n[1959];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1958] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1958] <= mem_n[1958];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1957] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1957] <= mem_n[1957];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1956] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1956] <= mem_n[1956];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1955] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1955] <= mem_n[1955];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1954] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1954] <= mem_n[1954];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1953] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1953] <= mem_n[1953];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1952] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1952] <= mem_n[1952];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1951] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1951] <= mem_n[1951];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1950] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1950] <= mem_n[1950];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1949] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1949] <= mem_n[1949];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1948] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1948] <= mem_n[1948];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1947] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1947] <= mem_n[1947];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1946] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1946] <= mem_n[1946];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1945] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1945] <= mem_n[1945];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1944] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1944] <= mem_n[1944];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1943] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1943] <= mem_n[1943];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1942] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1942] <= mem_n[1942];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1941] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1941] <= mem_n[1941];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1940] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1940] <= mem_n[1940];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1939] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1939] <= mem_n[1939];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1938] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1938] <= mem_n[1938];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1937] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1937] <= mem_n[1937];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1936] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1936] <= mem_n[1936];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1935] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1935] <= mem_n[1935];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1934] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1934] <= mem_n[1934];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1933] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1933] <= mem_n[1933];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1932] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1932] <= mem_n[1932];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1931] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1931] <= mem_n[1931];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1930] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1930] <= mem_n[1930];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1929] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1929] <= mem_n[1929];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1928] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1928] <= mem_n[1928];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1927] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1927] <= mem_n[1927];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1926] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1926] <= mem_n[1926];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1925] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1925] <= mem_n[1925];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1924] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1924] <= mem_n[1924];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1923] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1923] <= mem_n[1923];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1922] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1922] <= mem_n[1922];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1921] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1921] <= mem_n[1921];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1920] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1920] <= mem_n[1920];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1919] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1919] <= mem_n[1919];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1918] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1918] <= mem_n[1918];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1917] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1917] <= mem_n[1917];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1916] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1916] <= mem_n[1916];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1915] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1915] <= mem_n[1915];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1914] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1914] <= mem_n[1914];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1913] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1913] <= mem_n[1913];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1912] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1912] <= mem_n[1912];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1911] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1911] <= mem_n[1911];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1910] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1910] <= mem_n[1910];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1909] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1909] <= mem_n[1909];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1908] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1908] <= mem_n[1908];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1907] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1907] <= mem_n[1907];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1906] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1906] <= mem_n[1906];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1905] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1905] <= mem_n[1905];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1904] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1904] <= mem_n[1904];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1903] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1903] <= mem_n[1903];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1902] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1902] <= mem_n[1902];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1901] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1901] <= mem_n[1901];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1900] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1900] <= mem_n[1900];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1899] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1899] <= mem_n[1899];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1898] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1898] <= mem_n[1898];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1897] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1897] <= mem_n[1897];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1896] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1896] <= mem_n[1896];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1895] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1895] <= mem_n[1895];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1894] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1894] <= mem_n[1894];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1893] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1893] <= mem_n[1893];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1892] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1892] <= mem_n[1892];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1891] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1891] <= mem_n[1891];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1890] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1890] <= mem_n[1890];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1889] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1889] <= mem_n[1889];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1888] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1888] <= mem_n[1888];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1887] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1887] <= mem_n[1887];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1886] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1886] <= mem_n[1886];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1885] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1885] <= mem_n[1885];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1884] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1884] <= mem_n[1884];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1883] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1883] <= mem_n[1883];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1882] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1882] <= mem_n[1882];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1881] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1881] <= mem_n[1881];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1880] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1880] <= mem_n[1880];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1879] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1879] <= mem_n[1879];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1878] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1878] <= mem_n[1878];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1877] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1877] <= mem_n[1877];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1876] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1876] <= mem_n[1876];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1875] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1875] <= mem_n[1875];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1874] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1874] <= mem_n[1874];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1873] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1873] <= mem_n[1873];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1872] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1872] <= mem_n[1872];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1871] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1871] <= mem_n[1871];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1870] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1870] <= mem_n[1870];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1869] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1869] <= mem_n[1869];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1868] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1868] <= mem_n[1868];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1867] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1867] <= mem_n[1867];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1866] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1866] <= mem_n[1866];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1865] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1865] <= mem_n[1865];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1864] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1864] <= mem_n[1864];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1863] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1863] <= mem_n[1863];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1862] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1862] <= mem_n[1862];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1861] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1861] <= mem_n[1861];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1860] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1860] <= mem_n[1860];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1859] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1859] <= mem_n[1859];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1858] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1858] <= mem_n[1858];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1857] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1857] <= mem_n[1857];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1856] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1856] <= mem_n[1856];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1855] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1855] <= mem_n[1855];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1854] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1854] <= mem_n[1854];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1853] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1853] <= mem_n[1853];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1852] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1852] <= mem_n[1852];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1851] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1851] <= mem_n[1851];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1850] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1850] <= mem_n[1850];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1849] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1849] <= mem_n[1849];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1848] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1848] <= mem_n[1848];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1847] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1847] <= mem_n[1847];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1846] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1846] <= mem_n[1846];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1845] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1845] <= mem_n[1845];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1844] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1844] <= mem_n[1844];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1843] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1843] <= mem_n[1843];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1842] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1842] <= mem_n[1842];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1841] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1841] <= mem_n[1841];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1840] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1840] <= mem_n[1840];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1839] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1839] <= mem_n[1839];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1838] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1838] <= mem_n[1838];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1837] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1837] <= mem_n[1837];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1836] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1836] <= mem_n[1836];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1835] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1835] <= mem_n[1835];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1834] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1834] <= mem_n[1834];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1833] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1833] <= mem_n[1833];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1832] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1832] <= mem_n[1832];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1831] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1831] <= mem_n[1831];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1830] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1830] <= mem_n[1830];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1829] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1829] <= mem_n[1829];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1828] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1828] <= mem_n[1828];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1827] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1827] <= mem_n[1827];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1826] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1826] <= mem_n[1826];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1825] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1825] <= mem_n[1825];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1824] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1824] <= mem_n[1824];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1823] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1823] <= mem_n[1823];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1822] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1822] <= mem_n[1822];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1821] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1821] <= mem_n[1821];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1820] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1820] <= mem_n[1820];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1819] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1819] <= mem_n[1819];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1818] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1818] <= mem_n[1818];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1817] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1817] <= mem_n[1817];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1816] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1816] <= mem_n[1816];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1815] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1815] <= mem_n[1815];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1814] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1814] <= mem_n[1814];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1813] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1813] <= mem_n[1813];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1812] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1812] <= mem_n[1812];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1811] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1811] <= mem_n[1811];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1810] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1810] <= mem_n[1810];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1809] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1809] <= mem_n[1809];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1808] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1808] <= mem_n[1808];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1807] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1807] <= mem_n[1807];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1806] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1806] <= mem_n[1806];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1805] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1805] <= mem_n[1805];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1804] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1804] <= mem_n[1804];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1803] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1803] <= mem_n[1803];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1802] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1802] <= mem_n[1802];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1801] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1801] <= mem_n[1801];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1800] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1800] <= mem_n[1800];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1799] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1799] <= mem_n[1799];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1798] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1798] <= mem_n[1798];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1797] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1797] <= mem_n[1797];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1796] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1796] <= mem_n[1796];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1795] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1795] <= mem_n[1795];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1794] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1794] <= mem_n[1794];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1793] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1793] <= mem_n[1793];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1792] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1792] <= mem_n[1792];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1791] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1791] <= mem_n[1791];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1790] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1790] <= mem_n[1790];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1789] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1789] <= mem_n[1789];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1788] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1788] <= mem_n[1788];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1787] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1787] <= mem_n[1787];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1786] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1786] <= mem_n[1786];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1785] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1785] <= mem_n[1785];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1784] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1784] <= mem_n[1784];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1783] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1783] <= mem_n[1783];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1782] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1782] <= mem_n[1782];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1781] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1781] <= mem_n[1781];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1780] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1780] <= mem_n[1780];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1779] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1779] <= mem_n[1779];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1778] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1778] <= mem_n[1778];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1777] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1777] <= mem_n[1777];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1776] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1776] <= mem_n[1776];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1775] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1775] <= mem_n[1775];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1774] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1774] <= mem_n[1774];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1773] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1773] <= mem_n[1773];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1772] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1772] <= mem_n[1772];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1771] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1771] <= mem_n[1771];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1770] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1770] <= mem_n[1770];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1769] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1769] <= mem_n[1769];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1768] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1768] <= mem_n[1768];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1767] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1767] <= mem_n[1767];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1766] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1766] <= mem_n[1766];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1765] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1765] <= mem_n[1765];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1764] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1764] <= mem_n[1764];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1763] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1763] <= mem_n[1763];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1762] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1762] <= mem_n[1762];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1761] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1761] <= mem_n[1761];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1760] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1760] <= mem_n[1760];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1759] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1759] <= mem_n[1759];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1758] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1758] <= mem_n[1758];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1757] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1757] <= mem_n[1757];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1756] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1756] <= mem_n[1756];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1755] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1755] <= mem_n[1755];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1754] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1754] <= mem_n[1754];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1753] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1753] <= mem_n[1753];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1752] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1752] <= mem_n[1752];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1751] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1751] <= mem_n[1751];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1750] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1750] <= mem_n[1750];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1749] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1749] <= mem_n[1749];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1748] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1748] <= mem_n[1748];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1747] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1747] <= mem_n[1747];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1746] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1746] <= mem_n[1746];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1745] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1745] <= mem_n[1745];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1744] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1744] <= mem_n[1744];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1743] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1743] <= mem_n[1743];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1742] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1742] <= mem_n[1742];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1741] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1741] <= mem_n[1741];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1740] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1740] <= mem_n[1740];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1739] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1739] <= mem_n[1739];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1738] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1738] <= mem_n[1738];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1737] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1737] <= mem_n[1737];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1736] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1736] <= mem_n[1736];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1735] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1735] <= mem_n[1735];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1734] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1734] <= mem_n[1734];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1733] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1733] <= mem_n[1733];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1732] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1732] <= mem_n[1732];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1731] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1731] <= mem_n[1731];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1730] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1730] <= mem_n[1730];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1729] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1729] <= mem_n[1729];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1728] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1728] <= mem_n[1728];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1727] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1727] <= mem_n[1727];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1726] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1726] <= mem_n[1726];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1725] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1725] <= mem_n[1725];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1724] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1724] <= mem_n[1724];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1723] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1723] <= mem_n[1723];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1722] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1722] <= mem_n[1722];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1721] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1721] <= mem_n[1721];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1720] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1720] <= mem_n[1720];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1719] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1719] <= mem_n[1719];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1718] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1718] <= mem_n[1718];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1717] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1717] <= mem_n[1717];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1716] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1716] <= mem_n[1716];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1715] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1715] <= mem_n[1715];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1714] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1714] <= mem_n[1714];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1713] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1713] <= mem_n[1713];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1712] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1712] <= mem_n[1712];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1711] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1711] <= mem_n[1711];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1710] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1710] <= mem_n[1710];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1709] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1709] <= mem_n[1709];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1708] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1708] <= mem_n[1708];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1707] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1707] <= mem_n[1707];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1706] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1706] <= mem_n[1706];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1705] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1705] <= mem_n[1705];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1704] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1704] <= mem_n[1704];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1703] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1703] <= mem_n[1703];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1702] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1702] <= mem_n[1702];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1701] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1701] <= mem_n[1701];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1700] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1700] <= mem_n[1700];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1699] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1699] <= mem_n[1699];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1698] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1698] <= mem_n[1698];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1697] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1697] <= mem_n[1697];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1696] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1696] <= mem_n[1696];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1695] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1695] <= mem_n[1695];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1694] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1694] <= mem_n[1694];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1693] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1693] <= mem_n[1693];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1692] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1692] <= mem_n[1692];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1691] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1691] <= mem_n[1691];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1690] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1690] <= mem_n[1690];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1689] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1689] <= mem_n[1689];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1688] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1688] <= mem_n[1688];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1687] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1687] <= mem_n[1687];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1686] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1686] <= mem_n[1686];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1685] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1685] <= mem_n[1685];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1684] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1684] <= mem_n[1684];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1683] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1683] <= mem_n[1683];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1682] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1682] <= mem_n[1682];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1681] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1681] <= mem_n[1681];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1680] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1680] <= mem_n[1680];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1679] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1679] <= mem_n[1679];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1678] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1678] <= mem_n[1678];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1677] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1677] <= mem_n[1677];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1676] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1676] <= mem_n[1676];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1675] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1675] <= mem_n[1675];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1674] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1674] <= mem_n[1674];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1673] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1673] <= mem_n[1673];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1672] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1672] <= mem_n[1672];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1671] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1671] <= mem_n[1671];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1670] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1670] <= mem_n[1670];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1669] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1669] <= mem_n[1669];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1668] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1668] <= mem_n[1668];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1667] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1667] <= mem_n[1667];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1666] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1666] <= mem_n[1666];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1665] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1665] <= mem_n[1665];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1664] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1664] <= mem_n[1664];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1663] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1663] <= mem_n[1663];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1662] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1662] <= mem_n[1662];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1661] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1661] <= mem_n[1661];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1660] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1660] <= mem_n[1660];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1659] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1659] <= mem_n[1659];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1658] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1658] <= mem_n[1658];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1657] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1657] <= mem_n[1657];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1656] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1656] <= mem_n[1656];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1655] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1655] <= mem_n[1655];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1654] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1654] <= mem_n[1654];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1653] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1653] <= mem_n[1653];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1652] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1652] <= mem_n[1652];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1651] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1651] <= mem_n[1651];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1650] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1650] <= mem_n[1650];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1649] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1649] <= mem_n[1649];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1648] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1648] <= mem_n[1648];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1647] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1647] <= mem_n[1647];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1646] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1646] <= mem_n[1646];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1645] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1645] <= mem_n[1645];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1644] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1644] <= mem_n[1644];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1643] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1643] <= mem_n[1643];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1642] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1642] <= mem_n[1642];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1641] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1641] <= mem_n[1641];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1640] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1640] <= mem_n[1640];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1639] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1639] <= mem_n[1639];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1638] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1638] <= mem_n[1638];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1637] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1637] <= mem_n[1637];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1636] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1636] <= mem_n[1636];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1635] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1635] <= mem_n[1635];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1634] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1634] <= mem_n[1634];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1633] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1633] <= mem_n[1633];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1632] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1632] <= mem_n[1632];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1631] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1631] <= mem_n[1631];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1630] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1630] <= mem_n[1630];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1629] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1629] <= mem_n[1629];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1628] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1628] <= mem_n[1628];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1627] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1627] <= mem_n[1627];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1626] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1626] <= mem_n[1626];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1625] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1625] <= mem_n[1625];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1624] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1624] <= mem_n[1624];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1623] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1623] <= mem_n[1623];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1622] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1622] <= mem_n[1622];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1621] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1621] <= mem_n[1621];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1620] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1620] <= mem_n[1620];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1619] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1619] <= mem_n[1619];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1618] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1618] <= mem_n[1618];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1617] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1617] <= mem_n[1617];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1616] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1616] <= mem_n[1616];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1615] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1615] <= mem_n[1615];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1614] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1614] <= mem_n[1614];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1613] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1613] <= mem_n[1613];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1612] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1612] <= mem_n[1612];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1611] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1611] <= mem_n[1611];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1610] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1610] <= mem_n[1610];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1609] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1609] <= mem_n[1609];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1608] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1608] <= mem_n[1608];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1607] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1607] <= mem_n[1607];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1606] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1606] <= mem_n[1606];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1605] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1605] <= mem_n[1605];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1604] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1604] <= mem_n[1604];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1603] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1603] <= mem_n[1603];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1602] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1602] <= mem_n[1602];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1601] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1601] <= mem_n[1601];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1600] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1600] <= mem_n[1600];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1599] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1599] <= mem_n[1599];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1598] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1598] <= mem_n[1598];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1597] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1597] <= mem_n[1597];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1596] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1596] <= mem_n[1596];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1595] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1595] <= mem_n[1595];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1594] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1594] <= mem_n[1594];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1593] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1593] <= mem_n[1593];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1592] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1592] <= mem_n[1592];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1591] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1591] <= mem_n[1591];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1590] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1590] <= mem_n[1590];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1589] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1589] <= mem_n[1589];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1588] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1588] <= mem_n[1588];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1587] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1587] <= mem_n[1587];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1586] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1586] <= mem_n[1586];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1585] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1585] <= mem_n[1585];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1584] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1584] <= mem_n[1584];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1583] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1583] <= mem_n[1583];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1582] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1582] <= mem_n[1582];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1581] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1581] <= mem_n[1581];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1580] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1580] <= mem_n[1580];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1579] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1579] <= mem_n[1579];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1578] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1578] <= mem_n[1578];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1577] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1577] <= mem_n[1577];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1576] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1576] <= mem_n[1576];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1575] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1575] <= mem_n[1575];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1574] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1574] <= mem_n[1574];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1573] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1573] <= mem_n[1573];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1572] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1572] <= mem_n[1572];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1571] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1571] <= mem_n[1571];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1570] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1570] <= mem_n[1570];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1569] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1569] <= mem_n[1569];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1568] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1568] <= mem_n[1568];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1567] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1567] <= mem_n[1567];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1566] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1566] <= mem_n[1566];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1565] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1565] <= mem_n[1565];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1564] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1564] <= mem_n[1564];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1563] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1563] <= mem_n[1563];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1562] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1562] <= mem_n[1562];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1561] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1561] <= mem_n[1561];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1560] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1560] <= mem_n[1560];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1559] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1559] <= mem_n[1559];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1558] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1558] <= mem_n[1558];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1557] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1557] <= mem_n[1557];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1556] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1556] <= mem_n[1556];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1555] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1555] <= mem_n[1555];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1554] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1554] <= mem_n[1554];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1553] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1553] <= mem_n[1553];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1552] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1552] <= mem_n[1552];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1551] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1551] <= mem_n[1551];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1550] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1550] <= mem_n[1550];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1549] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1549] <= mem_n[1549];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1548] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1548] <= mem_n[1548];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1547] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1547] <= mem_n[1547];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1546] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1546] <= mem_n[1546];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1545] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1545] <= mem_n[1545];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1544] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1544] <= mem_n[1544];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1543] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1543] <= mem_n[1543];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1542] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1542] <= mem_n[1542];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1541] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1541] <= mem_n[1541];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1540] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1540] <= mem_n[1540];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1539] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1539] <= mem_n[1539];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1538] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1538] <= mem_n[1538];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1537] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1537] <= mem_n[1537];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1536] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1536] <= mem_n[1536];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1535] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1535] <= mem_n[1535];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1534] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1534] <= mem_n[1534];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1533] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1533] <= mem_n[1533];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1532] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1532] <= mem_n[1532];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1531] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1531] <= mem_n[1531];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1530] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1530] <= mem_n[1530];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1529] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1529] <= mem_n[1529];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1528] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1528] <= mem_n[1528];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1527] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1527] <= mem_n[1527];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1526] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1526] <= mem_n[1526];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1525] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1525] <= mem_n[1525];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1524] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1524] <= mem_n[1524];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1523] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1523] <= mem_n[1523];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1522] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1522] <= mem_n[1522];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1521] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1521] <= mem_n[1521];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1520] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1520] <= mem_n[1520];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1519] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1519] <= mem_n[1519];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1518] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1518] <= mem_n[1518];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1517] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1517] <= mem_n[1517];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1516] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1516] <= mem_n[1516];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1515] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1515] <= mem_n[1515];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1514] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1514] <= mem_n[1514];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1513] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1513] <= mem_n[1513];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1512] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1512] <= mem_n[1512];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1511] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1511] <= mem_n[1511];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1510] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1510] <= mem_n[1510];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1509] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1509] <= mem_n[1509];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1508] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1508] <= mem_n[1508];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1507] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1507] <= mem_n[1507];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1506] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1506] <= mem_n[1506];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1505] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1505] <= mem_n[1505];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1504] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1504] <= mem_n[1504];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1503] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1503] <= mem_n[1503];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1502] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1502] <= mem_n[1502];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1501] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1501] <= mem_n[1501];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1500] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1500] <= mem_n[1500];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1499] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1499] <= mem_n[1499];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1498] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1498] <= mem_n[1498];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1497] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1497] <= mem_n[1497];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1496] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1496] <= mem_n[1496];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1495] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1495] <= mem_n[1495];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1494] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1494] <= mem_n[1494];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1493] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1493] <= mem_n[1493];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1492] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1492] <= mem_n[1492];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1491] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1491] <= mem_n[1491];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1490] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1490] <= mem_n[1490];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1489] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1489] <= mem_n[1489];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1488] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1488] <= mem_n[1488];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1487] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1487] <= mem_n[1487];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1486] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1486] <= mem_n[1486];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1485] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1485] <= mem_n[1485];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1484] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1484] <= mem_n[1484];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1483] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1483] <= mem_n[1483];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1482] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1482] <= mem_n[1482];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1481] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1481] <= mem_n[1481];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1480] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1480] <= mem_n[1480];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1479] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1479] <= mem_n[1479];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1478] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1478] <= mem_n[1478];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1477] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1477] <= mem_n[1477];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1476] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1476] <= mem_n[1476];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1475] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1475] <= mem_n[1475];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1474] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1474] <= mem_n[1474];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1473] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1473] <= mem_n[1473];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1472] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1472] <= mem_n[1472];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1471] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1471] <= mem_n[1471];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1470] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1470] <= mem_n[1470];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1469] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1469] <= mem_n[1469];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1468] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1468] <= mem_n[1468];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1467] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1467] <= mem_n[1467];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1466] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1466] <= mem_n[1466];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1465] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1465] <= mem_n[1465];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1464] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1464] <= mem_n[1464];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1463] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1463] <= mem_n[1463];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1462] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1462] <= mem_n[1462];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1461] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1461] <= mem_n[1461];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1460] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1460] <= mem_n[1460];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1459] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1459] <= mem_n[1459];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1458] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1458] <= mem_n[1458];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1457] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1457] <= mem_n[1457];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1456] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1456] <= mem_n[1456];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1455] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1455] <= mem_n[1455];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1454] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1454] <= mem_n[1454];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1453] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1453] <= mem_n[1453];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1452] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1452] <= mem_n[1452];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1451] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1451] <= mem_n[1451];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1450] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1450] <= mem_n[1450];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1449] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1449] <= mem_n[1449];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1448] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1448] <= mem_n[1448];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1447] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1447] <= mem_n[1447];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1446] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1446] <= mem_n[1446];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1445] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1445] <= mem_n[1445];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1444] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1444] <= mem_n[1444];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1443] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1443] <= mem_n[1443];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1442] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1442] <= mem_n[1442];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1441] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1441] <= mem_n[1441];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1440] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1440] <= mem_n[1440];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1439] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1439] <= mem_n[1439];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1438] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1438] <= mem_n[1438];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1437] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1437] <= mem_n[1437];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1436] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1436] <= mem_n[1436];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1435] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1435] <= mem_n[1435];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1434] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1434] <= mem_n[1434];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1433] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1433] <= mem_n[1433];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1432] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1432] <= mem_n[1432];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1431] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1431] <= mem_n[1431];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1430] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1430] <= mem_n[1430];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1429] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1429] <= mem_n[1429];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1428] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1428] <= mem_n[1428];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1427] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1427] <= mem_n[1427];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1426] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1426] <= mem_n[1426];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1425] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1425] <= mem_n[1425];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1424] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1424] <= mem_n[1424];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1423] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1423] <= mem_n[1423];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1422] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1422] <= mem_n[1422];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1421] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1421] <= mem_n[1421];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1420] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1420] <= mem_n[1420];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1419] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1419] <= mem_n[1419];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1418] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1418] <= mem_n[1418];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1417] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1417] <= mem_n[1417];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1416] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1416] <= mem_n[1416];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1415] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1415] <= mem_n[1415];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1414] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1414] <= mem_n[1414];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1413] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1413] <= mem_n[1413];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1412] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1412] <= mem_n[1412];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1411] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1411] <= mem_n[1411];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1410] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1410] <= mem_n[1410];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1409] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1409] <= mem_n[1409];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1408] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1408] <= mem_n[1408];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1407] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1407] <= mem_n[1407];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1406] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1406] <= mem_n[1406];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1405] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1405] <= mem_n[1405];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1404] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1404] <= mem_n[1404];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1403] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1403] <= mem_n[1403];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1402] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1402] <= mem_n[1402];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1401] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1401] <= mem_n[1401];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1400] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1400] <= mem_n[1400];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1399] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1399] <= mem_n[1399];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1398] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1398] <= mem_n[1398];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1397] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1397] <= mem_n[1397];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1396] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1396] <= mem_n[1396];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1395] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1395] <= mem_n[1395];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1394] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1394] <= mem_n[1394];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1393] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1393] <= mem_n[1393];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1392] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1392] <= mem_n[1392];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1391] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1391] <= mem_n[1391];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1390] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1390] <= mem_n[1390];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1389] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1389] <= mem_n[1389];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1388] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1388] <= mem_n[1388];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1387] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1387] <= mem_n[1387];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1386] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1386] <= mem_n[1386];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1385] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1385] <= mem_n[1385];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1384] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1384] <= mem_n[1384];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1383] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1383] <= mem_n[1383];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1382] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1382] <= mem_n[1382];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1381] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1381] <= mem_n[1381];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1380] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1380] <= mem_n[1380];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1379] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1379] <= mem_n[1379];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1378] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1378] <= mem_n[1378];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1377] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1377] <= mem_n[1377];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1376] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1376] <= mem_n[1376];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1375] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1375] <= mem_n[1375];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1374] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1374] <= mem_n[1374];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1373] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1373] <= mem_n[1373];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1372] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1372] <= mem_n[1372];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1371] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1371] <= mem_n[1371];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1370] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1370] <= mem_n[1370];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1369] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1369] <= mem_n[1369];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1368] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1368] <= mem_n[1368];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1367] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1367] <= mem_n[1367];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1366] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1366] <= mem_n[1366];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1365] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1365] <= mem_n[1365];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1364] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1364] <= mem_n[1364];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1363] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1363] <= mem_n[1363];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1362] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1362] <= mem_n[1362];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1361] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1361] <= mem_n[1361];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1360] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1360] <= mem_n[1360];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1359] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1359] <= mem_n[1359];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1358] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1358] <= mem_n[1358];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1357] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1357] <= mem_n[1357];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1356] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1356] <= mem_n[1356];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1355] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1355] <= mem_n[1355];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1354] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1354] <= mem_n[1354];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1353] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1353] <= mem_n[1353];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1352] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1352] <= mem_n[1352];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1351] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1351] <= mem_n[1351];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1350] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1350] <= mem_n[1350];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1349] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1349] <= mem_n[1349];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1348] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1348] <= mem_n[1348];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1347] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1347] <= mem_n[1347];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1346] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1346] <= mem_n[1346];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1345] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1345] <= mem_n[1345];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1344] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1344] <= mem_n[1344];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1343] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1343] <= mem_n[1343];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1342] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1342] <= mem_n[1342];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1341] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1341] <= mem_n[1341];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1340] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1340] <= mem_n[1340];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1339] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1339] <= mem_n[1339];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1338] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1338] <= mem_n[1338];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1337] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1337] <= mem_n[1337];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1336] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1336] <= mem_n[1336];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1335] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1335] <= mem_n[1335];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1334] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1334] <= mem_n[1334];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1333] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1333] <= mem_n[1333];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1332] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1332] <= mem_n[1332];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1331] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1331] <= mem_n[1331];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1330] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1330] <= mem_n[1330];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1329] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1329] <= mem_n[1329];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1328] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1328] <= mem_n[1328];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1327] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1327] <= mem_n[1327];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1326] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1326] <= mem_n[1326];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1325] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1325] <= mem_n[1325];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1324] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1324] <= mem_n[1324];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1323] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1323] <= mem_n[1323];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1322] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1322] <= mem_n[1322];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1321] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1321] <= mem_n[1321];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1320] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1320] <= mem_n[1320];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1319] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1319] <= mem_n[1319];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1318] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1318] <= mem_n[1318];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1317] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1317] <= mem_n[1317];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1316] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1316] <= mem_n[1316];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1315] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1315] <= mem_n[1315];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1314] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1314] <= mem_n[1314];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1313] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1313] <= mem_n[1313];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1312] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1312] <= mem_n[1312];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1311] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1311] <= mem_n[1311];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1310] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1310] <= mem_n[1310];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1309] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1309] <= mem_n[1309];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1308] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1308] <= mem_n[1308];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1307] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1307] <= mem_n[1307];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1306] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1306] <= mem_n[1306];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1305] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1305] <= mem_n[1305];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1304] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1304] <= mem_n[1304];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1303] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1303] <= mem_n[1303];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1302] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1302] <= mem_n[1302];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1301] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1301] <= mem_n[1301];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1300] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1300] <= mem_n[1300];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1299] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1299] <= mem_n[1299];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1298] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1298] <= mem_n[1298];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1297] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1297] <= mem_n[1297];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1296] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1296] <= mem_n[1296];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1295] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1295] <= mem_n[1295];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1294] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1294] <= mem_n[1294];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1293] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1293] <= mem_n[1293];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1292] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1292] <= mem_n[1292];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1291] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1291] <= mem_n[1291];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1290] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1290] <= mem_n[1290];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1289] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1289] <= mem_n[1289];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1288] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1288] <= mem_n[1288];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1287] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1287] <= mem_n[1287];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1286] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1286] <= mem_n[1286];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1285] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1285] <= mem_n[1285];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1284] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1284] <= mem_n[1284];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1283] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1283] <= mem_n[1283];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1282] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1282] <= mem_n[1282];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1281] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1281] <= mem_n[1281];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1280] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1280] <= mem_n[1280];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1279] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1279] <= mem_n[1279];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1278] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1278] <= mem_n[1278];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1277] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1277] <= mem_n[1277];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1276] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1276] <= mem_n[1276];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1275] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1275] <= mem_n[1275];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1274] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1274] <= mem_n[1274];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1273] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1273] <= mem_n[1273];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1272] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1272] <= mem_n[1272];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1271] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1271] <= mem_n[1271];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1270] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1270] <= mem_n[1270];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1269] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1269] <= mem_n[1269];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1268] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1268] <= mem_n[1268];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1267] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1267] <= mem_n[1267];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1266] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1266] <= mem_n[1266];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1265] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1265] <= mem_n[1265];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1264] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1264] <= mem_n[1264];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1263] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1263] <= mem_n[1263];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1262] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1262] <= mem_n[1262];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1261] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1261] <= mem_n[1261];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1260] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1260] <= mem_n[1260];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1259] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1259] <= mem_n[1259];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1258] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1258] <= mem_n[1258];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1257] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1257] <= mem_n[1257];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1256] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1256] <= mem_n[1256];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1255] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1255] <= mem_n[1255];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1254] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1254] <= mem_n[1254];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1253] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1253] <= mem_n[1253];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1252] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1252] <= mem_n[1252];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1251] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1251] <= mem_n[1251];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1250] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1250] <= mem_n[1250];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1249] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1249] <= mem_n[1249];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1248] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1248] <= mem_n[1248];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1247] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1247] <= mem_n[1247];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1246] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1246] <= mem_n[1246];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1245] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1245] <= mem_n[1245];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1244] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1244] <= mem_n[1244];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1243] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1243] <= mem_n[1243];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1242] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1242] <= mem_n[1242];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1241] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1241] <= mem_n[1241];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1240] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1240] <= mem_n[1240];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1239] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1239] <= mem_n[1239];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1238] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1238] <= mem_n[1238];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1237] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1237] <= mem_n[1237];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1236] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1236] <= mem_n[1236];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1235] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1235] <= mem_n[1235];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1234] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1234] <= mem_n[1234];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1233] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1233] <= mem_n[1233];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1232] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1232] <= mem_n[1232];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1231] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1231] <= mem_n[1231];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1230] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1230] <= mem_n[1230];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1229] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1229] <= mem_n[1229];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1228] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1228] <= mem_n[1228];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1227] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1227] <= mem_n[1227];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1226] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1226] <= mem_n[1226];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1225] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1225] <= mem_n[1225];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1224] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1224] <= mem_n[1224];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1223] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1223] <= mem_n[1223];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1222] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1222] <= mem_n[1222];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1221] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1221] <= mem_n[1221];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1220] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1220] <= mem_n[1220];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1219] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1219] <= mem_n[1219];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1218] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1218] <= mem_n[1218];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1217] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1217] <= mem_n[1217];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1216] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1216] <= mem_n[1216];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1215] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1215] <= mem_n[1215];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1214] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1214] <= mem_n[1214];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1213] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1213] <= mem_n[1213];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1212] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1212] <= mem_n[1212];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1211] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1211] <= mem_n[1211];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1210] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1210] <= mem_n[1210];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1209] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1209] <= mem_n[1209];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1208] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1208] <= mem_n[1208];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1207] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1207] <= mem_n[1207];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1206] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1206] <= mem_n[1206];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1205] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1205] <= mem_n[1205];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1204] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1204] <= mem_n[1204];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1203] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1203] <= mem_n[1203];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1202] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1202] <= mem_n[1202];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1201] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1201] <= mem_n[1201];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1200] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1200] <= mem_n[1200];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1199] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1199] <= mem_n[1199];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1198] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1198] <= mem_n[1198];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1197] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1197] <= mem_n[1197];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1196] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1196] <= mem_n[1196];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1195] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1195] <= mem_n[1195];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1194] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1194] <= mem_n[1194];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1193] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1193] <= mem_n[1193];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1192] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1192] <= mem_n[1192];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1191] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1191] <= mem_n[1191];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1190] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1190] <= mem_n[1190];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1189] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1189] <= mem_n[1189];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1188] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1188] <= mem_n[1188];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1187] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1187] <= mem_n[1187];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1186] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1186] <= mem_n[1186];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1185] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1185] <= mem_n[1185];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1184] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1184] <= mem_n[1184];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1183] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1183] <= mem_n[1183];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1182] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1182] <= mem_n[1182];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1181] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1181] <= mem_n[1181];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1180] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1180] <= mem_n[1180];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1179] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1179] <= mem_n[1179];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1178] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1178] <= mem_n[1178];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1177] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1177] <= mem_n[1177];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1176] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1176] <= mem_n[1176];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1175] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1175] <= mem_n[1175];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1174] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1174] <= mem_n[1174];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1173] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1173] <= mem_n[1173];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1172] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1172] <= mem_n[1172];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1171] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1171] <= mem_n[1171];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1170] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1170] <= mem_n[1170];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1169] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1169] <= mem_n[1169];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1168] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1168] <= mem_n[1168];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1167] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1167] <= mem_n[1167];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1166] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1166] <= mem_n[1166];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1165] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1165] <= mem_n[1165];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1164] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1164] <= mem_n[1164];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1163] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1163] <= mem_n[1163];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1162] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1162] <= mem_n[1162];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1161] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1161] <= mem_n[1161];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1160] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1160] <= mem_n[1160];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1159] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1159] <= mem_n[1159];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1158] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1158] <= mem_n[1158];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1157] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1157] <= mem_n[1157];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1156] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1156] <= mem_n[1156];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1155] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1155] <= mem_n[1155];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1154] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1154] <= mem_n[1154];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1153] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1153] <= mem_n[1153];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1152] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1152] <= mem_n[1152];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1151] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1151] <= mem_n[1151];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1150] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1150] <= mem_n[1150];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1149] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1149] <= mem_n[1149];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1148] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1148] <= mem_n[1148];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1147] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1147] <= mem_n[1147];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1146] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1146] <= mem_n[1146];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1145] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1145] <= mem_n[1145];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1144] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1144] <= mem_n[1144];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1143] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1143] <= mem_n[1143];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1142] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1142] <= mem_n[1142];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1141] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1141] <= mem_n[1141];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1140] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1140] <= mem_n[1140];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1139] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1139] <= mem_n[1139];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1138] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1138] <= mem_n[1138];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1137] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1137] <= mem_n[1137];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1136] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1136] <= mem_n[1136];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1135] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1135] <= mem_n[1135];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1134] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1134] <= mem_n[1134];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1133] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1133] <= mem_n[1133];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1132] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1132] <= mem_n[1132];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1131] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1131] <= mem_n[1131];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1130] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1130] <= mem_n[1130];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1129] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1129] <= mem_n[1129];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1128] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1128] <= mem_n[1128];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1127] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1127] <= mem_n[1127];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1126] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1126] <= mem_n[1126];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1125] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1125] <= mem_n[1125];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1124] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1124] <= mem_n[1124];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1123] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1123] <= mem_n[1123];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1122] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1122] <= mem_n[1122];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1121] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1121] <= mem_n[1121];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1120] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1120] <= mem_n[1120];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1119] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1119] <= mem_n[1119];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1118] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1118] <= mem_n[1118];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1117] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1117] <= mem_n[1117];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1116] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1116] <= mem_n[1116];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1115] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1115] <= mem_n[1115];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1114] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1114] <= mem_n[1114];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1113] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1113] <= mem_n[1113];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1112] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1112] <= mem_n[1112];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1111] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1111] <= mem_n[1111];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1110] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1110] <= mem_n[1110];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1109] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1109] <= mem_n[1109];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1108] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1108] <= mem_n[1108];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1107] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1107] <= mem_n[1107];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1106] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1106] <= mem_n[1106];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1105] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1105] <= mem_n[1105];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1104] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1104] <= mem_n[1104];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1103] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1103] <= mem_n[1103];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1102] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1102] <= mem_n[1102];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1101] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1101] <= mem_n[1101];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1100] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1100] <= mem_n[1100];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1099] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1099] <= mem_n[1099];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1098] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1098] <= mem_n[1098];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1097] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1097] <= mem_n[1097];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1096] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1096] <= mem_n[1096];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1095] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1095] <= mem_n[1095];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1094] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1094] <= mem_n[1094];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1093] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1093] <= mem_n[1093];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1092] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1092] <= mem_n[1092];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1091] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1091] <= mem_n[1091];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1090] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1090] <= mem_n[1090];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1089] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1089] <= mem_n[1089];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1088] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1088] <= mem_n[1088];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1087] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1087] <= mem_n[1087];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1086] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1086] <= mem_n[1086];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1085] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1085] <= mem_n[1085];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1084] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1084] <= mem_n[1084];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1083] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1083] <= mem_n[1083];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1082] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1082] <= mem_n[1082];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1081] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1081] <= mem_n[1081];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1080] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1080] <= mem_n[1080];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1079] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1079] <= mem_n[1079];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1078] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1078] <= mem_n[1078];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1077] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1077] <= mem_n[1077];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1076] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1076] <= mem_n[1076];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1075] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1075] <= mem_n[1075];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1074] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1074] <= mem_n[1074];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1073] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1073] <= mem_n[1073];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1072] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1072] <= mem_n[1072];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1071] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1071] <= mem_n[1071];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1070] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1070] <= mem_n[1070];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1069] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1069] <= mem_n[1069];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1068] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1068] <= mem_n[1068];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1067] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1067] <= mem_n[1067];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1066] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1066] <= mem_n[1066];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1065] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1065] <= mem_n[1065];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1064] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1064] <= mem_n[1064];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1063] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1063] <= mem_n[1063];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1062] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1062] <= mem_n[1062];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1061] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1061] <= mem_n[1061];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1060] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1060] <= mem_n[1060];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1059] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1059] <= mem_n[1059];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1058] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1058] <= mem_n[1058];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1057] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1057] <= mem_n[1057];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1056] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1056] <= mem_n[1056];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1055] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1055] <= mem_n[1055];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1054] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1054] <= mem_n[1054];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1053] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1053] <= mem_n[1053];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1052] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1052] <= mem_n[1052];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1051] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1051] <= mem_n[1051];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1050] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1050] <= mem_n[1050];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1049] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1049] <= mem_n[1049];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1048] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1048] <= mem_n[1048];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1047] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1047] <= mem_n[1047];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1046] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1046] <= mem_n[1046];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1045] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1045] <= mem_n[1045];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1044] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1044] <= mem_n[1044];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1043] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1043] <= mem_n[1043];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1042] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1042] <= mem_n[1042];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1041] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1041] <= mem_n[1041];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1040] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1040] <= mem_n[1040];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1039] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1039] <= mem_n[1039];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1038] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1038] <= mem_n[1038];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1037] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1037] <= mem_n[1037];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1036] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1036] <= mem_n[1036];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1035] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1035] <= mem_n[1035];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1034] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1034] <= mem_n[1034];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1033] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1033] <= mem_n[1033];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1032] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1032] <= mem_n[1032];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1031] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1031] <= mem_n[1031];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1030] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1030] <= mem_n[1030];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1029] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1029] <= mem_n[1029];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1028] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1028] <= mem_n[1028];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1027] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1027] <= mem_n[1027];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1026] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1026] <= mem_n[1026];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1025] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1025] <= mem_n[1025];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1024] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1024] <= mem_n[1024];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1023] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1023] <= mem_n[1023];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1022] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1022] <= mem_n[1022];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1021] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1021] <= mem_n[1021];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1020] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1020] <= mem_n[1020];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1019] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1019] <= mem_n[1019];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1018] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1018] <= mem_n[1018];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1017] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1017] <= mem_n[1017];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1016] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1016] <= mem_n[1016];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1015] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1015] <= mem_n[1015];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1014] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1014] <= mem_n[1014];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1013] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1013] <= mem_n[1013];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1012] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1012] <= mem_n[1012];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1011] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1011] <= mem_n[1011];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1010] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1010] <= mem_n[1010];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1009] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1009] <= mem_n[1009];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1008] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1008] <= mem_n[1008];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1007] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1007] <= mem_n[1007];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1006] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1006] <= mem_n[1006];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1005] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1005] <= mem_n[1005];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1004] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1004] <= mem_n[1004];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1003] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1003] <= mem_n[1003];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1002] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1002] <= mem_n[1002];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1001] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1001] <= mem_n[1001];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1000] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1000] <= mem_n[1000];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[999] <= 1'b0;
    end else if(1'b1) begin
      mem_q[999] <= mem_n[999];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[998] <= 1'b0;
    end else if(1'b1) begin
      mem_q[998] <= mem_n[998];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[997] <= 1'b0;
    end else if(1'b1) begin
      mem_q[997] <= mem_n[997];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[996] <= 1'b0;
    end else if(1'b1) begin
      mem_q[996] <= mem_n[996];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[995] <= 1'b0;
    end else if(1'b1) begin
      mem_q[995] <= mem_n[995];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[994] <= 1'b0;
    end else if(1'b1) begin
      mem_q[994] <= mem_n[994];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[993] <= 1'b0;
    end else if(1'b1) begin
      mem_q[993] <= mem_n[993];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[992] <= 1'b0;
    end else if(1'b1) begin
      mem_q[992] <= mem_n[992];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[991] <= 1'b0;
    end else if(1'b1) begin
      mem_q[991] <= mem_n[991];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[990] <= 1'b0;
    end else if(1'b1) begin
      mem_q[990] <= mem_n[990];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[989] <= 1'b0;
    end else if(1'b1) begin
      mem_q[989] <= mem_n[989];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[988] <= 1'b0;
    end else if(1'b1) begin
      mem_q[988] <= mem_n[988];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[987] <= 1'b0;
    end else if(1'b1) begin
      mem_q[987] <= mem_n[987];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[986] <= 1'b0;
    end else if(1'b1) begin
      mem_q[986] <= mem_n[986];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[985] <= 1'b0;
    end else if(1'b1) begin
      mem_q[985] <= mem_n[985];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[984] <= 1'b0;
    end else if(1'b1) begin
      mem_q[984] <= mem_n[984];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[983] <= 1'b0;
    end else if(1'b1) begin
      mem_q[983] <= mem_n[983];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[982] <= 1'b0;
    end else if(1'b1) begin
      mem_q[982] <= mem_n[982];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[981] <= 1'b0;
    end else if(1'b1) begin
      mem_q[981] <= mem_n[981];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[980] <= 1'b0;
    end else if(1'b1) begin
      mem_q[980] <= mem_n[980];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[979] <= 1'b0;
    end else if(1'b1) begin
      mem_q[979] <= mem_n[979];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[978] <= 1'b0;
    end else if(1'b1) begin
      mem_q[978] <= mem_n[978];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[977] <= 1'b0;
    end else if(1'b1) begin
      mem_q[977] <= mem_n[977];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[976] <= 1'b0;
    end else if(1'b1) begin
      mem_q[976] <= mem_n[976];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[975] <= 1'b0;
    end else if(1'b1) begin
      mem_q[975] <= mem_n[975];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[974] <= 1'b0;
    end else if(1'b1) begin
      mem_q[974] <= mem_n[974];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[973] <= 1'b0;
    end else if(1'b1) begin
      mem_q[973] <= mem_n[973];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[972] <= 1'b0;
    end else if(1'b1) begin
      mem_q[972] <= mem_n[972];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[971] <= 1'b0;
    end else if(1'b1) begin
      mem_q[971] <= mem_n[971];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[970] <= 1'b0;
    end else if(1'b1) begin
      mem_q[970] <= mem_n[970];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[969] <= 1'b0;
    end else if(1'b1) begin
      mem_q[969] <= mem_n[969];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[968] <= 1'b0;
    end else if(1'b1) begin
      mem_q[968] <= mem_n[968];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[967] <= 1'b0;
    end else if(1'b1) begin
      mem_q[967] <= mem_n[967];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[966] <= 1'b0;
    end else if(1'b1) begin
      mem_q[966] <= mem_n[966];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[965] <= 1'b0;
    end else if(1'b1) begin
      mem_q[965] <= mem_n[965];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[964] <= 1'b0;
    end else if(1'b1) begin
      mem_q[964] <= mem_n[964];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[963] <= 1'b0;
    end else if(1'b1) begin
      mem_q[963] <= mem_n[963];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[962] <= 1'b0;
    end else if(1'b1) begin
      mem_q[962] <= mem_n[962];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[961] <= 1'b0;
    end else if(1'b1) begin
      mem_q[961] <= mem_n[961];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[960] <= 1'b0;
    end else if(1'b1) begin
      mem_q[960] <= mem_n[960];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[959] <= 1'b0;
    end else if(1'b1) begin
      mem_q[959] <= mem_n[959];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[958] <= 1'b0;
    end else if(1'b1) begin
      mem_q[958] <= mem_n[958];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[957] <= 1'b0;
    end else if(1'b1) begin
      mem_q[957] <= mem_n[957];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[956] <= 1'b0;
    end else if(1'b1) begin
      mem_q[956] <= mem_n[956];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[955] <= 1'b0;
    end else if(1'b1) begin
      mem_q[955] <= mem_n[955];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[954] <= 1'b0;
    end else if(1'b1) begin
      mem_q[954] <= mem_n[954];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[953] <= 1'b0;
    end else if(1'b1) begin
      mem_q[953] <= mem_n[953];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[952] <= 1'b0;
    end else if(1'b1) begin
      mem_q[952] <= mem_n[952];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[951] <= 1'b0;
    end else if(1'b1) begin
      mem_q[951] <= mem_n[951];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[950] <= 1'b0;
    end else if(1'b1) begin
      mem_q[950] <= mem_n[950];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[949] <= 1'b0;
    end else if(1'b1) begin
      mem_q[949] <= mem_n[949];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[948] <= 1'b0;
    end else if(1'b1) begin
      mem_q[948] <= mem_n[948];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[947] <= 1'b0;
    end else if(1'b1) begin
      mem_q[947] <= mem_n[947];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[946] <= 1'b0;
    end else if(1'b1) begin
      mem_q[946] <= mem_n[946];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[945] <= 1'b0;
    end else if(1'b1) begin
      mem_q[945] <= mem_n[945];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[944] <= 1'b0;
    end else if(1'b1) begin
      mem_q[944] <= mem_n[944];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[943] <= 1'b0;
    end else if(1'b1) begin
      mem_q[943] <= mem_n[943];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[942] <= 1'b0;
    end else if(1'b1) begin
      mem_q[942] <= mem_n[942];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[941] <= 1'b0;
    end else if(1'b1) begin
      mem_q[941] <= mem_n[941];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[940] <= 1'b0;
    end else if(1'b1) begin
      mem_q[940] <= mem_n[940];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[939] <= 1'b0;
    end else if(1'b1) begin
      mem_q[939] <= mem_n[939];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[938] <= 1'b0;
    end else if(1'b1) begin
      mem_q[938] <= mem_n[938];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[937] <= 1'b0;
    end else if(1'b1) begin
      mem_q[937] <= mem_n[937];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[936] <= 1'b0;
    end else if(1'b1) begin
      mem_q[936] <= mem_n[936];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[935] <= 1'b0;
    end else if(1'b1) begin
      mem_q[935] <= mem_n[935];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[934] <= 1'b0;
    end else if(1'b1) begin
      mem_q[934] <= mem_n[934];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[933] <= 1'b0;
    end else if(1'b1) begin
      mem_q[933] <= mem_n[933];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[932] <= 1'b0;
    end else if(1'b1) begin
      mem_q[932] <= mem_n[932];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[931] <= 1'b0;
    end else if(1'b1) begin
      mem_q[931] <= mem_n[931];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[930] <= 1'b0;
    end else if(1'b1) begin
      mem_q[930] <= mem_n[930];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[929] <= 1'b0;
    end else if(1'b1) begin
      mem_q[929] <= mem_n[929];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[928] <= 1'b0;
    end else if(1'b1) begin
      mem_q[928] <= mem_n[928];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[927] <= 1'b0;
    end else if(1'b1) begin
      mem_q[927] <= mem_n[927];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[926] <= 1'b0;
    end else if(1'b1) begin
      mem_q[926] <= mem_n[926];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[925] <= 1'b0;
    end else if(1'b1) begin
      mem_q[925] <= mem_n[925];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[924] <= 1'b0;
    end else if(1'b1) begin
      mem_q[924] <= mem_n[924];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[923] <= 1'b0;
    end else if(1'b1) begin
      mem_q[923] <= mem_n[923];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[922] <= 1'b0;
    end else if(1'b1) begin
      mem_q[922] <= mem_n[922];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[921] <= 1'b0;
    end else if(1'b1) begin
      mem_q[921] <= mem_n[921];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[920] <= 1'b0;
    end else if(1'b1) begin
      mem_q[920] <= mem_n[920];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[919] <= 1'b0;
    end else if(1'b1) begin
      mem_q[919] <= mem_n[919];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[918] <= 1'b0;
    end else if(1'b1) begin
      mem_q[918] <= mem_n[918];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[917] <= 1'b0;
    end else if(1'b1) begin
      mem_q[917] <= mem_n[917];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[916] <= 1'b0;
    end else if(1'b1) begin
      mem_q[916] <= mem_n[916];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[915] <= 1'b0;
    end else if(1'b1) begin
      mem_q[915] <= mem_n[915];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[914] <= 1'b0;
    end else if(1'b1) begin
      mem_q[914] <= mem_n[914];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[913] <= 1'b0;
    end else if(1'b1) begin
      mem_q[913] <= mem_n[913];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[912] <= 1'b0;
    end else if(1'b1) begin
      mem_q[912] <= mem_n[912];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[911] <= 1'b0;
    end else if(1'b1) begin
      mem_q[911] <= mem_n[911];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[910] <= 1'b0;
    end else if(1'b1) begin
      mem_q[910] <= mem_n[910];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[909] <= 1'b0;
    end else if(1'b1) begin
      mem_q[909] <= mem_n[909];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[908] <= 1'b0;
    end else if(1'b1) begin
      mem_q[908] <= mem_n[908];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[907] <= 1'b0;
    end else if(1'b1) begin
      mem_q[907] <= mem_n[907];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[906] <= 1'b0;
    end else if(1'b1) begin
      mem_q[906] <= mem_n[906];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[905] <= 1'b0;
    end else if(1'b1) begin
      mem_q[905] <= mem_n[905];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[904] <= 1'b0;
    end else if(1'b1) begin
      mem_q[904] <= mem_n[904];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[903] <= 1'b0;
    end else if(1'b1) begin
      mem_q[903] <= mem_n[903];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[902] <= 1'b0;
    end else if(1'b1) begin
      mem_q[902] <= mem_n[902];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[901] <= 1'b0;
    end else if(1'b1) begin
      mem_q[901] <= mem_n[901];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[900] <= 1'b0;
    end else if(1'b1) begin
      mem_q[900] <= mem_n[900];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[899] <= 1'b0;
    end else if(1'b1) begin
      mem_q[899] <= mem_n[899];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[898] <= 1'b0;
    end else if(1'b1) begin
      mem_q[898] <= mem_n[898];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[897] <= 1'b0;
    end else if(1'b1) begin
      mem_q[897] <= mem_n[897];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[896] <= 1'b0;
    end else if(1'b1) begin
      mem_q[896] <= mem_n[896];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[895] <= 1'b0;
    end else if(1'b1) begin
      mem_q[895] <= mem_n[895];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[894] <= 1'b0;
    end else if(1'b1) begin
      mem_q[894] <= mem_n[894];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[893] <= 1'b0;
    end else if(1'b1) begin
      mem_q[893] <= mem_n[893];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[892] <= 1'b0;
    end else if(1'b1) begin
      mem_q[892] <= mem_n[892];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[891] <= 1'b0;
    end else if(1'b1) begin
      mem_q[891] <= mem_n[891];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[890] <= 1'b0;
    end else if(1'b1) begin
      mem_q[890] <= mem_n[890];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[889] <= 1'b0;
    end else if(1'b1) begin
      mem_q[889] <= mem_n[889];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[888] <= 1'b0;
    end else if(1'b1) begin
      mem_q[888] <= mem_n[888];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[887] <= 1'b0;
    end else if(1'b1) begin
      mem_q[887] <= mem_n[887];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[886] <= 1'b0;
    end else if(1'b1) begin
      mem_q[886] <= mem_n[886];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[885] <= 1'b0;
    end else if(1'b1) begin
      mem_q[885] <= mem_n[885];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[884] <= 1'b0;
    end else if(1'b1) begin
      mem_q[884] <= mem_n[884];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[883] <= 1'b0;
    end else if(1'b1) begin
      mem_q[883] <= mem_n[883];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[882] <= 1'b0;
    end else if(1'b1) begin
      mem_q[882] <= mem_n[882];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[881] <= 1'b0;
    end else if(1'b1) begin
      mem_q[881] <= mem_n[881];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[880] <= 1'b0;
    end else if(1'b1) begin
      mem_q[880] <= mem_n[880];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[879] <= 1'b0;
    end else if(1'b1) begin
      mem_q[879] <= mem_n[879];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[878] <= 1'b0;
    end else if(1'b1) begin
      mem_q[878] <= mem_n[878];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[877] <= 1'b0;
    end else if(1'b1) begin
      mem_q[877] <= mem_n[877];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[876] <= 1'b0;
    end else if(1'b1) begin
      mem_q[876] <= mem_n[876];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[875] <= 1'b0;
    end else if(1'b1) begin
      mem_q[875] <= mem_n[875];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[874] <= 1'b0;
    end else if(1'b1) begin
      mem_q[874] <= mem_n[874];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[873] <= 1'b0;
    end else if(1'b1) begin
      mem_q[873] <= mem_n[873];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[872] <= 1'b0;
    end else if(1'b1) begin
      mem_q[872] <= mem_n[872];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[871] <= 1'b0;
    end else if(1'b1) begin
      mem_q[871] <= mem_n[871];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[870] <= 1'b0;
    end else if(1'b1) begin
      mem_q[870] <= mem_n[870];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[869] <= 1'b0;
    end else if(1'b1) begin
      mem_q[869] <= mem_n[869];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[868] <= 1'b0;
    end else if(1'b1) begin
      mem_q[868] <= mem_n[868];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[867] <= 1'b0;
    end else if(1'b1) begin
      mem_q[867] <= mem_n[867];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[866] <= 1'b0;
    end else if(1'b1) begin
      mem_q[866] <= mem_n[866];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[865] <= 1'b0;
    end else if(1'b1) begin
      mem_q[865] <= mem_n[865];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[864] <= 1'b0;
    end else if(1'b1) begin
      mem_q[864] <= mem_n[864];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[863] <= 1'b0;
    end else if(1'b1) begin
      mem_q[863] <= mem_n[863];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[862] <= 1'b0;
    end else if(1'b1) begin
      mem_q[862] <= mem_n[862];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[861] <= 1'b0;
    end else if(1'b1) begin
      mem_q[861] <= mem_n[861];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[860] <= 1'b0;
    end else if(1'b1) begin
      mem_q[860] <= mem_n[860];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[859] <= 1'b0;
    end else if(1'b1) begin
      mem_q[859] <= mem_n[859];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[858] <= 1'b0;
    end else if(1'b1) begin
      mem_q[858] <= mem_n[858];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[857] <= 1'b0;
    end else if(1'b1) begin
      mem_q[857] <= mem_n[857];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[856] <= 1'b0;
    end else if(1'b1) begin
      mem_q[856] <= mem_n[856];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[855] <= 1'b0;
    end else if(1'b1) begin
      mem_q[855] <= mem_n[855];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[854] <= 1'b0;
    end else if(1'b1) begin
      mem_q[854] <= mem_n[854];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[853] <= 1'b0;
    end else if(1'b1) begin
      mem_q[853] <= mem_n[853];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[852] <= 1'b0;
    end else if(1'b1) begin
      mem_q[852] <= mem_n[852];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[851] <= 1'b0;
    end else if(1'b1) begin
      mem_q[851] <= mem_n[851];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[850] <= 1'b0;
    end else if(1'b1) begin
      mem_q[850] <= mem_n[850];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[849] <= 1'b0;
    end else if(1'b1) begin
      mem_q[849] <= mem_n[849];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[848] <= 1'b0;
    end else if(1'b1) begin
      mem_q[848] <= mem_n[848];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[847] <= 1'b0;
    end else if(1'b1) begin
      mem_q[847] <= mem_n[847];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[846] <= 1'b0;
    end else if(1'b1) begin
      mem_q[846] <= mem_n[846];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[845] <= 1'b0;
    end else if(1'b1) begin
      mem_q[845] <= mem_n[845];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[844] <= 1'b0;
    end else if(1'b1) begin
      mem_q[844] <= mem_n[844];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[843] <= 1'b0;
    end else if(1'b1) begin
      mem_q[843] <= mem_n[843];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[842] <= 1'b0;
    end else if(1'b1) begin
      mem_q[842] <= mem_n[842];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[841] <= 1'b0;
    end else if(1'b1) begin
      mem_q[841] <= mem_n[841];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[840] <= 1'b0;
    end else if(1'b1) begin
      mem_q[840] <= mem_n[840];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[839] <= 1'b0;
    end else if(1'b1) begin
      mem_q[839] <= mem_n[839];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[838] <= 1'b0;
    end else if(1'b1) begin
      mem_q[838] <= mem_n[838];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[837] <= 1'b0;
    end else if(1'b1) begin
      mem_q[837] <= mem_n[837];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[836] <= 1'b0;
    end else if(1'b1) begin
      mem_q[836] <= mem_n[836];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[835] <= 1'b0;
    end else if(1'b1) begin
      mem_q[835] <= mem_n[835];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[834] <= 1'b0;
    end else if(1'b1) begin
      mem_q[834] <= mem_n[834];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[833] <= 1'b0;
    end else if(1'b1) begin
      mem_q[833] <= mem_n[833];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[832] <= 1'b0;
    end else if(1'b1) begin
      mem_q[832] <= mem_n[832];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[831] <= 1'b0;
    end else if(1'b1) begin
      mem_q[831] <= mem_n[831];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[830] <= 1'b0;
    end else if(1'b1) begin
      mem_q[830] <= mem_n[830];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[829] <= 1'b0;
    end else if(1'b1) begin
      mem_q[829] <= mem_n[829];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[828] <= 1'b0;
    end else if(1'b1) begin
      mem_q[828] <= mem_n[828];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[827] <= 1'b0;
    end else if(1'b1) begin
      mem_q[827] <= mem_n[827];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[826] <= 1'b0;
    end else if(1'b1) begin
      mem_q[826] <= mem_n[826];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[825] <= 1'b0;
    end else if(1'b1) begin
      mem_q[825] <= mem_n[825];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[824] <= 1'b0;
    end else if(1'b1) begin
      mem_q[824] <= mem_n[824];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[823] <= 1'b0;
    end else if(1'b1) begin
      mem_q[823] <= mem_n[823];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[822] <= 1'b0;
    end else if(1'b1) begin
      mem_q[822] <= mem_n[822];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[821] <= 1'b0;
    end else if(1'b1) begin
      mem_q[821] <= mem_n[821];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[820] <= 1'b0;
    end else if(1'b1) begin
      mem_q[820] <= mem_n[820];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[819] <= 1'b0;
    end else if(1'b1) begin
      mem_q[819] <= mem_n[819];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[818] <= 1'b0;
    end else if(1'b1) begin
      mem_q[818] <= mem_n[818];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[817] <= 1'b0;
    end else if(1'b1) begin
      mem_q[817] <= mem_n[817];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[816] <= 1'b0;
    end else if(1'b1) begin
      mem_q[816] <= mem_n[816];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[815] <= 1'b0;
    end else if(1'b1) begin
      mem_q[815] <= mem_n[815];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[814] <= 1'b0;
    end else if(1'b1) begin
      mem_q[814] <= mem_n[814];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[813] <= 1'b0;
    end else if(1'b1) begin
      mem_q[813] <= mem_n[813];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[812] <= 1'b0;
    end else if(1'b1) begin
      mem_q[812] <= mem_n[812];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[811] <= 1'b0;
    end else if(1'b1) begin
      mem_q[811] <= mem_n[811];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[810] <= 1'b0;
    end else if(1'b1) begin
      mem_q[810] <= mem_n[810];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[809] <= 1'b0;
    end else if(1'b1) begin
      mem_q[809] <= mem_n[809];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[808] <= 1'b0;
    end else if(1'b1) begin
      mem_q[808] <= mem_n[808];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[807] <= 1'b0;
    end else if(1'b1) begin
      mem_q[807] <= mem_n[807];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[806] <= 1'b0;
    end else if(1'b1) begin
      mem_q[806] <= mem_n[806];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[805] <= 1'b0;
    end else if(1'b1) begin
      mem_q[805] <= mem_n[805];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[804] <= 1'b0;
    end else if(1'b1) begin
      mem_q[804] <= mem_n[804];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[803] <= 1'b0;
    end else if(1'b1) begin
      mem_q[803] <= mem_n[803];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[802] <= 1'b0;
    end else if(1'b1) begin
      mem_q[802] <= mem_n[802];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[801] <= 1'b0;
    end else if(1'b1) begin
      mem_q[801] <= mem_n[801];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[800] <= 1'b0;
    end else if(1'b1) begin
      mem_q[800] <= mem_n[800];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[799] <= 1'b0;
    end else if(1'b1) begin
      mem_q[799] <= mem_n[799];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[798] <= 1'b0;
    end else if(1'b1) begin
      mem_q[798] <= mem_n[798];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[797] <= 1'b0;
    end else if(1'b1) begin
      mem_q[797] <= mem_n[797];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[796] <= 1'b0;
    end else if(1'b1) begin
      mem_q[796] <= mem_n[796];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[795] <= 1'b0;
    end else if(1'b1) begin
      mem_q[795] <= mem_n[795];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[794] <= 1'b0;
    end else if(1'b1) begin
      mem_q[794] <= mem_n[794];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[793] <= 1'b0;
    end else if(1'b1) begin
      mem_q[793] <= mem_n[793];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[792] <= 1'b0;
    end else if(1'b1) begin
      mem_q[792] <= mem_n[792];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[791] <= 1'b0;
    end else if(1'b1) begin
      mem_q[791] <= mem_n[791];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[790] <= 1'b0;
    end else if(1'b1) begin
      mem_q[790] <= mem_n[790];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[789] <= 1'b0;
    end else if(1'b1) begin
      mem_q[789] <= mem_n[789];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[788] <= 1'b0;
    end else if(1'b1) begin
      mem_q[788] <= mem_n[788];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[787] <= 1'b0;
    end else if(1'b1) begin
      mem_q[787] <= mem_n[787];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[786] <= 1'b0;
    end else if(1'b1) begin
      mem_q[786] <= mem_n[786];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[785] <= 1'b0;
    end else if(1'b1) begin
      mem_q[785] <= mem_n[785];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[784] <= 1'b0;
    end else if(1'b1) begin
      mem_q[784] <= mem_n[784];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[783] <= 1'b0;
    end else if(1'b1) begin
      mem_q[783] <= mem_n[783];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[782] <= 1'b0;
    end else if(1'b1) begin
      mem_q[782] <= mem_n[782];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[781] <= 1'b0;
    end else if(1'b1) begin
      mem_q[781] <= mem_n[781];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[780] <= 1'b0;
    end else if(1'b1) begin
      mem_q[780] <= mem_n[780];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[779] <= 1'b0;
    end else if(1'b1) begin
      mem_q[779] <= mem_n[779];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[778] <= 1'b0;
    end else if(1'b1) begin
      mem_q[778] <= mem_n[778];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[777] <= 1'b0;
    end else if(1'b1) begin
      mem_q[777] <= mem_n[777];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[776] <= 1'b0;
    end else if(1'b1) begin
      mem_q[776] <= mem_n[776];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[775] <= 1'b0;
    end else if(1'b1) begin
      mem_q[775] <= mem_n[775];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[774] <= 1'b0;
    end else if(1'b1) begin
      mem_q[774] <= mem_n[774];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[773] <= 1'b0;
    end else if(1'b1) begin
      mem_q[773] <= mem_n[773];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[772] <= 1'b0;
    end else if(1'b1) begin
      mem_q[772] <= mem_n[772];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[771] <= 1'b0;
    end else if(1'b1) begin
      mem_q[771] <= mem_n[771];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[770] <= 1'b0;
    end else if(1'b1) begin
      mem_q[770] <= mem_n[770];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[769] <= 1'b0;
    end else if(1'b1) begin
      mem_q[769] <= mem_n[769];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[768] <= 1'b0;
    end else if(1'b1) begin
      mem_q[768] <= mem_n[768];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[767] <= 1'b0;
    end else if(1'b1) begin
      mem_q[767] <= mem_n[767];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[766] <= 1'b0;
    end else if(1'b1) begin
      mem_q[766] <= mem_n[766];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[765] <= 1'b0;
    end else if(1'b1) begin
      mem_q[765] <= mem_n[765];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[764] <= 1'b0;
    end else if(1'b1) begin
      mem_q[764] <= mem_n[764];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[763] <= 1'b0;
    end else if(1'b1) begin
      mem_q[763] <= mem_n[763];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[762] <= 1'b0;
    end else if(1'b1) begin
      mem_q[762] <= mem_n[762];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[761] <= 1'b0;
    end else if(1'b1) begin
      mem_q[761] <= mem_n[761];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[760] <= 1'b0;
    end else if(1'b1) begin
      mem_q[760] <= mem_n[760];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[759] <= 1'b0;
    end else if(1'b1) begin
      mem_q[759] <= mem_n[759];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[758] <= 1'b0;
    end else if(1'b1) begin
      mem_q[758] <= mem_n[758];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[757] <= 1'b0;
    end else if(1'b1) begin
      mem_q[757] <= mem_n[757];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[756] <= 1'b0;
    end else if(1'b1) begin
      mem_q[756] <= mem_n[756];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[755] <= 1'b0;
    end else if(1'b1) begin
      mem_q[755] <= mem_n[755];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[754] <= 1'b0;
    end else if(1'b1) begin
      mem_q[754] <= mem_n[754];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[753] <= 1'b0;
    end else if(1'b1) begin
      mem_q[753] <= mem_n[753];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[752] <= 1'b0;
    end else if(1'b1) begin
      mem_q[752] <= mem_n[752];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[751] <= 1'b0;
    end else if(1'b1) begin
      mem_q[751] <= mem_n[751];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[750] <= 1'b0;
    end else if(1'b1) begin
      mem_q[750] <= mem_n[750];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[749] <= 1'b0;
    end else if(1'b1) begin
      mem_q[749] <= mem_n[749];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[748] <= 1'b0;
    end else if(1'b1) begin
      mem_q[748] <= mem_n[748];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[747] <= 1'b0;
    end else if(1'b1) begin
      mem_q[747] <= mem_n[747];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[746] <= 1'b0;
    end else if(1'b1) begin
      mem_q[746] <= mem_n[746];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[745] <= 1'b0;
    end else if(1'b1) begin
      mem_q[745] <= mem_n[745];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[744] <= 1'b0;
    end else if(1'b1) begin
      mem_q[744] <= mem_n[744];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[743] <= 1'b0;
    end else if(1'b1) begin
      mem_q[743] <= mem_n[743];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[742] <= 1'b0;
    end else if(1'b1) begin
      mem_q[742] <= mem_n[742];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[741] <= 1'b0;
    end else if(1'b1) begin
      mem_q[741] <= mem_n[741];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[740] <= 1'b0;
    end else if(1'b1) begin
      mem_q[740] <= mem_n[740];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[739] <= 1'b0;
    end else if(1'b1) begin
      mem_q[739] <= mem_n[739];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[738] <= 1'b0;
    end else if(1'b1) begin
      mem_q[738] <= mem_n[738];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[737] <= 1'b0;
    end else if(1'b1) begin
      mem_q[737] <= mem_n[737];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[736] <= 1'b0;
    end else if(1'b1) begin
      mem_q[736] <= mem_n[736];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[735] <= 1'b0;
    end else if(1'b1) begin
      mem_q[735] <= mem_n[735];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[734] <= 1'b0;
    end else if(1'b1) begin
      mem_q[734] <= mem_n[734];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[733] <= 1'b0;
    end else if(1'b1) begin
      mem_q[733] <= mem_n[733];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[732] <= 1'b0;
    end else if(1'b1) begin
      mem_q[732] <= mem_n[732];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[731] <= 1'b0;
    end else if(1'b1) begin
      mem_q[731] <= mem_n[731];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[730] <= 1'b0;
    end else if(1'b1) begin
      mem_q[730] <= mem_n[730];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[729] <= 1'b0;
    end else if(1'b1) begin
      mem_q[729] <= mem_n[729];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[728] <= 1'b0;
    end else if(1'b1) begin
      mem_q[728] <= mem_n[728];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[727] <= 1'b0;
    end else if(1'b1) begin
      mem_q[727] <= mem_n[727];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[726] <= 1'b0;
    end else if(1'b1) begin
      mem_q[726] <= mem_n[726];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[725] <= 1'b0;
    end else if(1'b1) begin
      mem_q[725] <= mem_n[725];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[724] <= 1'b0;
    end else if(1'b1) begin
      mem_q[724] <= mem_n[724];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[723] <= 1'b0;
    end else if(1'b1) begin
      mem_q[723] <= mem_n[723];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[722] <= 1'b0;
    end else if(1'b1) begin
      mem_q[722] <= mem_n[722];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[721] <= 1'b0;
    end else if(1'b1) begin
      mem_q[721] <= mem_n[721];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[720] <= 1'b0;
    end else if(1'b1) begin
      mem_q[720] <= mem_n[720];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[719] <= 1'b0;
    end else if(1'b1) begin
      mem_q[719] <= mem_n[719];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[718] <= 1'b0;
    end else if(1'b1) begin
      mem_q[718] <= mem_n[718];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[717] <= 1'b0;
    end else if(1'b1) begin
      mem_q[717] <= mem_n[717];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[716] <= 1'b0;
    end else if(1'b1) begin
      mem_q[716] <= mem_n[716];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[715] <= 1'b0;
    end else if(1'b1) begin
      mem_q[715] <= mem_n[715];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[714] <= 1'b0;
    end else if(1'b1) begin
      mem_q[714] <= mem_n[714];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[713] <= 1'b0;
    end else if(1'b1) begin
      mem_q[713] <= mem_n[713];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[712] <= 1'b0;
    end else if(1'b1) begin
      mem_q[712] <= mem_n[712];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[711] <= 1'b0;
    end else if(1'b1) begin
      mem_q[711] <= mem_n[711];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[710] <= 1'b0;
    end else if(1'b1) begin
      mem_q[710] <= mem_n[710];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[709] <= 1'b0;
    end else if(1'b1) begin
      mem_q[709] <= mem_n[709];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[708] <= 1'b0;
    end else if(1'b1) begin
      mem_q[708] <= mem_n[708];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[707] <= 1'b0;
    end else if(1'b1) begin
      mem_q[707] <= mem_n[707];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[706] <= 1'b0;
    end else if(1'b1) begin
      mem_q[706] <= mem_n[706];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[705] <= 1'b0;
    end else if(1'b1) begin
      mem_q[705] <= mem_n[705];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[704] <= 1'b0;
    end else if(1'b1) begin
      mem_q[704] <= mem_n[704];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[703] <= 1'b0;
    end else if(1'b1) begin
      mem_q[703] <= mem_n[703];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[702] <= 1'b0;
    end else if(1'b1) begin
      mem_q[702] <= mem_n[702];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[701] <= 1'b0;
    end else if(1'b1) begin
      mem_q[701] <= mem_n[701];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[700] <= 1'b0;
    end else if(1'b1) begin
      mem_q[700] <= mem_n[700];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[699] <= 1'b0;
    end else if(1'b1) begin
      mem_q[699] <= mem_n[699];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[698] <= 1'b0;
    end else if(1'b1) begin
      mem_q[698] <= mem_n[698];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[697] <= 1'b0;
    end else if(1'b1) begin
      mem_q[697] <= mem_n[697];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[696] <= 1'b0;
    end else if(1'b1) begin
      mem_q[696] <= mem_n[696];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[695] <= 1'b0;
    end else if(1'b1) begin
      mem_q[695] <= mem_n[695];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[694] <= 1'b0;
    end else if(1'b1) begin
      mem_q[694] <= mem_n[694];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[693] <= 1'b0;
    end else if(1'b1) begin
      mem_q[693] <= mem_n[693];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[692] <= 1'b0;
    end else if(1'b1) begin
      mem_q[692] <= mem_n[692];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[691] <= 1'b0;
    end else if(1'b1) begin
      mem_q[691] <= mem_n[691];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[690] <= 1'b0;
    end else if(1'b1) begin
      mem_q[690] <= mem_n[690];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[689] <= 1'b0;
    end else if(1'b1) begin
      mem_q[689] <= mem_n[689];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[688] <= 1'b0;
    end else if(1'b1) begin
      mem_q[688] <= mem_n[688];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[687] <= 1'b0;
    end else if(1'b1) begin
      mem_q[687] <= mem_n[687];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[686] <= 1'b0;
    end else if(1'b1) begin
      mem_q[686] <= mem_n[686];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[685] <= 1'b0;
    end else if(1'b1) begin
      mem_q[685] <= mem_n[685];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[684] <= 1'b0;
    end else if(1'b1) begin
      mem_q[684] <= mem_n[684];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[683] <= 1'b0;
    end else if(1'b1) begin
      mem_q[683] <= mem_n[683];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[682] <= 1'b0;
    end else if(1'b1) begin
      mem_q[682] <= mem_n[682];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[681] <= 1'b0;
    end else if(1'b1) begin
      mem_q[681] <= mem_n[681];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[680] <= 1'b0;
    end else if(1'b1) begin
      mem_q[680] <= mem_n[680];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[679] <= 1'b0;
    end else if(1'b1) begin
      mem_q[679] <= mem_n[679];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[678] <= 1'b0;
    end else if(1'b1) begin
      mem_q[678] <= mem_n[678];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[677] <= 1'b0;
    end else if(1'b1) begin
      mem_q[677] <= mem_n[677];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[676] <= 1'b0;
    end else if(1'b1) begin
      mem_q[676] <= mem_n[676];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[675] <= 1'b0;
    end else if(1'b1) begin
      mem_q[675] <= mem_n[675];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[674] <= 1'b0;
    end else if(1'b1) begin
      mem_q[674] <= mem_n[674];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[673] <= 1'b0;
    end else if(1'b1) begin
      mem_q[673] <= mem_n[673];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[672] <= 1'b0;
    end else if(1'b1) begin
      mem_q[672] <= mem_n[672];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[671] <= 1'b0;
    end else if(1'b1) begin
      mem_q[671] <= mem_n[671];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[670] <= 1'b0;
    end else if(1'b1) begin
      mem_q[670] <= mem_n[670];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[669] <= 1'b0;
    end else if(1'b1) begin
      mem_q[669] <= mem_n[669];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[668] <= 1'b0;
    end else if(1'b1) begin
      mem_q[668] <= mem_n[668];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[667] <= 1'b0;
    end else if(1'b1) begin
      mem_q[667] <= mem_n[667];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[666] <= 1'b0;
    end else if(1'b1) begin
      mem_q[666] <= mem_n[666];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[665] <= 1'b0;
    end else if(1'b1) begin
      mem_q[665] <= mem_n[665];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[664] <= 1'b0;
    end else if(1'b1) begin
      mem_q[664] <= mem_n[664];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[663] <= 1'b0;
    end else if(1'b1) begin
      mem_q[663] <= mem_n[663];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[662] <= 1'b0;
    end else if(1'b1) begin
      mem_q[662] <= mem_n[662];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[661] <= 1'b0;
    end else if(1'b1) begin
      mem_q[661] <= mem_n[661];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[660] <= 1'b0;
    end else if(1'b1) begin
      mem_q[660] <= mem_n[660];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[659] <= 1'b0;
    end else if(1'b1) begin
      mem_q[659] <= mem_n[659];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[658] <= 1'b0;
    end else if(1'b1) begin
      mem_q[658] <= mem_n[658];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[657] <= 1'b0;
    end else if(1'b1) begin
      mem_q[657] <= mem_n[657];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[656] <= 1'b0;
    end else if(1'b1) begin
      mem_q[656] <= mem_n[656];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[655] <= 1'b0;
    end else if(1'b1) begin
      mem_q[655] <= mem_n[655];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[654] <= 1'b0;
    end else if(1'b1) begin
      mem_q[654] <= mem_n[654];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[653] <= 1'b0;
    end else if(1'b1) begin
      mem_q[653] <= mem_n[653];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[652] <= 1'b0;
    end else if(1'b1) begin
      mem_q[652] <= mem_n[652];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[651] <= 1'b0;
    end else if(1'b1) begin
      mem_q[651] <= mem_n[651];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[650] <= 1'b0;
    end else if(1'b1) begin
      mem_q[650] <= mem_n[650];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[649] <= 1'b0;
    end else if(1'b1) begin
      mem_q[649] <= mem_n[649];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[648] <= 1'b0;
    end else if(1'b1) begin
      mem_q[648] <= mem_n[648];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[647] <= 1'b0;
    end else if(1'b1) begin
      mem_q[647] <= mem_n[647];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[646] <= 1'b0;
    end else if(1'b1) begin
      mem_q[646] <= mem_n[646];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[645] <= 1'b0;
    end else if(1'b1) begin
      mem_q[645] <= mem_n[645];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[644] <= 1'b0;
    end else if(1'b1) begin
      mem_q[644] <= mem_n[644];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[643] <= 1'b0;
    end else if(1'b1) begin
      mem_q[643] <= mem_n[643];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[642] <= 1'b0;
    end else if(1'b1) begin
      mem_q[642] <= mem_n[642];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[641] <= 1'b0;
    end else if(1'b1) begin
      mem_q[641] <= mem_n[641];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[640] <= 1'b0;
    end else if(1'b1) begin
      mem_q[640] <= mem_n[640];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[639] <= 1'b0;
    end else if(1'b1) begin
      mem_q[639] <= mem_n[639];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[638] <= 1'b0;
    end else if(1'b1) begin
      mem_q[638] <= mem_n[638];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[637] <= 1'b0;
    end else if(1'b1) begin
      mem_q[637] <= mem_n[637];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[636] <= 1'b0;
    end else if(1'b1) begin
      mem_q[636] <= mem_n[636];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[635] <= 1'b0;
    end else if(1'b1) begin
      mem_q[635] <= mem_n[635];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[634] <= 1'b0;
    end else if(1'b1) begin
      mem_q[634] <= mem_n[634];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[633] <= 1'b0;
    end else if(1'b1) begin
      mem_q[633] <= mem_n[633];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[632] <= 1'b0;
    end else if(1'b1) begin
      mem_q[632] <= mem_n[632];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[631] <= 1'b0;
    end else if(1'b1) begin
      mem_q[631] <= mem_n[631];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[630] <= 1'b0;
    end else if(1'b1) begin
      mem_q[630] <= mem_n[630];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[629] <= 1'b0;
    end else if(1'b1) begin
      mem_q[629] <= mem_n[629];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[628] <= 1'b0;
    end else if(1'b1) begin
      mem_q[628] <= mem_n[628];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[627] <= 1'b0;
    end else if(1'b1) begin
      mem_q[627] <= mem_n[627];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[626] <= 1'b0;
    end else if(1'b1) begin
      mem_q[626] <= mem_n[626];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[625] <= 1'b0;
    end else if(1'b1) begin
      mem_q[625] <= mem_n[625];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[624] <= 1'b0;
    end else if(1'b1) begin
      mem_q[624] <= mem_n[624];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[623] <= 1'b0;
    end else if(1'b1) begin
      mem_q[623] <= mem_n[623];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[622] <= 1'b0;
    end else if(1'b1) begin
      mem_q[622] <= mem_n[622];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[621] <= 1'b0;
    end else if(1'b1) begin
      mem_q[621] <= mem_n[621];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[620] <= 1'b0;
    end else if(1'b1) begin
      mem_q[620] <= mem_n[620];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[619] <= 1'b0;
    end else if(1'b1) begin
      mem_q[619] <= mem_n[619];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[618] <= 1'b0;
    end else if(1'b1) begin
      mem_q[618] <= mem_n[618];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[617] <= 1'b0;
    end else if(1'b1) begin
      mem_q[617] <= mem_n[617];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[616] <= 1'b0;
    end else if(1'b1) begin
      mem_q[616] <= mem_n[616];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[615] <= 1'b0;
    end else if(1'b1) begin
      mem_q[615] <= mem_n[615];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[614] <= 1'b0;
    end else if(1'b1) begin
      mem_q[614] <= mem_n[614];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[613] <= 1'b0;
    end else if(1'b1) begin
      mem_q[613] <= mem_n[613];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[612] <= 1'b0;
    end else if(1'b1) begin
      mem_q[612] <= mem_n[612];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[611] <= 1'b0;
    end else if(1'b1) begin
      mem_q[611] <= mem_n[611];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[610] <= 1'b0;
    end else if(1'b1) begin
      mem_q[610] <= mem_n[610];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[609] <= 1'b0;
    end else if(1'b1) begin
      mem_q[609] <= mem_n[609];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[608] <= 1'b0;
    end else if(1'b1) begin
      mem_q[608] <= mem_n[608];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[607] <= 1'b0;
    end else if(1'b1) begin
      mem_q[607] <= mem_n[607];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[606] <= 1'b0;
    end else if(1'b1) begin
      mem_q[606] <= mem_n[606];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[605] <= 1'b0;
    end else if(1'b1) begin
      mem_q[605] <= mem_n[605];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[604] <= 1'b0;
    end else if(1'b1) begin
      mem_q[604] <= mem_n[604];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[603] <= 1'b0;
    end else if(1'b1) begin
      mem_q[603] <= mem_n[603];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[602] <= 1'b0;
    end else if(1'b1) begin
      mem_q[602] <= mem_n[602];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[601] <= 1'b0;
    end else if(1'b1) begin
      mem_q[601] <= mem_n[601];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[600] <= 1'b0;
    end else if(1'b1) begin
      mem_q[600] <= mem_n[600];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[599] <= 1'b0;
    end else if(1'b1) begin
      mem_q[599] <= mem_n[599];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[598] <= 1'b0;
    end else if(1'b1) begin
      mem_q[598] <= mem_n[598];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[597] <= 1'b0;
    end else if(1'b1) begin
      mem_q[597] <= mem_n[597];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[596] <= 1'b0;
    end else if(1'b1) begin
      mem_q[596] <= mem_n[596];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[595] <= 1'b0;
    end else if(1'b1) begin
      mem_q[595] <= mem_n[595];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[594] <= 1'b0;
    end else if(1'b1) begin
      mem_q[594] <= mem_n[594];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[593] <= 1'b0;
    end else if(1'b1) begin
      mem_q[593] <= mem_n[593];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[592] <= 1'b0;
    end else if(1'b1) begin
      mem_q[592] <= mem_n[592];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[591] <= 1'b0;
    end else if(1'b1) begin
      mem_q[591] <= mem_n[591];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[590] <= 1'b0;
    end else if(1'b1) begin
      mem_q[590] <= mem_n[590];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[589] <= 1'b0;
    end else if(1'b1) begin
      mem_q[589] <= mem_n[589];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[588] <= 1'b0;
    end else if(1'b1) begin
      mem_q[588] <= mem_n[588];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[587] <= 1'b0;
    end else if(1'b1) begin
      mem_q[587] <= mem_n[587];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[586] <= 1'b0;
    end else if(1'b1) begin
      mem_q[586] <= mem_n[586];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[585] <= 1'b0;
    end else if(1'b1) begin
      mem_q[585] <= mem_n[585];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[584] <= 1'b0;
    end else if(1'b1) begin
      mem_q[584] <= mem_n[584];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[583] <= 1'b0;
    end else if(1'b1) begin
      mem_q[583] <= mem_n[583];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[582] <= 1'b0;
    end else if(1'b1) begin
      mem_q[582] <= mem_n[582];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[581] <= 1'b0;
    end else if(1'b1) begin
      mem_q[581] <= mem_n[581];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[580] <= 1'b0;
    end else if(1'b1) begin
      mem_q[580] <= mem_n[580];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[579] <= 1'b0;
    end else if(1'b1) begin
      mem_q[579] <= mem_n[579];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[578] <= 1'b0;
    end else if(1'b1) begin
      mem_q[578] <= mem_n[578];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[577] <= 1'b0;
    end else if(1'b1) begin
      mem_q[577] <= mem_n[577];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[576] <= 1'b0;
    end else if(1'b1) begin
      mem_q[576] <= mem_n[576];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[575] <= 1'b0;
    end else if(1'b1) begin
      mem_q[575] <= mem_n[575];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[574] <= 1'b0;
    end else if(1'b1) begin
      mem_q[574] <= mem_n[574];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[573] <= 1'b0;
    end else if(1'b1) begin
      mem_q[573] <= mem_n[573];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[572] <= 1'b0;
    end else if(1'b1) begin
      mem_q[572] <= mem_n[572];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[571] <= 1'b0;
    end else if(1'b1) begin
      mem_q[571] <= mem_n[571];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[570] <= 1'b0;
    end else if(1'b1) begin
      mem_q[570] <= mem_n[570];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[569] <= 1'b0;
    end else if(1'b1) begin
      mem_q[569] <= mem_n[569];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[568] <= 1'b0;
    end else if(1'b1) begin
      mem_q[568] <= mem_n[568];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[567] <= 1'b0;
    end else if(1'b1) begin
      mem_q[567] <= mem_n[567];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[566] <= 1'b0;
    end else if(1'b1) begin
      mem_q[566] <= mem_n[566];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[565] <= 1'b0;
    end else if(1'b1) begin
      mem_q[565] <= mem_n[565];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[564] <= 1'b0;
    end else if(1'b1) begin
      mem_q[564] <= mem_n[564];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[563] <= 1'b0;
    end else if(1'b1) begin
      mem_q[563] <= mem_n[563];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[562] <= 1'b0;
    end else if(1'b1) begin
      mem_q[562] <= mem_n[562];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[561] <= 1'b0;
    end else if(1'b1) begin
      mem_q[561] <= mem_n[561];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[560] <= 1'b0;
    end else if(1'b1) begin
      mem_q[560] <= mem_n[560];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[559] <= 1'b0;
    end else if(1'b1) begin
      mem_q[559] <= mem_n[559];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[558] <= 1'b0;
    end else if(1'b1) begin
      mem_q[558] <= mem_n[558];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[557] <= 1'b0;
    end else if(1'b1) begin
      mem_q[557] <= mem_n[557];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[556] <= 1'b0;
    end else if(1'b1) begin
      mem_q[556] <= mem_n[556];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[555] <= 1'b0;
    end else if(1'b1) begin
      mem_q[555] <= mem_n[555];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[554] <= 1'b0;
    end else if(1'b1) begin
      mem_q[554] <= mem_n[554];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[553] <= 1'b0;
    end else if(1'b1) begin
      mem_q[553] <= mem_n[553];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[552] <= 1'b0;
    end else if(1'b1) begin
      mem_q[552] <= mem_n[552];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[551] <= 1'b0;
    end else if(1'b1) begin
      mem_q[551] <= mem_n[551];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[550] <= 1'b0;
    end else if(1'b1) begin
      mem_q[550] <= mem_n[550];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[549] <= 1'b0;
    end else if(1'b1) begin
      mem_q[549] <= mem_n[549];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[548] <= 1'b0;
    end else if(1'b1) begin
      mem_q[548] <= mem_n[548];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[547] <= 1'b0;
    end else if(1'b1) begin
      mem_q[547] <= mem_n[547];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[546] <= 1'b0;
    end else if(1'b1) begin
      mem_q[546] <= mem_n[546];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[545] <= 1'b0;
    end else if(1'b1) begin
      mem_q[545] <= mem_n[545];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[544] <= 1'b0;
    end else if(1'b1) begin
      mem_q[544] <= mem_n[544];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[543] <= 1'b0;
    end else if(1'b1) begin
      mem_q[543] <= mem_n[543];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[542] <= 1'b0;
    end else if(1'b1) begin
      mem_q[542] <= mem_n[542];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[541] <= 1'b0;
    end else if(1'b1) begin
      mem_q[541] <= mem_n[541];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[540] <= 1'b0;
    end else if(1'b1) begin
      mem_q[540] <= mem_n[540];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[539] <= 1'b0;
    end else if(1'b1) begin
      mem_q[539] <= mem_n[539];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[538] <= 1'b0;
    end else if(1'b1) begin
      mem_q[538] <= mem_n[538];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[537] <= 1'b0;
    end else if(1'b1) begin
      mem_q[537] <= mem_n[537];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[536] <= 1'b0;
    end else if(1'b1) begin
      mem_q[536] <= mem_n[536];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[535] <= 1'b0;
    end else if(1'b1) begin
      mem_q[535] <= mem_n[535];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[534] <= 1'b0;
    end else if(1'b1) begin
      mem_q[534] <= mem_n[534];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[533] <= 1'b0;
    end else if(1'b1) begin
      mem_q[533] <= mem_n[533];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[532] <= 1'b0;
    end else if(1'b1) begin
      mem_q[532] <= mem_n[532];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[531] <= 1'b0;
    end else if(1'b1) begin
      mem_q[531] <= mem_n[531];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[530] <= 1'b0;
    end else if(1'b1) begin
      mem_q[530] <= mem_n[530];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[529] <= 1'b0;
    end else if(1'b1) begin
      mem_q[529] <= mem_n[529];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[528] <= 1'b0;
    end else if(1'b1) begin
      mem_q[528] <= mem_n[528];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[527] <= 1'b0;
    end else if(1'b1) begin
      mem_q[527] <= mem_n[527];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[526] <= 1'b0;
    end else if(1'b1) begin
      mem_q[526] <= mem_n[526];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[525] <= 1'b0;
    end else if(1'b1) begin
      mem_q[525] <= mem_n[525];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[524] <= 1'b0;
    end else if(1'b1) begin
      mem_q[524] <= mem_n[524];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[523] <= 1'b0;
    end else if(1'b1) begin
      mem_q[523] <= mem_n[523];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[522] <= 1'b0;
    end else if(1'b1) begin
      mem_q[522] <= mem_n[522];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[521] <= 1'b0;
    end else if(1'b1) begin
      mem_q[521] <= mem_n[521];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[520] <= 1'b0;
    end else if(1'b1) begin
      mem_q[520] <= mem_n[520];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[519] <= 1'b0;
    end else if(1'b1) begin
      mem_q[519] <= mem_n[519];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[518] <= 1'b0;
    end else if(1'b1) begin
      mem_q[518] <= mem_n[518];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[517] <= 1'b0;
    end else if(1'b1) begin
      mem_q[517] <= mem_n[517];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[516] <= 1'b0;
    end else if(1'b1) begin
      mem_q[516] <= mem_n[516];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[515] <= 1'b0;
    end else if(1'b1) begin
      mem_q[515] <= mem_n[515];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[514] <= 1'b0;
    end else if(1'b1) begin
      mem_q[514] <= mem_n[514];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[513] <= 1'b0;
    end else if(1'b1) begin
      mem_q[513] <= mem_n[513];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[512] <= 1'b0;
    end else if(1'b1) begin
      mem_q[512] <= mem_n[512];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[511] <= 1'b0;
    end else if(1'b1) begin
      mem_q[511] <= mem_n[511];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[510] <= 1'b0;
    end else if(1'b1) begin
      mem_q[510] <= mem_n[510];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[509] <= 1'b0;
    end else if(1'b1) begin
      mem_q[509] <= mem_n[509];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[508] <= 1'b0;
    end else if(1'b1) begin
      mem_q[508] <= mem_n[508];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[507] <= 1'b0;
    end else if(1'b1) begin
      mem_q[507] <= mem_n[507];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[506] <= 1'b0;
    end else if(1'b1) begin
      mem_q[506] <= mem_n[506];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[505] <= 1'b0;
    end else if(1'b1) begin
      mem_q[505] <= mem_n[505];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[504] <= 1'b0;
    end else if(1'b1) begin
      mem_q[504] <= mem_n[504];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[503] <= 1'b0;
    end else if(1'b1) begin
      mem_q[503] <= mem_n[503];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[502] <= 1'b0;
    end else if(1'b1) begin
      mem_q[502] <= mem_n[502];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[501] <= 1'b0;
    end else if(1'b1) begin
      mem_q[501] <= mem_n[501];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[500] <= 1'b0;
    end else if(1'b1) begin
      mem_q[500] <= mem_n[500];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[499] <= 1'b0;
    end else if(1'b1) begin
      mem_q[499] <= mem_n[499];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[498] <= 1'b0;
    end else if(1'b1) begin
      mem_q[498] <= mem_n[498];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[497] <= 1'b0;
    end else if(1'b1) begin
      mem_q[497] <= mem_n[497];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[496] <= 1'b0;
    end else if(1'b1) begin
      mem_q[496] <= mem_n[496];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[495] <= 1'b0;
    end else if(1'b1) begin
      mem_q[495] <= mem_n[495];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[494] <= 1'b0;
    end else if(1'b1) begin
      mem_q[494] <= mem_n[494];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[493] <= 1'b0;
    end else if(1'b1) begin
      mem_q[493] <= mem_n[493];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[492] <= 1'b0;
    end else if(1'b1) begin
      mem_q[492] <= mem_n[492];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[491] <= 1'b0;
    end else if(1'b1) begin
      mem_q[491] <= mem_n[491];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[490] <= 1'b0;
    end else if(1'b1) begin
      mem_q[490] <= mem_n[490];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[489] <= 1'b0;
    end else if(1'b1) begin
      mem_q[489] <= mem_n[489];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[488] <= 1'b0;
    end else if(1'b1) begin
      mem_q[488] <= mem_n[488];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[487] <= 1'b0;
    end else if(1'b1) begin
      mem_q[487] <= mem_n[487];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[486] <= 1'b0;
    end else if(1'b1) begin
      mem_q[486] <= mem_n[486];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[485] <= 1'b0;
    end else if(1'b1) begin
      mem_q[485] <= mem_n[485];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[484] <= 1'b0;
    end else if(1'b1) begin
      mem_q[484] <= mem_n[484];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[483] <= 1'b0;
    end else if(1'b1) begin
      mem_q[483] <= mem_n[483];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[482] <= 1'b0;
    end else if(1'b1) begin
      mem_q[482] <= mem_n[482];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[481] <= 1'b0;
    end else if(1'b1) begin
      mem_q[481] <= mem_n[481];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[480] <= 1'b0;
    end else if(1'b1) begin
      mem_q[480] <= mem_n[480];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[479] <= 1'b0;
    end else if(1'b1) begin
      mem_q[479] <= mem_n[479];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[478] <= 1'b0;
    end else if(1'b1) begin
      mem_q[478] <= mem_n[478];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[477] <= 1'b0;
    end else if(1'b1) begin
      mem_q[477] <= mem_n[477];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[476] <= 1'b0;
    end else if(1'b1) begin
      mem_q[476] <= mem_n[476];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[475] <= 1'b0;
    end else if(1'b1) begin
      mem_q[475] <= mem_n[475];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[474] <= 1'b0;
    end else if(1'b1) begin
      mem_q[474] <= mem_n[474];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[473] <= 1'b0;
    end else if(1'b1) begin
      mem_q[473] <= mem_n[473];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[472] <= 1'b0;
    end else if(1'b1) begin
      mem_q[472] <= mem_n[472];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[471] <= 1'b0;
    end else if(1'b1) begin
      mem_q[471] <= mem_n[471];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[470] <= 1'b0;
    end else if(1'b1) begin
      mem_q[470] <= mem_n[470];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[469] <= 1'b0;
    end else if(1'b1) begin
      mem_q[469] <= mem_n[469];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[468] <= 1'b0;
    end else if(1'b1) begin
      mem_q[468] <= mem_n[468];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[467] <= 1'b0;
    end else if(1'b1) begin
      mem_q[467] <= mem_n[467];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[466] <= 1'b0;
    end else if(1'b1) begin
      mem_q[466] <= mem_n[466];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[465] <= 1'b0;
    end else if(1'b1) begin
      mem_q[465] <= mem_n[465];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[464] <= 1'b0;
    end else if(1'b1) begin
      mem_q[464] <= mem_n[464];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[463] <= 1'b0;
    end else if(1'b1) begin
      mem_q[463] <= mem_n[463];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[462] <= 1'b0;
    end else if(1'b1) begin
      mem_q[462] <= mem_n[462];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[461] <= 1'b0;
    end else if(1'b1) begin
      mem_q[461] <= mem_n[461];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[460] <= 1'b0;
    end else if(1'b1) begin
      mem_q[460] <= mem_n[460];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[459] <= 1'b0;
    end else if(1'b1) begin
      mem_q[459] <= mem_n[459];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[458] <= 1'b0;
    end else if(1'b1) begin
      mem_q[458] <= mem_n[458];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[457] <= 1'b0;
    end else if(1'b1) begin
      mem_q[457] <= mem_n[457];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[456] <= 1'b0;
    end else if(1'b1) begin
      mem_q[456] <= mem_n[456];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[455] <= 1'b0;
    end else if(1'b1) begin
      mem_q[455] <= mem_n[455];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[454] <= 1'b0;
    end else if(1'b1) begin
      mem_q[454] <= mem_n[454];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[453] <= 1'b0;
    end else if(1'b1) begin
      mem_q[453] <= mem_n[453];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[452] <= 1'b0;
    end else if(1'b1) begin
      mem_q[452] <= mem_n[452];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[451] <= 1'b0;
    end else if(1'b1) begin
      mem_q[451] <= mem_n[451];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[450] <= 1'b0;
    end else if(1'b1) begin
      mem_q[450] <= mem_n[450];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[449] <= 1'b0;
    end else if(1'b1) begin
      mem_q[449] <= mem_n[449];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[448] <= 1'b0;
    end else if(1'b1) begin
      mem_q[448] <= mem_n[448];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[447] <= 1'b0;
    end else if(1'b1) begin
      mem_q[447] <= mem_n[447];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[446] <= 1'b0;
    end else if(1'b1) begin
      mem_q[446] <= mem_n[446];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[445] <= 1'b0;
    end else if(1'b1) begin
      mem_q[445] <= mem_n[445];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[444] <= 1'b0;
    end else if(1'b1) begin
      mem_q[444] <= mem_n[444];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[443] <= 1'b0;
    end else if(1'b1) begin
      mem_q[443] <= mem_n[443];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[442] <= 1'b0;
    end else if(1'b1) begin
      mem_q[442] <= mem_n[442];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[441] <= 1'b0;
    end else if(1'b1) begin
      mem_q[441] <= mem_n[441];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[440] <= 1'b0;
    end else if(1'b1) begin
      mem_q[440] <= mem_n[440];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[439] <= 1'b0;
    end else if(1'b1) begin
      mem_q[439] <= mem_n[439];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[438] <= 1'b0;
    end else if(1'b1) begin
      mem_q[438] <= mem_n[438];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[437] <= 1'b0;
    end else if(1'b1) begin
      mem_q[437] <= mem_n[437];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[436] <= 1'b0;
    end else if(1'b1) begin
      mem_q[436] <= mem_n[436];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[435] <= 1'b0;
    end else if(1'b1) begin
      mem_q[435] <= mem_n[435];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[434] <= 1'b0;
    end else if(1'b1) begin
      mem_q[434] <= mem_n[434];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[433] <= 1'b0;
    end else if(1'b1) begin
      mem_q[433] <= mem_n[433];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[432] <= 1'b0;
    end else if(1'b1) begin
      mem_q[432] <= mem_n[432];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[431] <= 1'b0;
    end else if(1'b1) begin
      mem_q[431] <= mem_n[431];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[430] <= 1'b0;
    end else if(1'b1) begin
      mem_q[430] <= mem_n[430];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[429] <= 1'b0;
    end else if(1'b1) begin
      mem_q[429] <= mem_n[429];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[428] <= 1'b0;
    end else if(1'b1) begin
      mem_q[428] <= mem_n[428];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[427] <= 1'b0;
    end else if(1'b1) begin
      mem_q[427] <= mem_n[427];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[426] <= 1'b0;
    end else if(1'b1) begin
      mem_q[426] <= mem_n[426];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[425] <= 1'b0;
    end else if(1'b1) begin
      mem_q[425] <= mem_n[425];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[424] <= 1'b0;
    end else if(1'b1) begin
      mem_q[424] <= mem_n[424];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[423] <= 1'b0;
    end else if(1'b1) begin
      mem_q[423] <= mem_n[423];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[422] <= 1'b0;
    end else if(1'b1) begin
      mem_q[422] <= mem_n[422];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[421] <= 1'b0;
    end else if(1'b1) begin
      mem_q[421] <= mem_n[421];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[420] <= 1'b0;
    end else if(1'b1) begin
      mem_q[420] <= mem_n[420];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[419] <= 1'b0;
    end else if(1'b1) begin
      mem_q[419] <= mem_n[419];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[418] <= 1'b0;
    end else if(1'b1) begin
      mem_q[418] <= mem_n[418];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[417] <= 1'b0;
    end else if(1'b1) begin
      mem_q[417] <= mem_n[417];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[416] <= 1'b0;
    end else if(1'b1) begin
      mem_q[416] <= mem_n[416];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[415] <= 1'b0;
    end else if(1'b1) begin
      mem_q[415] <= mem_n[415];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[414] <= 1'b0;
    end else if(1'b1) begin
      mem_q[414] <= mem_n[414];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[413] <= 1'b0;
    end else if(1'b1) begin
      mem_q[413] <= mem_n[413];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[412] <= 1'b0;
    end else if(1'b1) begin
      mem_q[412] <= mem_n[412];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[411] <= 1'b0;
    end else if(1'b1) begin
      mem_q[411] <= mem_n[411];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[410] <= 1'b0;
    end else if(1'b1) begin
      mem_q[410] <= mem_n[410];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[409] <= 1'b0;
    end else if(1'b1) begin
      mem_q[409] <= mem_n[409];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[408] <= 1'b0;
    end else if(1'b1) begin
      mem_q[408] <= mem_n[408];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[407] <= 1'b0;
    end else if(1'b1) begin
      mem_q[407] <= mem_n[407];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[406] <= 1'b0;
    end else if(1'b1) begin
      mem_q[406] <= mem_n[406];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[405] <= 1'b0;
    end else if(1'b1) begin
      mem_q[405] <= mem_n[405];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[404] <= 1'b0;
    end else if(1'b1) begin
      mem_q[404] <= mem_n[404];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[403] <= 1'b0;
    end else if(1'b1) begin
      mem_q[403] <= mem_n[403];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[402] <= 1'b0;
    end else if(1'b1) begin
      mem_q[402] <= mem_n[402];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[401] <= 1'b0;
    end else if(1'b1) begin
      mem_q[401] <= mem_n[401];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[400] <= 1'b0;
    end else if(1'b1) begin
      mem_q[400] <= mem_n[400];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[399] <= 1'b0;
    end else if(1'b1) begin
      mem_q[399] <= mem_n[399];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[398] <= 1'b0;
    end else if(1'b1) begin
      mem_q[398] <= mem_n[398];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[397] <= 1'b0;
    end else if(1'b1) begin
      mem_q[397] <= mem_n[397];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[396] <= 1'b0;
    end else if(1'b1) begin
      mem_q[396] <= mem_n[396];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[395] <= 1'b0;
    end else if(1'b1) begin
      mem_q[395] <= mem_n[395];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[394] <= 1'b0;
    end else if(1'b1) begin
      mem_q[394] <= mem_n[394];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[393] <= 1'b0;
    end else if(1'b1) begin
      mem_q[393] <= mem_n[393];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[392] <= 1'b0;
    end else if(1'b1) begin
      mem_q[392] <= mem_n[392];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[391] <= 1'b0;
    end else if(1'b1) begin
      mem_q[391] <= mem_n[391];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[390] <= 1'b0;
    end else if(1'b1) begin
      mem_q[390] <= mem_n[390];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[389] <= 1'b0;
    end else if(1'b1) begin
      mem_q[389] <= mem_n[389];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[388] <= 1'b0;
    end else if(1'b1) begin
      mem_q[388] <= mem_n[388];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[387] <= 1'b0;
    end else if(1'b1) begin
      mem_q[387] <= mem_n[387];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[386] <= 1'b0;
    end else if(1'b1) begin
      mem_q[386] <= mem_n[386];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[385] <= 1'b0;
    end else if(1'b1) begin
      mem_q[385] <= mem_n[385];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[384] <= 1'b0;
    end else if(1'b1) begin
      mem_q[384] <= mem_n[384];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[383] <= 1'b0;
    end else if(1'b1) begin
      mem_q[383] <= mem_n[383];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[382] <= 1'b0;
    end else if(1'b1) begin
      mem_q[382] <= mem_n[382];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[381] <= 1'b0;
    end else if(1'b1) begin
      mem_q[381] <= mem_n[381];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[380] <= 1'b0;
    end else if(1'b1) begin
      mem_q[380] <= mem_n[380];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[379] <= 1'b0;
    end else if(1'b1) begin
      mem_q[379] <= mem_n[379];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[378] <= 1'b0;
    end else if(1'b1) begin
      mem_q[378] <= mem_n[378];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[377] <= 1'b0;
    end else if(1'b1) begin
      mem_q[377] <= mem_n[377];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[376] <= 1'b0;
    end else if(1'b1) begin
      mem_q[376] <= mem_n[376];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[375] <= 1'b0;
    end else if(1'b1) begin
      mem_q[375] <= mem_n[375];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[374] <= 1'b0;
    end else if(1'b1) begin
      mem_q[374] <= mem_n[374];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[373] <= 1'b0;
    end else if(1'b1) begin
      mem_q[373] <= mem_n[373];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[372] <= 1'b0;
    end else if(1'b1) begin
      mem_q[372] <= mem_n[372];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[371] <= 1'b0;
    end else if(1'b1) begin
      mem_q[371] <= mem_n[371];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[370] <= 1'b0;
    end else if(1'b1) begin
      mem_q[370] <= mem_n[370];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[369] <= 1'b0;
    end else if(1'b1) begin
      mem_q[369] <= mem_n[369];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[368] <= 1'b0;
    end else if(1'b1) begin
      mem_q[368] <= mem_n[368];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[367] <= 1'b0;
    end else if(1'b1) begin
      mem_q[367] <= mem_n[367];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[366] <= 1'b0;
    end else if(1'b1) begin
      mem_q[366] <= mem_n[366];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[365] <= 1'b0;
    end else if(1'b1) begin
      mem_q[365] <= mem_n[365];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[364] <= 1'b0;
    end else if(1'b1) begin
      mem_q[364] <= mem_n[364];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[363] <= 1'b0;
    end else if(1'b1) begin
      mem_q[363] <= mem_n[363];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[362] <= 1'b0;
    end else if(1'b1) begin
      mem_q[362] <= mem_n[362];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[361] <= 1'b0;
    end else if(1'b1) begin
      mem_q[361] <= mem_n[361];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[360] <= 1'b0;
    end else if(1'b1) begin
      mem_q[360] <= mem_n[360];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[359] <= 1'b0;
    end else if(1'b1) begin
      mem_q[359] <= mem_n[359];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[358] <= 1'b0;
    end else if(1'b1) begin
      mem_q[358] <= mem_n[358];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[357] <= 1'b0;
    end else if(1'b1) begin
      mem_q[357] <= mem_n[357];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[356] <= 1'b0;
    end else if(1'b1) begin
      mem_q[356] <= mem_n[356];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[355] <= 1'b0;
    end else if(1'b1) begin
      mem_q[355] <= mem_n[355];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[354] <= 1'b0;
    end else if(1'b1) begin
      mem_q[354] <= mem_n[354];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[353] <= 1'b0;
    end else if(1'b1) begin
      mem_q[353] <= mem_n[353];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[352] <= 1'b0;
    end else if(1'b1) begin
      mem_q[352] <= mem_n[352];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[351] <= 1'b0;
    end else if(1'b1) begin
      mem_q[351] <= mem_n[351];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[350] <= 1'b0;
    end else if(1'b1) begin
      mem_q[350] <= mem_n[350];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[349] <= 1'b0;
    end else if(1'b1) begin
      mem_q[349] <= mem_n[349];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[348] <= 1'b0;
    end else if(1'b1) begin
      mem_q[348] <= mem_n[348];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[347] <= 1'b0;
    end else if(1'b1) begin
      mem_q[347] <= mem_n[347];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[346] <= 1'b0;
    end else if(1'b1) begin
      mem_q[346] <= mem_n[346];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[345] <= 1'b0;
    end else if(1'b1) begin
      mem_q[345] <= mem_n[345];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[344] <= 1'b0;
    end else if(1'b1) begin
      mem_q[344] <= mem_n[344];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[343] <= 1'b0;
    end else if(1'b1) begin
      mem_q[343] <= mem_n[343];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[342] <= 1'b0;
    end else if(1'b1) begin
      mem_q[342] <= mem_n[342];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[341] <= 1'b0;
    end else if(1'b1) begin
      mem_q[341] <= mem_n[341];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[340] <= 1'b0;
    end else if(1'b1) begin
      mem_q[340] <= mem_n[340];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[339] <= 1'b0;
    end else if(1'b1) begin
      mem_q[339] <= mem_n[339];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[338] <= 1'b0;
    end else if(1'b1) begin
      mem_q[338] <= mem_n[338];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[337] <= 1'b0;
    end else if(1'b1) begin
      mem_q[337] <= mem_n[337];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[336] <= 1'b0;
    end else if(1'b1) begin
      mem_q[336] <= mem_n[336];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[335] <= 1'b0;
    end else if(1'b1) begin
      mem_q[335] <= mem_n[335];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[334] <= 1'b0;
    end else if(1'b1) begin
      mem_q[334] <= mem_n[334];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[333] <= 1'b0;
    end else if(1'b1) begin
      mem_q[333] <= mem_n[333];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[332] <= 1'b0;
    end else if(1'b1) begin
      mem_q[332] <= mem_n[332];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[331] <= 1'b0;
    end else if(1'b1) begin
      mem_q[331] <= mem_n[331];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[330] <= 1'b0;
    end else if(1'b1) begin
      mem_q[330] <= mem_n[330];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[329] <= 1'b0;
    end else if(1'b1) begin
      mem_q[329] <= mem_n[329];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[328] <= 1'b0;
    end else if(1'b1) begin
      mem_q[328] <= mem_n[328];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[327] <= 1'b0;
    end else if(1'b1) begin
      mem_q[327] <= mem_n[327];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[326] <= 1'b0;
    end else if(1'b1) begin
      mem_q[326] <= mem_n[326];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[325] <= 1'b0;
    end else if(1'b1) begin
      mem_q[325] <= mem_n[325];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[324] <= 1'b0;
    end else if(1'b1) begin
      mem_q[324] <= mem_n[324];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[323] <= 1'b0;
    end else if(1'b1) begin
      mem_q[323] <= mem_n[323];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[322] <= 1'b0;
    end else if(1'b1) begin
      mem_q[322] <= mem_n[322];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[321] <= 1'b0;
    end else if(1'b1) begin
      mem_q[321] <= mem_n[321];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[320] <= 1'b0;
    end else if(1'b1) begin
      mem_q[320] <= mem_n[320];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[319] <= 1'b0;
    end else if(1'b1) begin
      mem_q[319] <= mem_n[319];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[318] <= 1'b0;
    end else if(1'b1) begin
      mem_q[318] <= mem_n[318];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[317] <= 1'b0;
    end else if(1'b1) begin
      mem_q[317] <= mem_n[317];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[316] <= 1'b0;
    end else if(1'b1) begin
      mem_q[316] <= mem_n[316];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[315] <= 1'b0;
    end else if(1'b1) begin
      mem_q[315] <= mem_n[315];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[314] <= 1'b0;
    end else if(1'b1) begin
      mem_q[314] <= mem_n[314];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[313] <= 1'b0;
    end else if(1'b1) begin
      mem_q[313] <= mem_n[313];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[312] <= 1'b0;
    end else if(1'b1) begin
      mem_q[312] <= mem_n[312];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[311] <= 1'b0;
    end else if(1'b1) begin
      mem_q[311] <= mem_n[311];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[310] <= 1'b0;
    end else if(1'b1) begin
      mem_q[310] <= mem_n[310];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[309] <= 1'b0;
    end else if(1'b1) begin
      mem_q[309] <= mem_n[309];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[308] <= 1'b0;
    end else if(1'b1) begin
      mem_q[308] <= mem_n[308];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[307] <= 1'b0;
    end else if(1'b1) begin
      mem_q[307] <= mem_n[307];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[306] <= 1'b0;
    end else if(1'b1) begin
      mem_q[306] <= mem_n[306];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[305] <= 1'b0;
    end else if(1'b1) begin
      mem_q[305] <= mem_n[305];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[304] <= 1'b0;
    end else if(1'b1) begin
      mem_q[304] <= mem_n[304];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[303] <= 1'b0;
    end else if(1'b1) begin
      mem_q[303] <= mem_n[303];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[302] <= 1'b0;
    end else if(1'b1) begin
      mem_q[302] <= mem_n[302];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[301] <= 1'b0;
    end else if(1'b1) begin
      mem_q[301] <= mem_n[301];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[300] <= 1'b0;
    end else if(1'b1) begin
      mem_q[300] <= mem_n[300];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[299] <= 1'b0;
    end else if(1'b1) begin
      mem_q[299] <= mem_n[299];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[298] <= 1'b0;
    end else if(1'b1) begin
      mem_q[298] <= mem_n[298];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[297] <= 1'b0;
    end else if(1'b1) begin
      mem_q[297] <= mem_n[297];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[296] <= 1'b0;
    end else if(1'b1) begin
      mem_q[296] <= mem_n[296];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[295] <= 1'b0;
    end else if(1'b1) begin
      mem_q[295] <= mem_n[295];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[294] <= 1'b0;
    end else if(1'b1) begin
      mem_q[294] <= mem_n[294];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[293] <= 1'b0;
    end else if(1'b1) begin
      mem_q[293] <= mem_n[293];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[292] <= 1'b0;
    end else if(1'b1) begin
      mem_q[292] <= mem_n[292];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[291] <= 1'b0;
    end else if(1'b1) begin
      mem_q[291] <= mem_n[291];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[290] <= 1'b0;
    end else if(1'b1) begin
      mem_q[290] <= mem_n[290];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[289] <= 1'b0;
    end else if(1'b1) begin
      mem_q[289] <= mem_n[289];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[288] <= 1'b0;
    end else if(1'b1) begin
      mem_q[288] <= mem_n[288];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[287] <= 1'b0;
    end else if(1'b1) begin
      mem_q[287] <= mem_n[287];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[286] <= 1'b0;
    end else if(1'b1) begin
      mem_q[286] <= mem_n[286];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[285] <= 1'b0;
    end else if(1'b1) begin
      mem_q[285] <= mem_n[285];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[284] <= 1'b0;
    end else if(1'b1) begin
      mem_q[284] <= mem_n[284];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[283] <= 1'b0;
    end else if(1'b1) begin
      mem_q[283] <= mem_n[283];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[282] <= 1'b0;
    end else if(1'b1) begin
      mem_q[282] <= mem_n[282];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[281] <= 1'b0;
    end else if(1'b1) begin
      mem_q[281] <= mem_n[281];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[280] <= 1'b0;
    end else if(1'b1) begin
      mem_q[280] <= mem_n[280];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[279] <= 1'b0;
    end else if(1'b1) begin
      mem_q[279] <= mem_n[279];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[278] <= 1'b0;
    end else if(1'b1) begin
      mem_q[278] <= mem_n[278];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[277] <= 1'b0;
    end else if(1'b1) begin
      mem_q[277] <= mem_n[277];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[276] <= 1'b0;
    end else if(1'b1) begin
      mem_q[276] <= mem_n[276];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[275] <= 1'b0;
    end else if(1'b1) begin
      mem_q[275] <= mem_n[275];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[274] <= 1'b0;
    end else if(1'b1) begin
      mem_q[274] <= mem_n[274];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[273] <= 1'b0;
    end else if(1'b1) begin
      mem_q[273] <= mem_n[273];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[272] <= 1'b0;
    end else if(1'b1) begin
      mem_q[272] <= mem_n[272];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[271] <= 1'b0;
    end else if(1'b1) begin
      mem_q[271] <= mem_n[271];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[270] <= 1'b0;
    end else if(1'b1) begin
      mem_q[270] <= mem_n[270];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[269] <= 1'b0;
    end else if(1'b1) begin
      mem_q[269] <= mem_n[269];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[268] <= 1'b0;
    end else if(1'b1) begin
      mem_q[268] <= mem_n[268];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[267] <= 1'b0;
    end else if(1'b1) begin
      mem_q[267] <= mem_n[267];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[266] <= 1'b0;
    end else if(1'b1) begin
      mem_q[266] <= mem_n[266];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[265] <= 1'b0;
    end else if(1'b1) begin
      mem_q[265] <= mem_n[265];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[264] <= 1'b0;
    end else if(1'b1) begin
      mem_q[264] <= mem_n[264];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[263] <= 1'b0;
    end else if(1'b1) begin
      mem_q[263] <= mem_n[263];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[262] <= 1'b0;
    end else if(1'b1) begin
      mem_q[262] <= mem_n[262];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[261] <= 1'b0;
    end else if(1'b1) begin
      mem_q[261] <= mem_n[261];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[260] <= 1'b0;
    end else if(1'b1) begin
      mem_q[260] <= mem_n[260];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[259] <= 1'b0;
    end else if(1'b1) begin
      mem_q[259] <= mem_n[259];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[258] <= 1'b0;
    end else if(1'b1) begin
      mem_q[258] <= mem_n[258];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[257] <= 1'b0;
    end else if(1'b1) begin
      mem_q[257] <= mem_n[257];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[256] <= 1'b0;
    end else if(1'b1) begin
      mem_q[256] <= mem_n[256];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[255] <= 1'b0;
    end else if(1'b1) begin
      mem_q[255] <= mem_n[255];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[254] <= 1'b0;
    end else if(1'b1) begin
      mem_q[254] <= mem_n[254];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[253] <= 1'b0;
    end else if(1'b1) begin
      mem_q[253] <= mem_n[253];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[252] <= 1'b0;
    end else if(1'b1) begin
      mem_q[252] <= mem_n[252];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[251] <= 1'b0;
    end else if(1'b1) begin
      mem_q[251] <= mem_n[251];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[250] <= 1'b0;
    end else if(1'b1) begin
      mem_q[250] <= mem_n[250];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[249] <= 1'b0;
    end else if(1'b1) begin
      mem_q[249] <= mem_n[249];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[248] <= 1'b0;
    end else if(1'b1) begin
      mem_q[248] <= mem_n[248];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[247] <= 1'b0;
    end else if(1'b1) begin
      mem_q[247] <= mem_n[247];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[246] <= 1'b0;
    end else if(1'b1) begin
      mem_q[246] <= mem_n[246];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[245] <= 1'b0;
    end else if(1'b1) begin
      mem_q[245] <= mem_n[245];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[244] <= 1'b0;
    end else if(1'b1) begin
      mem_q[244] <= mem_n[244];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[243] <= 1'b0;
    end else if(1'b1) begin
      mem_q[243] <= mem_n[243];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[242] <= 1'b0;
    end else if(1'b1) begin
      mem_q[242] <= mem_n[242];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[241] <= 1'b0;
    end else if(1'b1) begin
      mem_q[241] <= mem_n[241];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[240] <= 1'b0;
    end else if(1'b1) begin
      mem_q[240] <= mem_n[240];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[239] <= 1'b0;
    end else if(1'b1) begin
      mem_q[239] <= mem_n[239];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[238] <= 1'b0;
    end else if(1'b1) begin
      mem_q[238] <= mem_n[238];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[237] <= 1'b0;
    end else if(1'b1) begin
      mem_q[237] <= mem_n[237];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[236] <= 1'b0;
    end else if(1'b1) begin
      mem_q[236] <= mem_n[236];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[235] <= 1'b0;
    end else if(1'b1) begin
      mem_q[235] <= mem_n[235];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[234] <= 1'b0;
    end else if(1'b1) begin
      mem_q[234] <= mem_n[234];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[233] <= 1'b0;
    end else if(1'b1) begin
      mem_q[233] <= mem_n[233];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[232] <= 1'b0;
    end else if(1'b1) begin
      mem_q[232] <= mem_n[232];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[231] <= 1'b0;
    end else if(1'b1) begin
      mem_q[231] <= mem_n[231];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[230] <= 1'b0;
    end else if(1'b1) begin
      mem_q[230] <= mem_n[230];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[229] <= 1'b0;
    end else if(1'b1) begin
      mem_q[229] <= mem_n[229];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[228] <= 1'b0;
    end else if(1'b1) begin
      mem_q[228] <= mem_n[228];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[227] <= 1'b0;
    end else if(1'b1) begin
      mem_q[227] <= mem_n[227];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[226] <= 1'b0;
    end else if(1'b1) begin
      mem_q[226] <= mem_n[226];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[225] <= 1'b0;
    end else if(1'b1) begin
      mem_q[225] <= mem_n[225];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[224] <= 1'b0;
    end else if(1'b1) begin
      mem_q[224] <= mem_n[224];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[223] <= 1'b0;
    end else if(1'b1) begin
      mem_q[223] <= mem_n[223];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[222] <= 1'b0;
    end else if(1'b1) begin
      mem_q[222] <= mem_n[222];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[221] <= 1'b0;
    end else if(1'b1) begin
      mem_q[221] <= mem_n[221];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[220] <= 1'b0;
    end else if(1'b1) begin
      mem_q[220] <= mem_n[220];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[219] <= 1'b0;
    end else if(1'b1) begin
      mem_q[219] <= mem_n[219];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[218] <= 1'b0;
    end else if(1'b1) begin
      mem_q[218] <= mem_n[218];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[217] <= 1'b0;
    end else if(1'b1) begin
      mem_q[217] <= mem_n[217];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[216] <= 1'b0;
    end else if(1'b1) begin
      mem_q[216] <= mem_n[216];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[215] <= 1'b0;
    end else if(1'b1) begin
      mem_q[215] <= mem_n[215];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[214] <= 1'b0;
    end else if(1'b1) begin
      mem_q[214] <= mem_n[214];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[213] <= 1'b0;
    end else if(1'b1) begin
      mem_q[213] <= mem_n[213];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[212] <= 1'b0;
    end else if(1'b1) begin
      mem_q[212] <= mem_n[212];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[211] <= 1'b0;
    end else if(1'b1) begin
      mem_q[211] <= mem_n[211];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[210] <= 1'b0;
    end else if(1'b1) begin
      mem_q[210] <= mem_n[210];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[209] <= 1'b0;
    end else if(1'b1) begin
      mem_q[209] <= mem_n[209];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[208] <= 1'b0;
    end else if(1'b1) begin
      mem_q[208] <= mem_n[208];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[207] <= 1'b0;
    end else if(1'b1) begin
      mem_q[207] <= mem_n[207];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[206] <= 1'b0;
    end else if(1'b1) begin
      mem_q[206] <= mem_n[206];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[205] <= 1'b0;
    end else if(1'b1) begin
      mem_q[205] <= mem_n[205];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[204] <= 1'b0;
    end else if(1'b1) begin
      mem_q[204] <= mem_n[204];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[203] <= 1'b0;
    end else if(1'b1) begin
      mem_q[203] <= mem_n[203];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[202] <= 1'b0;
    end else if(1'b1) begin
      mem_q[202] <= mem_n[202];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[201] <= 1'b0;
    end else if(1'b1) begin
      mem_q[201] <= mem_n[201];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[200] <= 1'b0;
    end else if(1'b1) begin
      mem_q[200] <= mem_n[200];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[199] <= 1'b0;
    end else if(1'b1) begin
      mem_q[199] <= mem_n[199];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[198] <= 1'b0;
    end else if(1'b1) begin
      mem_q[198] <= mem_n[198];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[197] <= 1'b0;
    end else if(1'b1) begin
      mem_q[197] <= mem_n[197];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[196] <= 1'b0;
    end else if(1'b1) begin
      mem_q[196] <= mem_n[196];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[195] <= 1'b0;
    end else if(1'b1) begin
      mem_q[195] <= mem_n[195];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[194] <= 1'b0;
    end else if(1'b1) begin
      mem_q[194] <= mem_n[194];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[193] <= 1'b0;
    end else if(1'b1) begin
      mem_q[193] <= mem_n[193];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[192] <= 1'b0;
    end else if(1'b1) begin
      mem_q[192] <= mem_n[192];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[191] <= 1'b0;
    end else if(1'b1) begin
      mem_q[191] <= mem_n[191];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[190] <= 1'b0;
    end else if(1'b1) begin
      mem_q[190] <= mem_n[190];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[189] <= 1'b0;
    end else if(1'b1) begin
      mem_q[189] <= mem_n[189];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[188] <= 1'b0;
    end else if(1'b1) begin
      mem_q[188] <= mem_n[188];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[187] <= 1'b0;
    end else if(1'b1) begin
      mem_q[187] <= mem_n[187];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[186] <= 1'b0;
    end else if(1'b1) begin
      mem_q[186] <= mem_n[186];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[185] <= 1'b0;
    end else if(1'b1) begin
      mem_q[185] <= mem_n[185];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[184] <= 1'b0;
    end else if(1'b1) begin
      mem_q[184] <= mem_n[184];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[183] <= 1'b0;
    end else if(1'b1) begin
      mem_q[183] <= mem_n[183];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[182] <= 1'b0;
    end else if(1'b1) begin
      mem_q[182] <= mem_n[182];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[181] <= 1'b0;
    end else if(1'b1) begin
      mem_q[181] <= mem_n[181];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[180] <= 1'b0;
    end else if(1'b1) begin
      mem_q[180] <= mem_n[180];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[179] <= 1'b0;
    end else if(1'b1) begin
      mem_q[179] <= mem_n[179];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[178] <= 1'b0;
    end else if(1'b1) begin
      mem_q[178] <= mem_n[178];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[177] <= 1'b0;
    end else if(1'b1) begin
      mem_q[177] <= mem_n[177];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[176] <= 1'b0;
    end else if(1'b1) begin
      mem_q[176] <= mem_n[176];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[175] <= 1'b0;
    end else if(1'b1) begin
      mem_q[175] <= mem_n[175];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[174] <= 1'b0;
    end else if(1'b1) begin
      mem_q[174] <= mem_n[174];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[173] <= 1'b0;
    end else if(1'b1) begin
      mem_q[173] <= mem_n[173];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[172] <= 1'b0;
    end else if(1'b1) begin
      mem_q[172] <= mem_n[172];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[171] <= 1'b0;
    end else if(1'b1) begin
      mem_q[171] <= mem_n[171];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[170] <= 1'b0;
    end else if(1'b1) begin
      mem_q[170] <= mem_n[170];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[169] <= 1'b0;
    end else if(1'b1) begin
      mem_q[169] <= mem_n[169];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[168] <= 1'b0;
    end else if(1'b1) begin
      mem_q[168] <= mem_n[168];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[167] <= 1'b0;
    end else if(1'b1) begin
      mem_q[167] <= mem_n[167];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[166] <= 1'b0;
    end else if(1'b1) begin
      mem_q[166] <= mem_n[166];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[165] <= 1'b0;
    end else if(1'b1) begin
      mem_q[165] <= mem_n[165];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[164] <= 1'b0;
    end else if(1'b1) begin
      mem_q[164] <= mem_n[164];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[163] <= 1'b0;
    end else if(1'b1) begin
      mem_q[163] <= mem_n[163];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[162] <= 1'b0;
    end else if(1'b1) begin
      mem_q[162] <= mem_n[162];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[161] <= 1'b0;
    end else if(1'b1) begin
      mem_q[161] <= mem_n[161];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[160] <= 1'b0;
    end else if(1'b1) begin
      mem_q[160] <= mem_n[160];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[159] <= 1'b0;
    end else if(1'b1) begin
      mem_q[159] <= mem_n[159];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[158] <= 1'b0;
    end else if(1'b1) begin
      mem_q[158] <= mem_n[158];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[157] <= 1'b0;
    end else if(1'b1) begin
      mem_q[157] <= mem_n[157];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[156] <= 1'b0;
    end else if(1'b1) begin
      mem_q[156] <= mem_n[156];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[155] <= 1'b0;
    end else if(1'b1) begin
      mem_q[155] <= mem_n[155];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[154] <= 1'b0;
    end else if(1'b1) begin
      mem_q[154] <= mem_n[154];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[153] <= 1'b0;
    end else if(1'b1) begin
      mem_q[153] <= mem_n[153];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[152] <= 1'b0;
    end else if(1'b1) begin
      mem_q[152] <= mem_n[152];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[151] <= 1'b0;
    end else if(1'b1) begin
      mem_q[151] <= mem_n[151];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[150] <= 1'b0;
    end else if(1'b1) begin
      mem_q[150] <= mem_n[150];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[149] <= 1'b0;
    end else if(1'b1) begin
      mem_q[149] <= mem_n[149];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[148] <= 1'b0;
    end else if(1'b1) begin
      mem_q[148] <= mem_n[148];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[147] <= 1'b0;
    end else if(1'b1) begin
      mem_q[147] <= mem_n[147];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[146] <= 1'b0;
    end else if(1'b1) begin
      mem_q[146] <= mem_n[146];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[145] <= 1'b0;
    end else if(1'b1) begin
      mem_q[145] <= mem_n[145];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[144] <= 1'b0;
    end else if(1'b1) begin
      mem_q[144] <= mem_n[144];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[143] <= 1'b0;
    end else if(1'b1) begin
      mem_q[143] <= mem_n[143];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[142] <= 1'b0;
    end else if(1'b1) begin
      mem_q[142] <= mem_n[142];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[141] <= 1'b0;
    end else if(1'b1) begin
      mem_q[141] <= mem_n[141];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[140] <= 1'b0;
    end else if(1'b1) begin
      mem_q[140] <= mem_n[140];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[139] <= 1'b0;
    end else if(1'b1) begin
      mem_q[139] <= mem_n[139];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[138] <= 1'b0;
    end else if(1'b1) begin
      mem_q[138] <= mem_n[138];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[137] <= 1'b0;
    end else if(1'b1) begin
      mem_q[137] <= mem_n[137];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[136] <= 1'b0;
    end else if(1'b1) begin
      mem_q[136] <= mem_n[136];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[135] <= 1'b0;
    end else if(1'b1) begin
      mem_q[135] <= mem_n[135];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[134] <= 1'b0;
    end else if(1'b1) begin
      mem_q[134] <= mem_n[134];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[133] <= 1'b0;
    end else if(1'b1) begin
      mem_q[133] <= mem_n[133];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[132] <= 1'b0;
    end else if(1'b1) begin
      mem_q[132] <= mem_n[132];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[131] <= 1'b0;
    end else if(1'b1) begin
      mem_q[131] <= mem_n[131];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[130] <= 1'b0;
    end else if(1'b1) begin
      mem_q[130] <= mem_n[130];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[129] <= 1'b0;
    end else if(1'b1) begin
      mem_q[129] <= mem_n[129];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[128] <= 1'b0;
    end else if(1'b1) begin
      mem_q[128] <= mem_n[128];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[127] <= 1'b0;
    end else if(1'b1) begin
      mem_q[127] <= mem_n[127];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[126] <= 1'b0;
    end else if(1'b1) begin
      mem_q[126] <= mem_n[126];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[125] <= 1'b0;
    end else if(1'b1) begin
      mem_q[125] <= mem_n[125];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[124] <= 1'b0;
    end else if(1'b1) begin
      mem_q[124] <= mem_n[124];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[123] <= 1'b0;
    end else if(1'b1) begin
      mem_q[123] <= mem_n[123];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[122] <= 1'b0;
    end else if(1'b1) begin
      mem_q[122] <= mem_n[122];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[121] <= 1'b0;
    end else if(1'b1) begin
      mem_q[121] <= mem_n[121];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[120] <= 1'b0;
    end else if(1'b1) begin
      mem_q[120] <= mem_n[120];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[119] <= 1'b0;
    end else if(1'b1) begin
      mem_q[119] <= mem_n[119];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[118] <= 1'b0;
    end else if(1'b1) begin
      mem_q[118] <= mem_n[118];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[117] <= 1'b0;
    end else if(1'b1) begin
      mem_q[117] <= mem_n[117];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[116] <= 1'b0;
    end else if(1'b1) begin
      mem_q[116] <= mem_n[116];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[115] <= 1'b0;
    end else if(1'b1) begin
      mem_q[115] <= mem_n[115];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[114] <= 1'b0;
    end else if(1'b1) begin
      mem_q[114] <= mem_n[114];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[113] <= 1'b0;
    end else if(1'b1) begin
      mem_q[113] <= mem_n[113];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[112] <= 1'b0;
    end else if(1'b1) begin
      mem_q[112] <= mem_n[112];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[111] <= 1'b0;
    end else if(1'b1) begin
      mem_q[111] <= mem_n[111];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[110] <= 1'b0;
    end else if(1'b1) begin
      mem_q[110] <= mem_n[110];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[109] <= 1'b0;
    end else if(1'b1) begin
      mem_q[109] <= mem_n[109];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[108] <= 1'b0;
    end else if(1'b1) begin
      mem_q[108] <= mem_n[108];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[107] <= 1'b0;
    end else if(1'b1) begin
      mem_q[107] <= mem_n[107];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[106] <= 1'b0;
    end else if(1'b1) begin
      mem_q[106] <= mem_n[106];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[105] <= 1'b0;
    end else if(1'b1) begin
      mem_q[105] <= mem_n[105];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[104] <= 1'b0;
    end else if(1'b1) begin
      mem_q[104] <= mem_n[104];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[103] <= 1'b0;
    end else if(1'b1) begin
      mem_q[103] <= mem_n[103];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[102] <= 1'b0;
    end else if(1'b1) begin
      mem_q[102] <= mem_n[102];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[101] <= 1'b0;
    end else if(1'b1) begin
      mem_q[101] <= mem_n[101];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[100] <= 1'b0;
    end else if(1'b1) begin
      mem_q[100] <= mem_n[100];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[99] <= 1'b0;
    end else if(1'b1) begin
      mem_q[99] <= mem_n[99];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[98] <= 1'b0;
    end else if(1'b1) begin
      mem_q[98] <= mem_n[98];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[97] <= 1'b0;
    end else if(1'b1) begin
      mem_q[97] <= mem_n[97];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[96] <= 1'b0;
    end else if(1'b1) begin
      mem_q[96] <= mem_n[96];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[95] <= 1'b0;
    end else if(1'b1) begin
      mem_q[95] <= mem_n[95];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[94] <= 1'b0;
    end else if(1'b1) begin
      mem_q[94] <= mem_n[94];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[93] <= 1'b0;
    end else if(1'b1) begin
      mem_q[93] <= mem_n[93];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[92] <= 1'b0;
    end else if(1'b1) begin
      mem_q[92] <= mem_n[92];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[91] <= 1'b0;
    end else if(1'b1) begin
      mem_q[91] <= mem_n[91];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[90] <= 1'b0;
    end else if(1'b1) begin
      mem_q[90] <= mem_n[90];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[89] <= 1'b0;
    end else if(1'b1) begin
      mem_q[89] <= mem_n[89];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[88] <= 1'b0;
    end else if(1'b1) begin
      mem_q[88] <= mem_n[88];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[87] <= 1'b0;
    end else if(1'b1) begin
      mem_q[87] <= mem_n[87];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[86] <= 1'b0;
    end else if(1'b1) begin
      mem_q[86] <= mem_n[86];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[85] <= 1'b0;
    end else if(1'b1) begin
      mem_q[85] <= mem_n[85];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[84] <= 1'b0;
    end else if(1'b1) begin
      mem_q[84] <= mem_n[84];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[83] <= 1'b0;
    end else if(1'b1) begin
      mem_q[83] <= mem_n[83];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[82] <= 1'b0;
    end else if(1'b1) begin
      mem_q[82] <= mem_n[82];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[81] <= 1'b0;
    end else if(1'b1) begin
      mem_q[81] <= mem_n[81];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[80] <= 1'b0;
    end else if(1'b1) begin
      mem_q[80] <= mem_n[80];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[79] <= 1'b0;
    end else if(1'b1) begin
      mem_q[79] <= mem_n[79];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[78] <= 1'b0;
    end else if(1'b1) begin
      mem_q[78] <= mem_n[78];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[77] <= 1'b0;
    end else if(1'b1) begin
      mem_q[77] <= mem_n[77];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[76] <= 1'b0;
    end else if(1'b1) begin
      mem_q[76] <= mem_n[76];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[75] <= 1'b0;
    end else if(1'b1) begin
      mem_q[75] <= mem_n[75];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[74] <= 1'b0;
    end else if(1'b1) begin
      mem_q[74] <= mem_n[74];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[73] <= 1'b0;
    end else if(1'b1) begin
      mem_q[73] <= mem_n[73];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[72] <= 1'b0;
    end else if(1'b1) begin
      mem_q[72] <= mem_n[72];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[71] <= 1'b0;
    end else if(1'b1) begin
      mem_q[71] <= mem_n[71];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[70] <= 1'b0;
    end else if(1'b1) begin
      mem_q[70] <= mem_n[70];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[69] <= 1'b0;
    end else if(1'b1) begin
      mem_q[69] <= mem_n[69];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[68] <= 1'b0;
    end else if(1'b1) begin
      mem_q[68] <= mem_n[68];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[67] <= 1'b0;
    end else if(1'b1) begin
      mem_q[67] <= mem_n[67];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[66] <= 1'b0;
    end else if(1'b1) begin
      mem_q[66] <= mem_n[66];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[65] <= 1'b0;
    end else if(1'b1) begin
      mem_q[65] <= mem_n[65];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[64] <= 1'b0;
    end else if(1'b1) begin
      mem_q[64] <= mem_n[64];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[63] <= 1'b0;
    end else if(1'b1) begin
      mem_q[63] <= mem_n[63];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[62] <= 1'b0;
    end else if(1'b1) begin
      mem_q[62] <= mem_n[62];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[61] <= 1'b0;
    end else if(1'b1) begin
      mem_q[61] <= mem_n[61];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[60] <= 1'b0;
    end else if(1'b1) begin
      mem_q[60] <= mem_n[60];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[59] <= 1'b0;
    end else if(1'b1) begin
      mem_q[59] <= mem_n[59];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[58] <= 1'b0;
    end else if(1'b1) begin
      mem_q[58] <= mem_n[58];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[57] <= 1'b0;
    end else if(1'b1) begin
      mem_q[57] <= mem_n[57];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[56] <= 1'b0;
    end else if(1'b1) begin
      mem_q[56] <= mem_n[56];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[55] <= 1'b0;
    end else if(1'b1) begin
      mem_q[55] <= mem_n[55];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[54] <= 1'b0;
    end else if(1'b1) begin
      mem_q[54] <= mem_n[54];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[53] <= 1'b0;
    end else if(1'b1) begin
      mem_q[53] <= mem_n[53];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[52] <= 1'b0;
    end else if(1'b1) begin
      mem_q[52] <= mem_n[52];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[51] <= 1'b0;
    end else if(1'b1) begin
      mem_q[51] <= mem_n[51];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[50] <= 1'b0;
    end else if(1'b1) begin
      mem_q[50] <= mem_n[50];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[49] <= 1'b0;
    end else if(1'b1) begin
      mem_q[49] <= mem_n[49];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[48] <= 1'b0;
    end else if(1'b1) begin
      mem_q[48] <= mem_n[48];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[47] <= 1'b0;
    end else if(1'b1) begin
      mem_q[47] <= mem_n[47];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[46] <= 1'b0;
    end else if(1'b1) begin
      mem_q[46] <= mem_n[46];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[45] <= 1'b0;
    end else if(1'b1) begin
      mem_q[45] <= mem_n[45];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[44] <= 1'b0;
    end else if(1'b1) begin
      mem_q[44] <= mem_n[44];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[43] <= 1'b0;
    end else if(1'b1) begin
      mem_q[43] <= mem_n[43];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[42] <= 1'b0;
    end else if(1'b1) begin
      mem_q[42] <= mem_n[42];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[41] <= 1'b0;
    end else if(1'b1) begin
      mem_q[41] <= mem_n[41];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[40] <= 1'b0;
    end else if(1'b1) begin
      mem_q[40] <= mem_n[40];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[39] <= 1'b0;
    end else if(1'b1) begin
      mem_q[39] <= mem_n[39];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[38] <= 1'b0;
    end else if(1'b1) begin
      mem_q[38] <= mem_n[38];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[37] <= 1'b0;
    end else if(1'b1) begin
      mem_q[37] <= mem_n[37];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[36] <= 1'b0;
    end else if(1'b1) begin
      mem_q[36] <= mem_n[36];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[35] <= 1'b0;
    end else if(1'b1) begin
      mem_q[35] <= mem_n[35];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[34] <= 1'b0;
    end else if(1'b1) begin
      mem_q[34] <= mem_n[34];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[33] <= 1'b0;
    end else if(1'b1) begin
      mem_q[33] <= mem_n[33];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[32] <= 1'b0;
    end else if(1'b1) begin
      mem_q[32] <= mem_n[32];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[31] <= 1'b0;
    end else if(1'b1) begin
      mem_q[31] <= mem_n[31];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[30] <= 1'b0;
    end else if(1'b1) begin
      mem_q[30] <= mem_n[30];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[29] <= 1'b0;
    end else if(1'b1) begin
      mem_q[29] <= mem_n[29];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[28] <= 1'b0;
    end else if(1'b1) begin
      mem_q[28] <= mem_n[28];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[27] <= 1'b0;
    end else if(1'b1) begin
      mem_q[27] <= mem_n[27];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[26] <= 1'b0;
    end else if(1'b1) begin
      mem_q[26] <= mem_n[26];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[25] <= 1'b0;
    end else if(1'b1) begin
      mem_q[25] <= mem_n[25];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[24] <= 1'b0;
    end else if(1'b1) begin
      mem_q[24] <= mem_n[24];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[23] <= 1'b0;
    end else if(1'b1) begin
      mem_q[23] <= mem_n[23];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[22] <= 1'b0;
    end else if(1'b1) begin
      mem_q[22] <= mem_n[22];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[21] <= 1'b0;
    end else if(1'b1) begin
      mem_q[21] <= mem_n[21];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[20] <= 1'b0;
    end else if(1'b1) begin
      mem_q[20] <= mem_n[20];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[19] <= 1'b0;
    end else if(1'b1) begin
      mem_q[19] <= mem_n[19];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[18] <= 1'b0;
    end else if(1'b1) begin
      mem_q[18] <= mem_n[18];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[17] <= 1'b0;
    end else if(1'b1) begin
      mem_q[17] <= mem_n[17];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[16] <= 1'b0;
    end else if(1'b1) begin
      mem_q[16] <= mem_n[16];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[15] <= 1'b0;
    end else if(1'b1) begin
      mem_q[15] <= mem_n[15];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[14] <= 1'b0;
    end else if(1'b1) begin
      mem_q[14] <= mem_n[14];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[13] <= 1'b0;
    end else if(1'b1) begin
      mem_q[13] <= mem_n[13];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[12] <= 1'b0;
    end else if(1'b1) begin
      mem_q[12] <= mem_n[12];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[11] <= 1'b0;
    end else if(1'b1) begin
      mem_q[11] <= mem_n[11];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[10] <= 1'b0;
    end else if(1'b1) begin
      mem_q[10] <= mem_n[10];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[9] <= 1'b0;
    end else if(1'b1) begin
      mem_q[9] <= mem_n[9];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[8] <= 1'b0;
    end else if(1'b1) begin
      mem_q[8] <= mem_n[8];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[7] <= 1'b0;
    end else if(1'b1) begin
      mem_q[7] <= mem_n[7];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[6] <= 1'b0;
    end else if(1'b1) begin
      mem_q[6] <= mem_n[6];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[5] <= 1'b0;
    end else if(1'b1) begin
      mem_q[5] <= mem_n[5];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[4] <= 1'b0;
    end else if(1'b1) begin
      mem_q[4] <= mem_n[4];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[3] <= 1'b0;
    end else if(1'b1) begin
      mem_q[3] <= mem_n[3];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[2] <= 1'b0;
    end else if(1'b1) begin
      mem_q[2] <= mem_n[2];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[1] <= 1'b0;
    end else if(1'b1) begin
      mem_q[1] <= mem_n[1];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      mem_q[0] <= 1'b0;
    end else if(1'b1) begin
      mem_q[0] <= mem_n[0];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      issue_cnt_q[2] <= 1'b0;
    end else if(1'b1) begin
      issue_cnt_q[2] <= issue_cnt_n[2];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      issue_cnt_q[1] <= 1'b0;
    end else if(1'b1) begin
      issue_cnt_q[1] <= issue_cnt_n[1];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      issue_cnt_q[0] <= 1'b0;
    end else if(1'b1) begin
      issue_cnt_q[0] <= issue_cnt_n[0];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      commit_pointer_q[2] <= 1'b0;
    end else if(1'b1) begin
      commit_pointer_q[2] <= commit_pointer_n[2];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      commit_pointer_q[1] <= 1'b0;
    end else if(1'b1) begin
      commit_pointer_q[1] <= commit_pointer_n[1];
    end 
  end


  always @(posedge clk_i or posedge N38659) begin
    if(N38659) begin
      commit_pointer_q[0] <= 1'b0;
    end else if(1'b1) begin
      commit_pointer_q[0] <= commit_pointer_n[0];
    end 
  end

  assign N38662 = rs1_i[4] | rs1_i[5];
  assign N38663 = rs1_i[3] | N38662;
  assign N38664 = rs1_i[2] | N38663;
  assign N38665 = rs1_i[1] | N38664;
  assign N38666 = rs1_i[0] | N38665;
  assign N38667 = ~N38666;
  assign N38668 = rs2_i[4] | rs2_i[5];
  assign N38669 = rs2_i[3] | N38668;
  assign N38670 = rs2_i[2] | N38669;
  assign N38671 = rs2_i[1] | N38670;
  assign N38672 = rs2_i[0] | N38671;
  assign N38673 = ~N38672;
  assign N38674 = issue_cnt_q[1] & issue_cnt_q[2];
  assign sb_full_o = issue_cnt_q[0] & N38674;
  assign { N866, N865, N864 } = commit_pointer_q + 1'b1;
  assign { N28857, N28856, N28855 } = commit_pointer_q + 1'b1;
  assign { N28884, N28883, N28882 } = commit_pointer_q + 1'b1;
  assign { N28830, N28829, N28828 } = commit_pointer_q + 1'b1;
  assign { N28911, N28910, N28909 } = { N28852, N28851, N28850 } + 1'b1;
  assign { N887, N886, N885 } = issue_cnt_q + 1'b1;
  assign { N3810, N3809, N3808 } = issue_instr_o[297:295] + 1'b1;
  assign { N28833, N28832, N28831 } = { N3813, N3812, N3811 } - commit_ack_i[0];
  assign { N28914, N28913, N28912 } = { N28833, N28832, N28831 } - commit_ack_i[1];
  assign N38676 = issue_instr_o[295] & issue_instr_o[296];
  assign N895 = N38676 & issue_instr_o[297];
  assign N38677 = N0 & issue_instr_o[296];
  assign N0 = ~issue_instr_o[295];
  assign N894 = N38677 & issue_instr_o[297];
  assign N38678 = issue_instr_o[295] & N1;
  assign N1 = ~issue_instr_o[296];
  assign N893 = N38678 & issue_instr_o[297];
  assign N38679 = N2 & N3;
  assign N2 = ~issue_instr_o[295];
  assign N3 = ~issue_instr_o[296];
  assign N892 = N38679 & issue_instr_o[297];
  assign N38680 = issue_instr_o[295] & issue_instr_o[296];
  assign N891 = N38680 & N4;
  assign N4 = ~issue_instr_o[297];
  assign N38681 = N5 & issue_instr_o[296];
  assign N5 = ~issue_instr_o[295];
  assign N890 = N38681 & N6;
  assign N6 = ~issue_instr_o[297];
  assign N38682 = issue_instr_o[295] & N7;
  assign N7 = ~issue_instr_o[296];
  assign N889 = N38682 & N8;
  assign N8 = ~issue_instr_o[297];
  assign N38683 = N9 & N10;
  assign N9 = ~issue_instr_o[295];
  assign N10 = ~issue_instr_o[296];
  assign N888 = N38683 & N11;
  assign N11 = ~issue_instr_o[297];
  assign N38684 = trans_id_i[0] & trans_id_i[1];
  assign N5919 = N38684 & trans_id_i[2];
  assign N38685 = N12 & trans_id_i[1];
  assign N12 = ~trans_id_i[0];
  assign N5918 = N38685 & trans_id_i[2];
  assign N38686 = trans_id_i[0] & N13;
  assign N13 = ~trans_id_i[1];
  assign N5917 = N38686 & trans_id_i[2];
  assign N38687 = N14 & N15;
  assign N14 = ~trans_id_i[0];
  assign N15 = ~trans_id_i[1];
  assign N5916 = N38687 & trans_id_i[2];
  assign N5915 = N38684 & N16;
  assign N16 = ~trans_id_i[2];
  assign N5914 = N38685 & N17;
  assign N17 = ~trans_id_i[2];
  assign N5913 = N38686 & N18;
  assign N18 = ~trans_id_i[2];
  assign N5912 = N38687 & N19;
  assign N19 = ~trans_id_i[2];
  assign N38688 = trans_id_i[3] & trans_id_i[4];
  assign N12154 = N38688 & trans_id_i[5];
  assign N38689 = N20 & trans_id_i[4];
  assign N20 = ~trans_id_i[3];
  assign N12153 = N38689 & trans_id_i[5];
  assign N38690 = trans_id_i[3] & N21;
  assign N21 = ~trans_id_i[4];
  assign N12152 = N38690 & trans_id_i[5];
  assign N38691 = N22 & N23;
  assign N22 = ~trans_id_i[3];
  assign N23 = ~trans_id_i[4];
  assign N12151 = N38691 & trans_id_i[5];
  assign N12150 = N38688 & N24;
  assign N24 = ~trans_id_i[5];
  assign N12149 = N38689 & N25;
  assign N25 = ~trans_id_i[5];
  assign N12148 = N38690 & N26;
  assign N26 = ~trans_id_i[5];
  assign N12147 = N38691 & N27;
  assign N27 = ~trans_id_i[5];
  assign N38692 = trans_id_i[6] & trans_id_i[7];
  assign N18389 = N38692 & trans_id_i[8];
  assign N38693 = N28 & trans_id_i[7];
  assign N28 = ~trans_id_i[6];
  assign N18388 = N38693 & trans_id_i[8];
  assign N38694 = trans_id_i[6] & N29;
  assign N29 = ~trans_id_i[7];
  assign N18387 = N38694 & trans_id_i[8];
  assign N38695 = N30 & N31;
  assign N30 = ~trans_id_i[6];
  assign N31 = ~trans_id_i[7];
  assign N18386 = N38695 & trans_id_i[8];
  assign N18385 = N38692 & N32;
  assign N32 = ~trans_id_i[8];
  assign N18384 = N38693 & N33;
  assign N33 = ~trans_id_i[8];
  assign N18383 = N38694 & N34;
  assign N34 = ~trans_id_i[8];
  assign N18382 = N38695 & N35;
  assign N35 = ~trans_id_i[8];
  assign N38696 = trans_id_i[9] & trans_id_i[10];
  assign N24624 = N38696 & trans_id_i[11];
  assign N38697 = N36 & trans_id_i[10];
  assign N36 = ~trans_id_i[9];
  assign N24623 = N38697 & trans_id_i[11];
  assign N38698 = trans_id_i[9] & N37;
  assign N37 = ~trans_id_i[10];
  assign N24622 = N38698 & trans_id_i[11];
  assign N38699 = N38 & N39;
  assign N38 = ~trans_id_i[9];
  assign N39 = ~trans_id_i[10];
  assign N24621 = N38699 & trans_id_i[11];
  assign N24620 = N38696 & N40;
  assign N40 = ~trans_id_i[11];
  assign N24619 = N38697 & N41;
  assign N41 = ~trans_id_i[11];
  assign N24618 = N38698 & N42;
  assign N42 = ~trans_id_i[11];
  assign N24617 = N38699 & N43;
  assign N43 = ~trans_id_i[11];
  assign N38700 = commit_pointer_q[0] & commit_pointer_q[1];
  assign N28787 = N38700 & commit_pointer_q[2];
  assign N38701 = N44 & commit_pointer_q[1];
  assign N44 = ~commit_pointer_q[0];
  assign N28786 = N38701 & commit_pointer_q[2];
  assign N38702 = commit_pointer_q[0] & N45;
  assign N45 = ~commit_pointer_q[1];
  assign N28785 = N38702 & commit_pointer_q[2];
  assign N38703 = N46 & N47;
  assign N46 = ~commit_pointer_q[0];
  assign N47 = ~commit_pointer_q[1];
  assign N28784 = N38703 & commit_pointer_q[2];
  assign N38704 = commit_pointer_q[0] & commit_pointer_q[1];
  assign N28783 = N38704 & N48;
  assign N48 = ~commit_pointer_q[2];
  assign N38705 = N49 & commit_pointer_q[1];
  assign N49 = ~commit_pointer_q[0];
  assign N28782 = N38705 & N50;
  assign N50 = ~commit_pointer_q[2];
  assign N38706 = commit_pointer_q[0] & N51;
  assign N51 = ~commit_pointer_q[1];
  assign N28781 = N38706 & N52;
  assign N52 = ~commit_pointer_q[2];
  assign N38707 = N53 & N54;
  assign N53 = ~commit_pointer_q[0];
  assign N54 = ~commit_pointer_q[1];
  assign N28780 = N38707 & N55;
  assign N55 = ~commit_pointer_q[2];
  assign N38708 = commit_pointer_q[0] & commit_pointer_q[1];
  assign N28811 = N38708 & commit_pointer_q[2];
  assign N38709 = N56 & commit_pointer_q[1];
  assign N56 = ~commit_pointer_q[0];
  assign N28810 = N38709 & commit_pointer_q[2];
  assign N38710 = commit_pointer_q[0] & N57;
  assign N57 = ~commit_pointer_q[1];
  assign N28809 = N38710 & commit_pointer_q[2];
  assign N38711 = N58 & N59;
  assign N58 = ~commit_pointer_q[0];
  assign N59 = ~commit_pointer_q[1];
  assign N28808 = N38711 & commit_pointer_q[2];
  assign N38712 = commit_pointer_q[0] & commit_pointer_q[1];
  assign N28807 = N38712 & N60;
  assign N60 = ~commit_pointer_q[2];
  assign N38713 = N61 & commit_pointer_q[1];
  assign N61 = ~commit_pointer_q[0];
  assign N28806 = N38713 & N62;
  assign N62 = ~commit_pointer_q[2];
  assign N38714 = commit_pointer_q[0] & N63;
  assign N63 = ~commit_pointer_q[1];
  assign N28805 = N38714 & N64;
  assign N64 = ~commit_pointer_q[2];
  assign N38715 = N65 & N66;
  assign N65 = ~commit_pointer_q[0];
  assign N66 = ~commit_pointer_q[1];
  assign N28804 = N38715 & N67;
  assign N67 = ~commit_pointer_q[2];
  assign N38716 = N28855 & N28856;
  assign N28865 = N38716 & N28857;
  assign N38717 = N68 & N28856;
  assign N68 = ~N28855;
  assign N28864 = N38717 & N28857;
  assign N38718 = N28855 & N69;
  assign N69 = ~N28856;
  assign N28863 = N38718 & N28857;
  assign N38719 = N70 & N71;
  assign N70 = ~N28855;
  assign N71 = ~N28856;
  assign N28862 = N38719 & N28857;
  assign N28861 = N38716 & N72;
  assign N72 = ~N28857;
  assign N28860 = N38717 & N73;
  assign N73 = ~N28857;
  assign N28859 = N38718 & N74;
  assign N74 = ~N28857;
  assign N28858 = N38719 & N75;
  assign N75 = ~N28857;
  assign N38720 = N28882 & N28883;
  assign N28892 = N38720 & N28884;
  assign N38721 = N76 & N28883;
  assign N76 = ~N28882;
  assign N28891 = N38721 & N28884;
  assign N38722 = N28882 & N77;
  assign N77 = ~N28883;
  assign N28890 = N38722 & N28884;
  assign N38723 = N78 & N79;
  assign N78 = ~N28882;
  assign N79 = ~N28883;
  assign N28889 = N38723 & N28884;
  assign N28888 = N38720 & N80;
  assign N80 = ~N28884;
  assign N28887 = N38721 & N81;
  assign N81 = ~N28884;
  assign N28886 = N38722 & N82;
  assign N82 = ~N28884;
  assign N28885 = N38723 & N83;
  assign N83 = ~N28884;
  assign N38724 = ~mem_q[271];
  assign N38725 = mem_q[269] & mem_q[270];
  assign N38726 = N84 & mem_q[270];
  assign N84 = ~mem_q[269];
  assign N38727 = mem_q[269] & N85;
  assign N85 = ~mem_q[270];
  assign N38728 = N86 & N87;
  assign N86 = ~mem_q[269];
  assign N87 = ~mem_q[270];
  assign N38729 = mem_q[271] & N38725;
  assign N38730 = mem_q[271] & N38726;
  assign N38731 = mem_q[271] & N38727;
  assign N38732 = mem_q[271] & N38728;
  assign N38733 = N38724 & N38725;
  assign N38734 = N38724 & N38726;
  assign N38735 = N38724 & N38727;
  assign N38736 = N38724 & N38728;
  assign N38737 = ~mem_q[268];
  assign N38738 = mem_q[266] & mem_q[267];
  assign N38739 = N88 & mem_q[267];
  assign N88 = ~mem_q[266];
  assign N38740 = mem_q[266] & N89;
  assign N89 = ~mem_q[267];
  assign N38741 = N90 & N91;
  assign N90 = ~mem_q[266];
  assign N91 = ~mem_q[267];
  assign N38742 = mem_q[268] & N38738;
  assign N38743 = mem_q[268] & N38739;
  assign N38744 = mem_q[268] & N38740;
  assign N38745 = mem_q[268] & N38741;
  assign N38746 = N38737 & N38738;
  assign N38747 = N38737 & N38739;
  assign N38748 = N38737 & N38740;
  assign N38749 = N38737 & N38741;
  assign N28998 = N38729 & N38742;
  assign N28997 = N38729 & N38743;
  assign N28996 = N38729 & N38744;
  assign N28995 = N38729 & N38745;
  assign N28994 = N38729 & N38746;
  assign N28993 = N38729 & N38747;
  assign N28992 = N38729 & N38748;
  assign N28991 = N38729 & N38749;
  assign N28990 = N38730 & N38742;
  assign N28989 = N38730 & N38743;
  assign N28988 = N38730 & N38744;
  assign N28987 = N38730 & N38745;
  assign N28986 = N38730 & N38746;
  assign N28985 = N38730 & N38747;
  assign N28984 = N38730 & N38748;
  assign N28983 = N38730 & N38749;
  assign N28982 = N38731 & N38742;
  assign N28981 = N38731 & N38743;
  assign N28980 = N38731 & N38744;
  assign N28979 = N38731 & N38745;
  assign N28978 = N38731 & N38746;
  assign N28977 = N38731 & N38747;
  assign N28976 = N38731 & N38748;
  assign N28975 = N38731 & N38749;
  assign N28974 = N38732 & N38742;
  assign N28973 = N38732 & N38743;
  assign N28972 = N38732 & N38744;
  assign N28971 = N38732 & N38745;
  assign N28970 = N38732 & N38746;
  assign N28969 = N38732 & N38747;
  assign N28968 = N38732 & N38748;
  assign N28967 = N38732 & N38749;
  assign N28966 = N38733 & N38742;
  assign N28965 = N38733 & N38743;
  assign N28964 = N38733 & N38744;
  assign N28963 = N38733 & N38745;
  assign N28962 = N38733 & N38746;
  assign N28961 = N38733 & N38747;
  assign N28960 = N38733 & N38748;
  assign N28959 = N38733 & N38749;
  assign N28958 = N38734 & N38742;
  assign N28957 = N38734 & N38743;
  assign N28956 = N38734 & N38744;
  assign N28955 = N38734 & N38745;
  assign N28954 = N38734 & N38746;
  assign N28953 = N38734 & N38747;
  assign N28952 = N38734 & N38748;
  assign N28951 = N38734 & N38749;
  assign N28950 = N38735 & N38742;
  assign N28949 = N38735 & N38743;
  assign N28948 = N38735 & N38744;
  assign N28947 = N38735 & N38745;
  assign N28946 = N38735 & N38746;
  assign N28945 = N38735 & N38747;
  assign N28944 = N38735 & N38748;
  assign N28943 = N38735 & N38749;
  assign N28942 = N38736 & N38742;
  assign N28941 = N38736 & N38743;
  assign N28940 = N38736 & N38744;
  assign N28939 = N38736 & N38745;
  assign N28938 = N38736 & N38746;
  assign N28937 = N38736 & N38747;
  assign N28936 = N38736 & N38748;
  assign N38750 = ~mem_q[634];
  assign N38751 = mem_q[632] & mem_q[633];
  assign N38752 = N92 & mem_q[633];
  assign N92 = ~mem_q[632];
  assign N38753 = mem_q[632] & N93;
  assign N93 = ~mem_q[633];
  assign N38754 = N94 & N95;
  assign N94 = ~mem_q[632];
  assign N95 = ~mem_q[633];
  assign N38755 = mem_q[634] & N38751;
  assign N38756 = mem_q[634] & N38752;
  assign N38757 = mem_q[634] & N38753;
  assign N38758 = mem_q[634] & N38754;
  assign N38759 = N38750 & N38751;
  assign N38760 = N38750 & N38752;
  assign N38761 = N38750 & N38753;
  assign N38762 = N38750 & N38754;
  assign N38763 = ~mem_q[631];
  assign N38764 = mem_q[629] & mem_q[630];
  assign N38765 = N96 & mem_q[630];
  assign N96 = ~mem_q[629];
  assign N38766 = mem_q[629] & N97;
  assign N97 = ~mem_q[630];
  assign N38767 = N98 & N99;
  assign N98 = ~mem_q[629];
  assign N99 = ~mem_q[630];
  assign N38768 = mem_q[631] & N38764;
  assign N38769 = mem_q[631] & N38765;
  assign N38770 = mem_q[631] & N38766;
  assign N38771 = mem_q[631] & N38767;
  assign N38772 = N38763 & N38764;
  assign N38773 = N38763 & N38765;
  assign N38774 = N38763 & N38766;
  assign N38775 = N38763 & N38767;
  assign N29629 = N38755 & N38768;
  assign N29628 = N38755 & N38769;
  assign N29627 = N38755 & N38770;
  assign N29626 = N38755 & N38771;
  assign N29625 = N38755 & N38772;
  assign N29624 = N38755 & N38773;
  assign N29623 = N38755 & N38774;
  assign N29622 = N38755 & N38775;
  assign N29621 = N38756 & N38768;
  assign N29620 = N38756 & N38769;
  assign N29619 = N38756 & N38770;
  assign N29618 = N38756 & N38771;
  assign N29617 = N38756 & N38772;
  assign N29616 = N38756 & N38773;
  assign N29615 = N38756 & N38774;
  assign N29614 = N38756 & N38775;
  assign N29613 = N38757 & N38768;
  assign N29612 = N38757 & N38769;
  assign N29611 = N38757 & N38770;
  assign N29610 = N38757 & N38771;
  assign N29609 = N38757 & N38772;
  assign N29608 = N38757 & N38773;
  assign N29607 = N38757 & N38774;
  assign N29606 = N38757 & N38775;
  assign N29605 = N38758 & N38768;
  assign N29604 = N38758 & N38769;
  assign N29603 = N38758 & N38770;
  assign N29602 = N38758 & N38771;
  assign N29601 = N38758 & N38772;
  assign N29600 = N38758 & N38773;
  assign N29599 = N38758 & N38774;
  assign N29598 = N38758 & N38775;
  assign N29597 = N38759 & N38768;
  assign N29596 = N38759 & N38769;
  assign N29595 = N38759 & N38770;
  assign N29594 = N38759 & N38771;
  assign N29593 = N38759 & N38772;
  assign N29592 = N38759 & N38773;
  assign N29591 = N38759 & N38774;
  assign N29590 = N38759 & N38775;
  assign N29589 = N38760 & N38768;
  assign N29588 = N38760 & N38769;
  assign N29587 = N38760 & N38770;
  assign N29586 = N38760 & N38771;
  assign N29585 = N38760 & N38772;
  assign N29584 = N38760 & N38773;
  assign N29583 = N38760 & N38774;
  assign N29582 = N38760 & N38775;
  assign N29581 = N38761 & N38768;
  assign N29580 = N38761 & N38769;
  assign N29579 = N38761 & N38770;
  assign N29578 = N38761 & N38771;
  assign N29577 = N38761 & N38772;
  assign N29576 = N38761 & N38773;
  assign N29575 = N38761 & N38774;
  assign N29574 = N38761 & N38775;
  assign N29573 = N38762 & N38768;
  assign N29572 = N38762 & N38769;
  assign N29571 = N38762 & N38770;
  assign N29570 = N38762 & N38771;
  assign N29569 = N38762 & N38772;
  assign N29568 = N38762 & N38773;
  assign N29567 = N38762 & N38774;
  assign N38776 = ~mem_q[997];
  assign N38777 = mem_q[995] & mem_q[996];
  assign N38778 = N100 & mem_q[996];
  assign N100 = ~mem_q[995];
  assign N38779 = mem_q[995] & N101;
  assign N101 = ~mem_q[996];
  assign N38780 = N102 & N103;
  assign N102 = ~mem_q[995];
  assign N103 = ~mem_q[996];
  assign N38781 = mem_q[997] & N38777;
  assign N38782 = mem_q[997] & N38778;
  assign N38783 = mem_q[997] & N38779;
  assign N38784 = mem_q[997] & N38780;
  assign N38785 = N38776 & N38777;
  assign N38786 = N38776 & N38778;
  assign N38787 = N38776 & N38779;
  assign N38788 = N38776 & N38780;
  assign N38789 = ~mem_q[994];
  assign N38790 = mem_q[992] & mem_q[993];
  assign N38791 = N104 & mem_q[993];
  assign N104 = ~mem_q[992];
  assign N38792 = mem_q[992] & N105;
  assign N105 = ~mem_q[993];
  assign N38793 = N106 & N107;
  assign N106 = ~mem_q[992];
  assign N107 = ~mem_q[993];
  assign N38794 = mem_q[994] & N38790;
  assign N38795 = mem_q[994] & N38791;
  assign N38796 = mem_q[994] & N38792;
  assign N38797 = mem_q[994] & N38793;
  assign N38798 = N38789 & N38790;
  assign N38799 = N38789 & N38791;
  assign N38800 = N38789 & N38792;
  assign N38801 = N38789 & N38793;
  assign N30260 = N38781 & N38794;
  assign N30259 = N38781 & N38795;
  assign N30258 = N38781 & N38796;
  assign N30257 = N38781 & N38797;
  assign N30256 = N38781 & N38798;
  assign N30255 = N38781 & N38799;
  assign N30254 = N38781 & N38800;
  assign N30253 = N38781 & N38801;
  assign N30252 = N38782 & N38794;
  assign N30251 = N38782 & N38795;
  assign N30250 = N38782 & N38796;
  assign N30249 = N38782 & N38797;
  assign N30248 = N38782 & N38798;
  assign N30247 = N38782 & N38799;
  assign N30246 = N38782 & N38800;
  assign N30245 = N38782 & N38801;
  assign N30244 = N38783 & N38794;
  assign N30243 = N38783 & N38795;
  assign N30242 = N38783 & N38796;
  assign N30241 = N38783 & N38797;
  assign N30240 = N38783 & N38798;
  assign N30239 = N38783 & N38799;
  assign N30238 = N38783 & N38800;
  assign N30237 = N38783 & N38801;
  assign N30236 = N38784 & N38794;
  assign N30235 = N38784 & N38795;
  assign N30234 = N38784 & N38796;
  assign N30233 = N38784 & N38797;
  assign N30232 = N38784 & N38798;
  assign N30231 = N38784 & N38799;
  assign N30230 = N38784 & N38800;
  assign N30229 = N38784 & N38801;
  assign N30228 = N38785 & N38794;
  assign N30227 = N38785 & N38795;
  assign N30226 = N38785 & N38796;
  assign N30225 = N38785 & N38797;
  assign N30224 = N38785 & N38798;
  assign N30223 = N38785 & N38799;
  assign N30222 = N38785 & N38800;
  assign N30221 = N38785 & N38801;
  assign N30220 = N38786 & N38794;
  assign N30219 = N38786 & N38795;
  assign N30218 = N38786 & N38796;
  assign N30217 = N38786 & N38797;
  assign N30216 = N38786 & N38798;
  assign N30215 = N38786 & N38799;
  assign N30214 = N38786 & N38800;
  assign N30213 = N38786 & N38801;
  assign N30212 = N38787 & N38794;
  assign N30211 = N38787 & N38795;
  assign N30210 = N38787 & N38796;
  assign N30209 = N38787 & N38797;
  assign N30208 = N38787 & N38798;
  assign N30207 = N38787 & N38799;
  assign N30206 = N38787 & N38800;
  assign N30205 = N38787 & N38801;
  assign N30204 = N38788 & N38794;
  assign N30203 = N38788 & N38795;
  assign N30202 = N38788 & N38796;
  assign N30201 = N38788 & N38797;
  assign N30200 = N38788 & N38798;
  assign N30199 = N38788 & N38799;
  assign N30198 = N38788 & N38800;
  assign N38802 = ~mem_q[1360];
  assign N38803 = mem_q[1358] & mem_q[1359];
  assign N38804 = N108 & mem_q[1359];
  assign N108 = ~mem_q[1358];
  assign N38805 = mem_q[1358] & N109;
  assign N109 = ~mem_q[1359];
  assign N38806 = N110 & N111;
  assign N110 = ~mem_q[1358];
  assign N111 = ~mem_q[1359];
  assign N38807 = mem_q[1360] & N38803;
  assign N38808 = mem_q[1360] & N38804;
  assign N38809 = mem_q[1360] & N38805;
  assign N38810 = mem_q[1360] & N38806;
  assign N38811 = N38802 & N38803;
  assign N38812 = N38802 & N38804;
  assign N38813 = N38802 & N38805;
  assign N38814 = N38802 & N38806;
  assign N38815 = ~mem_q[1357];
  assign N38816 = mem_q[1355] & mem_q[1356];
  assign N38817 = N112 & mem_q[1356];
  assign N112 = ~mem_q[1355];
  assign N38818 = mem_q[1355] & N113;
  assign N113 = ~mem_q[1356];
  assign N38819 = N114 & N115;
  assign N114 = ~mem_q[1355];
  assign N115 = ~mem_q[1356];
  assign N38820 = mem_q[1357] & N38816;
  assign N38821 = mem_q[1357] & N38817;
  assign N38822 = mem_q[1357] & N38818;
  assign N38823 = mem_q[1357] & N38819;
  assign N38824 = N38815 & N38816;
  assign N38825 = N38815 & N38817;
  assign N38826 = N38815 & N38818;
  assign N38827 = N38815 & N38819;
  assign N30891 = N38807 & N38820;
  assign N30890 = N38807 & N38821;
  assign N30889 = N38807 & N38822;
  assign N30888 = N38807 & N38823;
  assign N30887 = N38807 & N38824;
  assign N30886 = N38807 & N38825;
  assign N30885 = N38807 & N38826;
  assign N30884 = N38807 & N38827;
  assign N30883 = N38808 & N38820;
  assign N30882 = N38808 & N38821;
  assign N30881 = N38808 & N38822;
  assign N30880 = N38808 & N38823;
  assign N30879 = N38808 & N38824;
  assign N30878 = N38808 & N38825;
  assign N30877 = N38808 & N38826;
  assign N30876 = N38808 & N38827;
  assign N30875 = N38809 & N38820;
  assign N30874 = N38809 & N38821;
  assign N30873 = N38809 & N38822;
  assign N30872 = N38809 & N38823;
  assign N30871 = N38809 & N38824;
  assign N30870 = N38809 & N38825;
  assign N30869 = N38809 & N38826;
  assign N30868 = N38809 & N38827;
  assign N30867 = N38810 & N38820;
  assign N30866 = N38810 & N38821;
  assign N30865 = N38810 & N38822;
  assign N30864 = N38810 & N38823;
  assign N30863 = N38810 & N38824;
  assign N30862 = N38810 & N38825;
  assign N30861 = N38810 & N38826;
  assign N30860 = N38810 & N38827;
  assign N30859 = N38811 & N38820;
  assign N30858 = N38811 & N38821;
  assign N30857 = N38811 & N38822;
  assign N30856 = N38811 & N38823;
  assign N30855 = N38811 & N38824;
  assign N30854 = N38811 & N38825;
  assign N30853 = N38811 & N38826;
  assign N30852 = N38811 & N38827;
  assign N30851 = N38812 & N38820;
  assign N30850 = N38812 & N38821;
  assign N30849 = N38812 & N38822;
  assign N30848 = N38812 & N38823;
  assign N30847 = N38812 & N38824;
  assign N30846 = N38812 & N38825;
  assign N30845 = N38812 & N38826;
  assign N30844 = N38812 & N38827;
  assign N30843 = N38813 & N38820;
  assign N30842 = N38813 & N38821;
  assign N30841 = N38813 & N38822;
  assign N30840 = N38813 & N38823;
  assign N30839 = N38813 & N38824;
  assign N30838 = N38813 & N38825;
  assign N30837 = N38813 & N38826;
  assign N30836 = N38813 & N38827;
  assign N30835 = N38814 & N38820;
  assign N30834 = N38814 & N38821;
  assign N30833 = N38814 & N38822;
  assign N30832 = N38814 & N38823;
  assign N30831 = N38814 & N38824;
  assign N30830 = N38814 & N38825;
  assign N30829 = N38814 & N38826;
  assign N38828 = ~mem_q[1723];
  assign N38829 = mem_q[1721] & mem_q[1722];
  assign N38830 = N116 & mem_q[1722];
  assign N116 = ~mem_q[1721];
  assign N38831 = mem_q[1721] & N117;
  assign N117 = ~mem_q[1722];
  assign N38832 = N118 & N119;
  assign N118 = ~mem_q[1721];
  assign N119 = ~mem_q[1722];
  assign N38833 = mem_q[1723] & N38829;
  assign N38834 = mem_q[1723] & N38830;
  assign N38835 = mem_q[1723] & N38831;
  assign N38836 = mem_q[1723] & N38832;
  assign N38837 = N38828 & N38829;
  assign N38838 = N38828 & N38830;
  assign N38839 = N38828 & N38831;
  assign N38840 = N38828 & N38832;
  assign N38841 = ~mem_q[1720];
  assign N38842 = mem_q[1718] & mem_q[1719];
  assign N38843 = N120 & mem_q[1719];
  assign N120 = ~mem_q[1718];
  assign N38844 = mem_q[1718] & N121;
  assign N121 = ~mem_q[1719];
  assign N38845 = N122 & N123;
  assign N122 = ~mem_q[1718];
  assign N123 = ~mem_q[1719];
  assign N38846 = mem_q[1720] & N38842;
  assign N38847 = mem_q[1720] & N38843;
  assign N38848 = mem_q[1720] & N38844;
  assign N38849 = mem_q[1720] & N38845;
  assign N38850 = N38841 & N38842;
  assign N38851 = N38841 & N38843;
  assign N38852 = N38841 & N38844;
  assign N38853 = N38841 & N38845;
  assign N31522 = N38833 & N38846;
  assign N31521 = N38833 & N38847;
  assign N31520 = N38833 & N38848;
  assign N31519 = N38833 & N38849;
  assign N31518 = N38833 & N38850;
  assign N31517 = N38833 & N38851;
  assign N31516 = N38833 & N38852;
  assign N31515 = N38833 & N38853;
  assign N31514 = N38834 & N38846;
  assign N31513 = N38834 & N38847;
  assign N31512 = N38834 & N38848;
  assign N31511 = N38834 & N38849;
  assign N31510 = N38834 & N38850;
  assign N31509 = N38834 & N38851;
  assign N31508 = N38834 & N38852;
  assign N31507 = N38834 & N38853;
  assign N31506 = N38835 & N38846;
  assign N31505 = N38835 & N38847;
  assign N31504 = N38835 & N38848;
  assign N31503 = N38835 & N38849;
  assign N31502 = N38835 & N38850;
  assign N31501 = N38835 & N38851;
  assign N31500 = N38835 & N38852;
  assign N31499 = N38835 & N38853;
  assign N31498 = N38836 & N38846;
  assign N31497 = N38836 & N38847;
  assign N31496 = N38836 & N38848;
  assign N31495 = N38836 & N38849;
  assign N31494 = N38836 & N38850;
  assign N31493 = N38836 & N38851;
  assign N31492 = N38836 & N38852;
  assign N31491 = N38836 & N38853;
  assign N31490 = N38837 & N38846;
  assign N31489 = N38837 & N38847;
  assign N31488 = N38837 & N38848;
  assign N31487 = N38837 & N38849;
  assign N31486 = N38837 & N38850;
  assign N31485 = N38837 & N38851;
  assign N31484 = N38837 & N38852;
  assign N31483 = N38837 & N38853;
  assign N31482 = N38838 & N38846;
  assign N31481 = N38838 & N38847;
  assign N31480 = N38838 & N38848;
  assign N31479 = N38838 & N38849;
  assign N31478 = N38838 & N38850;
  assign N31477 = N38838 & N38851;
  assign N31476 = N38838 & N38852;
  assign N31475 = N38838 & N38853;
  assign N31474 = N38839 & N38846;
  assign N31473 = N38839 & N38847;
  assign N31472 = N38839 & N38848;
  assign N31471 = N38839 & N38849;
  assign N31470 = N38839 & N38850;
  assign N31469 = N38839 & N38851;
  assign N31468 = N38839 & N38852;
  assign N31467 = N38839 & N38853;
  assign N31466 = N38840 & N38846;
  assign N31465 = N38840 & N38847;
  assign N31464 = N38840 & N38848;
  assign N31463 = N38840 & N38849;
  assign N31462 = N38840 & N38850;
  assign N31461 = N38840 & N38851;
  assign N31460 = N38840 & N38852;
  assign N38854 = ~mem_q[2086];
  assign N38855 = mem_q[2084] & mem_q[2085];
  assign N38856 = N124 & mem_q[2085];
  assign N124 = ~mem_q[2084];
  assign N38857 = mem_q[2084] & N125;
  assign N125 = ~mem_q[2085];
  assign N38858 = N126 & N127;
  assign N126 = ~mem_q[2084];
  assign N127 = ~mem_q[2085];
  assign N38859 = mem_q[2086] & N38855;
  assign N38860 = mem_q[2086] & N38856;
  assign N38861 = mem_q[2086] & N38857;
  assign N38862 = mem_q[2086] & N38858;
  assign N38863 = N38854 & N38855;
  assign N38864 = N38854 & N38856;
  assign N38865 = N38854 & N38857;
  assign N38866 = N38854 & N38858;
  assign N38867 = ~mem_q[2083];
  assign N38868 = mem_q[2081] & mem_q[2082];
  assign N38869 = N128 & mem_q[2082];
  assign N128 = ~mem_q[2081];
  assign N38870 = mem_q[2081] & N129;
  assign N129 = ~mem_q[2082];
  assign N38871 = N130 & N131;
  assign N130 = ~mem_q[2081];
  assign N131 = ~mem_q[2082];
  assign N38872 = mem_q[2083] & N38868;
  assign N38873 = mem_q[2083] & N38869;
  assign N38874 = mem_q[2083] & N38870;
  assign N38875 = mem_q[2083] & N38871;
  assign N38876 = N38867 & N38868;
  assign N38877 = N38867 & N38869;
  assign N38878 = N38867 & N38870;
  assign N38879 = N38867 & N38871;
  assign N32153 = N38859 & N38872;
  assign N32152 = N38859 & N38873;
  assign N32151 = N38859 & N38874;
  assign N32150 = N38859 & N38875;
  assign N32149 = N38859 & N38876;
  assign N32148 = N38859 & N38877;
  assign N32147 = N38859 & N38878;
  assign N32146 = N38859 & N38879;
  assign N32145 = N38860 & N38872;
  assign N32144 = N38860 & N38873;
  assign N32143 = N38860 & N38874;
  assign N32142 = N38860 & N38875;
  assign N32141 = N38860 & N38876;
  assign N32140 = N38860 & N38877;
  assign N32139 = N38860 & N38878;
  assign N32138 = N38860 & N38879;
  assign N32137 = N38861 & N38872;
  assign N32136 = N38861 & N38873;
  assign N32135 = N38861 & N38874;
  assign N32134 = N38861 & N38875;
  assign N32133 = N38861 & N38876;
  assign N32132 = N38861 & N38877;
  assign N32131 = N38861 & N38878;
  assign N32130 = N38861 & N38879;
  assign N32129 = N38862 & N38872;
  assign N32128 = N38862 & N38873;
  assign N32127 = N38862 & N38874;
  assign N32126 = N38862 & N38875;
  assign N32125 = N38862 & N38876;
  assign N32124 = N38862 & N38877;
  assign N32123 = N38862 & N38878;
  assign N32122 = N38862 & N38879;
  assign N32121 = N38863 & N38872;
  assign N32120 = N38863 & N38873;
  assign N32119 = N38863 & N38874;
  assign N32118 = N38863 & N38875;
  assign N32117 = N38863 & N38876;
  assign N32116 = N38863 & N38877;
  assign N32115 = N38863 & N38878;
  assign N32114 = N38863 & N38879;
  assign N32113 = N38864 & N38872;
  assign N32112 = N38864 & N38873;
  assign N32111 = N38864 & N38874;
  assign N32110 = N38864 & N38875;
  assign N32109 = N38864 & N38876;
  assign N32108 = N38864 & N38877;
  assign N32107 = N38864 & N38878;
  assign N32106 = N38864 & N38879;
  assign N32105 = N38865 & N38872;
  assign N32104 = N38865 & N38873;
  assign N32103 = N38865 & N38874;
  assign N32102 = N38865 & N38875;
  assign N32101 = N38865 & N38876;
  assign N32100 = N38865 & N38877;
  assign N32099 = N38865 & N38878;
  assign N32098 = N38865 & N38879;
  assign N32097 = N38866 & N38872;
  assign N32096 = N38866 & N38873;
  assign N32095 = N38866 & N38874;
  assign N32094 = N38866 & N38875;
  assign N32093 = N38866 & N38876;
  assign N32092 = N38866 & N38877;
  assign N32091 = N38866 & N38878;
  assign N38880 = ~mem_q[2449];
  assign N38881 = mem_q[2447] & mem_q[2448];
  assign N38882 = N132 & mem_q[2448];
  assign N132 = ~mem_q[2447];
  assign N38883 = mem_q[2447] & N133;
  assign N133 = ~mem_q[2448];
  assign N38884 = N134 & N135;
  assign N134 = ~mem_q[2447];
  assign N135 = ~mem_q[2448];
  assign N38885 = mem_q[2449] & N38881;
  assign N38886 = mem_q[2449] & N38882;
  assign N38887 = mem_q[2449] & N38883;
  assign N38888 = mem_q[2449] & N38884;
  assign N38889 = N38880 & N38881;
  assign N38890 = N38880 & N38882;
  assign N38891 = N38880 & N38883;
  assign N38892 = N38880 & N38884;
  assign N38893 = ~mem_q[2446];
  assign N38894 = mem_q[2444] & mem_q[2445];
  assign N38895 = N136 & mem_q[2445];
  assign N136 = ~mem_q[2444];
  assign N38896 = mem_q[2444] & N137;
  assign N137 = ~mem_q[2445];
  assign N38897 = N138 & N139;
  assign N138 = ~mem_q[2444];
  assign N139 = ~mem_q[2445];
  assign N38898 = mem_q[2446] & N38894;
  assign N38899 = mem_q[2446] & N38895;
  assign N38900 = mem_q[2446] & N38896;
  assign N38901 = mem_q[2446] & N38897;
  assign N38902 = N38893 & N38894;
  assign N38903 = N38893 & N38895;
  assign N38904 = N38893 & N38896;
  assign N38905 = N38893 & N38897;
  assign N32784 = N38885 & N38898;
  assign N32783 = N38885 & N38899;
  assign N32782 = N38885 & N38900;
  assign N32781 = N38885 & N38901;
  assign N32780 = N38885 & N38902;
  assign N32779 = N38885 & N38903;
  assign N32778 = N38885 & N38904;
  assign N32777 = N38885 & N38905;
  assign N32776 = N38886 & N38898;
  assign N32775 = N38886 & N38899;
  assign N32774 = N38886 & N38900;
  assign N32773 = N38886 & N38901;
  assign N32772 = N38886 & N38902;
  assign N32771 = N38886 & N38903;
  assign N32770 = N38886 & N38904;
  assign N32769 = N38886 & N38905;
  assign N32768 = N38887 & N38898;
  assign N32767 = N38887 & N38899;
  assign N32766 = N38887 & N38900;
  assign N32765 = N38887 & N38901;
  assign N32764 = N38887 & N38902;
  assign N32763 = N38887 & N38903;
  assign N32762 = N38887 & N38904;
  assign N32761 = N38887 & N38905;
  assign N32760 = N38888 & N38898;
  assign N32759 = N38888 & N38899;
  assign N32758 = N38888 & N38900;
  assign N32757 = N38888 & N38901;
  assign N32756 = N38888 & N38902;
  assign N32755 = N38888 & N38903;
  assign N32754 = N38888 & N38904;
  assign N32753 = N38888 & N38905;
  assign N32752 = N38889 & N38898;
  assign N32751 = N38889 & N38899;
  assign N32750 = N38889 & N38900;
  assign N32749 = N38889 & N38901;
  assign N32748 = N38889 & N38902;
  assign N32747 = N38889 & N38903;
  assign N32746 = N38889 & N38904;
  assign N32745 = N38889 & N38905;
  assign N32744 = N38890 & N38898;
  assign N32743 = N38890 & N38899;
  assign N32742 = N38890 & N38900;
  assign N32741 = N38890 & N38901;
  assign N32740 = N38890 & N38902;
  assign N32739 = N38890 & N38903;
  assign N32738 = N38890 & N38904;
  assign N32737 = N38890 & N38905;
  assign N32736 = N38891 & N38898;
  assign N32735 = N38891 & N38899;
  assign N32734 = N38891 & N38900;
  assign N32733 = N38891 & N38901;
  assign N32732 = N38891 & N38902;
  assign N32731 = N38891 & N38903;
  assign N32730 = N38891 & N38904;
  assign N32729 = N38891 & N38905;
  assign N32728 = N38892 & N38898;
  assign N32727 = N38892 & N38899;
  assign N32726 = N38892 & N38900;
  assign N32725 = N38892 & N38901;
  assign N32724 = N38892 & N38902;
  assign N32723 = N38892 & N38903;
  assign N32722 = N38892 & N38904;
  assign N38906 = ~mem_q[2812];
  assign N38907 = mem_q[2810] & mem_q[2811];
  assign N38908 = N140 & mem_q[2811];
  assign N140 = ~mem_q[2810];
  assign N38909 = mem_q[2810] & N141;
  assign N141 = ~mem_q[2811];
  assign N38910 = N142 & N143;
  assign N142 = ~mem_q[2810];
  assign N143 = ~mem_q[2811];
  assign N38911 = mem_q[2812] & N38907;
  assign N38912 = mem_q[2812] & N38908;
  assign N38913 = mem_q[2812] & N38909;
  assign N38914 = mem_q[2812] & N38910;
  assign N38915 = N38906 & N38907;
  assign N38916 = N38906 & N38908;
  assign N38917 = N38906 & N38909;
  assign N38918 = N38906 & N38910;
  assign N38919 = ~mem_q[2809];
  assign N38920 = mem_q[2807] & mem_q[2808];
  assign N38921 = N144 & mem_q[2808];
  assign N144 = ~mem_q[2807];
  assign N38922 = mem_q[2807] & N145;
  assign N145 = ~mem_q[2808];
  assign N38923 = N146 & N147;
  assign N146 = ~mem_q[2807];
  assign N147 = ~mem_q[2808];
  assign N38924 = mem_q[2809] & N38920;
  assign N38925 = mem_q[2809] & N38921;
  assign N38926 = mem_q[2809] & N38922;
  assign N38927 = mem_q[2809] & N38923;
  assign N38928 = N38919 & N38920;
  assign N38929 = N38919 & N38921;
  assign N38930 = N38919 & N38922;
  assign N38931 = N38919 & N38923;
  assign N33415 = N38911 & N38924;
  assign N33414 = N38911 & N38925;
  assign N33413 = N38911 & N38926;
  assign N33412 = N38911 & N38927;
  assign N33411 = N38911 & N38928;
  assign N33410 = N38911 & N38929;
  assign N33409 = N38911 & N38930;
  assign N33408 = N38911 & N38931;
  assign N33407 = N38912 & N38924;
  assign N33406 = N38912 & N38925;
  assign N33405 = N38912 & N38926;
  assign N33404 = N38912 & N38927;
  assign N33403 = N38912 & N38928;
  assign N33402 = N38912 & N38929;
  assign N33401 = N38912 & N38930;
  assign N33400 = N38912 & N38931;
  assign N33399 = N38913 & N38924;
  assign N33398 = N38913 & N38925;
  assign N33397 = N38913 & N38926;
  assign N33396 = N38913 & N38927;
  assign N33395 = N38913 & N38928;
  assign N33394 = N38913 & N38929;
  assign N33393 = N38913 & N38930;
  assign N33392 = N38913 & N38931;
  assign N33391 = N38914 & N38924;
  assign N33390 = N38914 & N38925;
  assign N33389 = N38914 & N38926;
  assign N33388 = N38914 & N38927;
  assign N33387 = N38914 & N38928;
  assign N33386 = N38914 & N38929;
  assign N33385 = N38914 & N38930;
  assign N33384 = N38914 & N38931;
  assign N33383 = N38915 & N38924;
  assign N33382 = N38915 & N38925;
  assign N33381 = N38915 & N38926;
  assign N33380 = N38915 & N38927;
  assign N33379 = N38915 & N38928;
  assign N33378 = N38915 & N38929;
  assign N33377 = N38915 & N38930;
  assign N33376 = N38915 & N38931;
  assign N33375 = N38916 & N38924;
  assign N33374 = N38916 & N38925;
  assign N33373 = N38916 & N38926;
  assign N33372 = N38916 & N38927;
  assign N33371 = N38916 & N38928;
  assign N33370 = N38916 & N38929;
  assign N33369 = N38916 & N38930;
  assign N33368 = N38916 & N38931;
  assign N33367 = N38917 & N38924;
  assign N33366 = N38917 & N38925;
  assign N33365 = N38917 & N38926;
  assign N33364 = N38917 & N38927;
  assign N33363 = N38917 & N38928;
  assign N33362 = N38917 & N38929;
  assign N33361 = N38917 & N38930;
  assign N33360 = N38917 & N38931;
  assign N33359 = N38918 & N38924;
  assign N33358 = N38918 & N38925;
  assign N33357 = N38918 & N38926;
  assign N33356 = N38918 & N38927;
  assign N33355 = N38918 & N38928;
  assign N33354 = N38918 & N38929;
  assign N33353 = N38918 & N38930;
  assign { N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897 } = (N148)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N896)? { mem_q[0:0], mem_q[1:1], mem_q[2:2], mem_q[3:3], mem_q[4:4], mem_q[5:5], mem_q[6:6], mem_q[7:7], mem_q[8:8], mem_q[9:9], mem_q[10:10], mem_q[11:11], mem_q[12:12], mem_q[13:13], mem_q[14:14], mem_q[15:15], mem_q[16:16], mem_q[17:17], mem_q[18:18], mem_q[19:19], mem_q[20:20], mem_q[21:21], mem_q[22:22], mem_q[23:23], mem_q[24:24], mem_q[25:25], mem_q[26:26], mem_q[27:27], mem_q[28:28], mem_q[29:29], mem_q[30:30], mem_q[31:31], mem_q[32:32], mem_q[33:33], mem_q[34:34], mem_q[35:35], mem_q[36:36], mem_q[37:37], mem_q[38:38], mem_q[39:39], mem_q[40:40], mem_q[41:41], mem_q[42:42], mem_q[43:43], mem_q[44:44], mem_q[45:45], mem_q[46:46], mem_q[47:47], mem_q[48:48], mem_q[49:49], mem_q[50:50], mem_q[51:51], mem_q[52:52], mem_q[53:53], mem_q[54:54], mem_q[55:55], mem_q[56:56], mem_q[57:57], mem_q[58:58], mem_q[59:59], mem_q[60:60], mem_q[61:61], mem_q[62:62], mem_q[63:63], mem_q[64:64], mem_q[65:65], mem_q[66:66], mem_q[67:67], mem_q[68:68], mem_q[69:69], mem_q[70:70], mem_q[71:71], mem_q[72:72], mem_q[73:73], mem_q[74:74], mem_q[75:75], mem_q[76:76], mem_q[77:77], mem_q[78:78], mem_q[79:79], mem_q[80:80], mem_q[81:81], mem_q[82:82], mem_q[83:83], mem_q[84:84], mem_q[85:85], mem_q[86:86], mem_q[87:87], mem_q[88:88], mem_q[89:89], mem_q[90:90], mem_q[91:91], mem_q[92:92], mem_q[93:93], mem_q[94:94], mem_q[95:95], mem_q[96:96], mem_q[97:97], mem_q[98:98], mem_q[99:99], mem_q[100:100], mem_q[101:101], mem_q[102:102], mem_q[103:103], mem_q[104:104], mem_q[105:105], mem_q[106:106], mem_q[107:107], mem_q[108:108], mem_q[109:109], mem_q[110:110], mem_q[111:111], mem_q[112:112], mem_q[113:113], mem_q[114:114], mem_q[115:115], mem_q[116:116], mem_q[117:117], mem_q[118:118], mem_q[119:119], mem_q[120:120], mem_q[121:121], mem_q[122:122], mem_q[123:123], mem_q[124:124], mem_q[125:125], mem_q[126:126], mem_q[127:127], mem_q[128:128], mem_q[129:129], mem_q[130:130], mem_q[131:131], mem_q[132:132], mem_q[133:133], mem_q[134:134], mem_q[135:135], mem_q[136:136], mem_q[137:137], mem_q[138:138], mem_q[139:139], mem_q[140:140], mem_q[141:141], mem_q[142:142], mem_q[143:143], mem_q[144:144], mem_q[145:145], mem_q[146:146], mem_q[147:147], mem_q[148:148], mem_q[149:149], mem_q[150:150], mem_q[151:151], mem_q[152:152], mem_q[153:153], mem_q[154:154], mem_q[155:155], mem_q[156:156], mem_q[157:157], mem_q[158:158], mem_q[159:159], mem_q[160:160], mem_q[161:161], mem_q[162:162], mem_q[163:163], mem_q[164:164], mem_q[165:165], mem_q[166:166], mem_q[167:167], mem_q[168:168], mem_q[169:169], mem_q[170:170], mem_q[171:171], mem_q[172:172], mem_q[173:173], mem_q[174:174], mem_q[175:175], mem_q[176:176], mem_q[177:177], mem_q[178:178], mem_q[179:179], mem_q[180:180], mem_q[181:181], mem_q[182:182], mem_q[183:183], mem_q[184:184], mem_q[185:185], mem_q[186:186], mem_q[187:187], mem_q[188:188], mem_q[189:189], mem_q[190:190], mem_q[191:191], mem_q[192:192], mem_q[193:193], mem_q[194:194], mem_q[195:195], mem_q[196:196], mem_q[197:197], mem_q[198:198], mem_q[199:199], mem_q[200:200], mem_q[201:201], mem_q[202:202], mem_q[203:203], mem_q[204:204], mem_q[205:205], mem_q[206:206], mem_q[207:207], mem_q[208:208], mem_q[209:209], mem_q[210:210], mem_q[211:211], mem_q[212:212], mem_q[213:213], mem_q[214:214], mem_q[215:215], mem_q[216:216], mem_q[217:217], mem_q[218:218], mem_q[219:219], mem_q[220:220], mem_q[221:221], mem_q[222:222], mem_q[223:223], mem_q[224:224], mem_q[225:225], mem_q[226:226], mem_q[227:227], mem_q[228:228], mem_q[229:229], mem_q[230:230], mem_q[231:231], mem_q[232:232], mem_q[233:233], mem_q[234:234], mem_q[235:235], mem_q[236:236], mem_q[237:237], mem_q[238:238], mem_q[239:239], mem_q[240:240], mem_q[241:241], mem_q[242:242], mem_q[243:243], mem_q[244:244], mem_q[245:245], mem_q[246:246], mem_q[247:247], mem_q[248:248], mem_q[249:249], mem_q[250:250], mem_q[251:251], mem_q[252:252], mem_q[253:253], mem_q[254:254], mem_q[255:255], mem_q[256:256], mem_q[257:257], mem_q[258:258], mem_q[259:259], mem_q[260:260], mem_q[261:261], mem_q[262:262], mem_q[263:263], mem_q[264:264], mem_q[265:265], mem_q[266:266], mem_q[267:267], mem_q[268:268], mem_q[269:269], mem_q[270:270], mem_q[271:271], mem_q[272:272], mem_q[273:273], mem_q[274:274], mem_q[275:275], mem_q[276:276], mem_q[277:277], mem_q[278:278], mem_q[279:279], mem_q[280:280], mem_q[281:281], mem_q[282:282], mem_q[283:283], mem_q[284:284], mem_q[285:285], mem_q[286:286], mem_q[287:287], mem_q[288:288], mem_q[289:289], mem_q[290:290], mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294], mem_q[295:295], mem_q[296:296], mem_q[297:297], mem_q[298:298], mem_q[299:299], mem_q[300:300], mem_q[301:301], mem_q[302:302], mem_q[303:303], mem_q[304:304], mem_q[305:305], mem_q[306:306], mem_q[307:307], mem_q[308:308], mem_q[309:309], mem_q[310:310], mem_q[311:311], mem_q[312:312], mem_q[313:313], mem_q[314:314], mem_q[315:315], mem_q[316:316], mem_q[317:317], mem_q[318:318], mem_q[319:319], mem_q[320:320], mem_q[321:321], mem_q[322:322], mem_q[323:323], mem_q[324:324], mem_q[325:325], mem_q[326:326], mem_q[327:327], mem_q[328:328], mem_q[329:329], mem_q[330:330], mem_q[331:331], mem_q[332:332], mem_q[333:333], mem_q[334:334], mem_q[335:335], mem_q[336:336], mem_q[337:337], mem_q[338:338], mem_q[339:339], mem_q[340:340], mem_q[341:341], mem_q[342:342], mem_q[343:343], mem_q[344:344], mem_q[345:345], mem_q[346:346], mem_q[347:347], mem_q[348:348], mem_q[349:349], mem_q[350:350], mem_q[351:351], mem_q[352:352], mem_q[353:353], mem_q[354:354], mem_q[355:355], mem_q[356:356], mem_q[357:357], mem_q[358:358], mem_q[359:359], mem_q[360:360], mem_q[361:361], mem_q[362:362] } : 1'b0;
  assign N148 = N888;
  assign { N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261 } = (N149)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N1260)? { mem_q[363:363], mem_q[364:364], mem_q[365:365], mem_q[366:366], mem_q[367:367], mem_q[368:368], mem_q[369:369], mem_q[370:370], mem_q[371:371], mem_q[372:372], mem_q[373:373], mem_q[374:374], mem_q[375:375], mem_q[376:376], mem_q[377:377], mem_q[378:378], mem_q[379:379], mem_q[380:380], mem_q[381:381], mem_q[382:382], mem_q[383:383], mem_q[384:384], mem_q[385:385], mem_q[386:386], mem_q[387:387], mem_q[388:388], mem_q[389:389], mem_q[390:390], mem_q[391:391], mem_q[392:392], mem_q[393:393], mem_q[394:394], mem_q[395:395], mem_q[396:396], mem_q[397:397], mem_q[398:398], mem_q[399:399], mem_q[400:400], mem_q[401:401], mem_q[402:402], mem_q[403:403], mem_q[404:404], mem_q[405:405], mem_q[406:406], mem_q[407:407], mem_q[408:408], mem_q[409:409], mem_q[410:410], mem_q[411:411], mem_q[412:412], mem_q[413:413], mem_q[414:414], mem_q[415:415], mem_q[416:416], mem_q[417:417], mem_q[418:418], mem_q[419:419], mem_q[420:420], mem_q[421:421], mem_q[422:422], mem_q[423:423], mem_q[424:424], mem_q[425:425], mem_q[426:426], mem_q[427:427], mem_q[428:428], mem_q[429:429], mem_q[430:430], mem_q[431:431], mem_q[432:432], mem_q[433:433], mem_q[434:434], mem_q[435:435], mem_q[436:436], mem_q[437:437], mem_q[438:438], mem_q[439:439], mem_q[440:440], mem_q[441:441], mem_q[442:442], mem_q[443:443], mem_q[444:444], mem_q[445:445], mem_q[446:446], mem_q[447:447], mem_q[448:448], mem_q[449:449], mem_q[450:450], mem_q[451:451], mem_q[452:452], mem_q[453:453], mem_q[454:454], mem_q[455:455], mem_q[456:456], mem_q[457:457], mem_q[458:458], mem_q[459:459], mem_q[460:460], mem_q[461:461], mem_q[462:462], mem_q[463:463], mem_q[464:464], mem_q[465:465], mem_q[466:466], mem_q[467:467], mem_q[468:468], mem_q[469:469], mem_q[470:470], mem_q[471:471], mem_q[472:472], mem_q[473:473], mem_q[474:474], mem_q[475:475], mem_q[476:476], mem_q[477:477], mem_q[478:478], mem_q[479:479], mem_q[480:480], mem_q[481:481], mem_q[482:482], mem_q[483:483], mem_q[484:484], mem_q[485:485], mem_q[486:486], mem_q[487:487], mem_q[488:488], mem_q[489:489], mem_q[490:490], mem_q[491:491], mem_q[492:492], mem_q[493:493], mem_q[494:494], mem_q[495:495], mem_q[496:496], mem_q[497:497], mem_q[498:498], mem_q[499:499], mem_q[500:500], mem_q[501:501], mem_q[502:502], mem_q[503:503], mem_q[504:504], mem_q[505:505], mem_q[506:506], mem_q[507:507], mem_q[508:508], mem_q[509:509], mem_q[510:510], mem_q[511:511], mem_q[512:512], mem_q[513:513], mem_q[514:514], mem_q[515:515], mem_q[516:516], mem_q[517:517], mem_q[518:518], mem_q[519:519], mem_q[520:520], mem_q[521:521], mem_q[522:522], mem_q[523:523], mem_q[524:524], mem_q[525:525], mem_q[526:526], mem_q[527:527], mem_q[528:528], mem_q[529:529], mem_q[530:530], mem_q[531:531], mem_q[532:532], mem_q[533:533], mem_q[534:534], mem_q[535:535], mem_q[536:536], mem_q[537:537], mem_q[538:538], mem_q[539:539], mem_q[540:540], mem_q[541:541], mem_q[542:542], mem_q[543:543], mem_q[544:544], mem_q[545:545], mem_q[546:546], mem_q[547:547], mem_q[548:548], mem_q[549:549], mem_q[550:550], mem_q[551:551], mem_q[552:552], mem_q[553:553], mem_q[554:554], mem_q[555:555], mem_q[556:556], mem_q[557:557], mem_q[558:558], mem_q[559:559], mem_q[560:560], mem_q[561:561], mem_q[562:562], mem_q[563:563], mem_q[564:564], mem_q[565:565], mem_q[566:566], mem_q[567:567], mem_q[568:568], mem_q[569:569], mem_q[570:570], mem_q[571:571], mem_q[572:572], mem_q[573:573], mem_q[574:574], mem_q[575:575], mem_q[576:576], mem_q[577:577], mem_q[578:578], mem_q[579:579], mem_q[580:580], mem_q[581:581], mem_q[582:582], mem_q[583:583], mem_q[584:584], mem_q[585:585], mem_q[586:586], mem_q[587:587], mem_q[588:588], mem_q[589:589], mem_q[590:590], mem_q[591:591], mem_q[592:592], mem_q[593:593], mem_q[594:594], mem_q[595:595], mem_q[596:596], mem_q[597:597], mem_q[598:598], mem_q[599:599], mem_q[600:600], mem_q[601:601], mem_q[602:602], mem_q[603:603], mem_q[604:604], mem_q[605:605], mem_q[606:606], mem_q[607:607], mem_q[608:608], mem_q[609:609], mem_q[610:610], mem_q[611:611], mem_q[612:612], mem_q[613:613], mem_q[614:614], mem_q[615:615], mem_q[616:616], mem_q[617:617], mem_q[618:618], mem_q[619:619], mem_q[620:620], mem_q[621:621], mem_q[622:622], mem_q[623:623], mem_q[624:624], mem_q[625:625], mem_q[626:626], mem_q[627:627], mem_q[628:628], mem_q[629:629], mem_q[630:630], mem_q[631:631], mem_q[632:632], mem_q[633:633], mem_q[634:634], mem_q[635:635], mem_q[636:636], mem_q[637:637], mem_q[638:638], mem_q[639:639], mem_q[640:640], mem_q[641:641], mem_q[642:642], mem_q[643:643], mem_q[644:644], mem_q[645:645], mem_q[646:646], mem_q[647:647], mem_q[648:648], mem_q[649:649], mem_q[650:650], mem_q[651:651], mem_q[652:652], mem_q[653:653], mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657], mem_q[658:658], mem_q[659:659], mem_q[660:660], mem_q[661:661], mem_q[662:662], mem_q[663:663], mem_q[664:664], mem_q[665:665], mem_q[666:666], mem_q[667:667], mem_q[668:668], mem_q[669:669], mem_q[670:670], mem_q[671:671], mem_q[672:672], mem_q[673:673], mem_q[674:674], mem_q[675:675], mem_q[676:676], mem_q[677:677], mem_q[678:678], mem_q[679:679], mem_q[680:680], mem_q[681:681], mem_q[682:682], mem_q[683:683], mem_q[684:684], mem_q[685:685], mem_q[686:686], mem_q[687:687], mem_q[688:688], mem_q[689:689], mem_q[690:690], mem_q[691:691], mem_q[692:692], mem_q[693:693], mem_q[694:694], mem_q[695:695], mem_q[696:696], mem_q[697:697], mem_q[698:698], mem_q[699:699], mem_q[700:700], mem_q[701:701], mem_q[702:702], mem_q[703:703], mem_q[704:704], mem_q[705:705], mem_q[706:706], mem_q[707:707], mem_q[708:708], mem_q[709:709], mem_q[710:710], mem_q[711:711], mem_q[712:712], mem_q[713:713], mem_q[714:714], mem_q[715:715], mem_q[716:716], mem_q[717:717], mem_q[718:718], mem_q[719:719], mem_q[720:720], mem_q[721:721], mem_q[722:722], mem_q[723:723], mem_q[724:724], mem_q[725:725] } : 1'b0;
  assign N149 = N889;
  assign { N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625 } = (N150)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N1624)? { mem_q[726:726], mem_q[727:727], mem_q[728:728], mem_q[729:729], mem_q[730:730], mem_q[731:731], mem_q[732:732], mem_q[733:733], mem_q[734:734], mem_q[735:735], mem_q[736:736], mem_q[737:737], mem_q[738:738], mem_q[739:739], mem_q[740:740], mem_q[741:741], mem_q[742:742], mem_q[743:743], mem_q[744:744], mem_q[745:745], mem_q[746:746], mem_q[747:747], mem_q[748:748], mem_q[749:749], mem_q[750:750], mem_q[751:751], mem_q[752:752], mem_q[753:753], mem_q[754:754], mem_q[755:755], mem_q[756:756], mem_q[757:757], mem_q[758:758], mem_q[759:759], mem_q[760:760], mem_q[761:761], mem_q[762:762], mem_q[763:763], mem_q[764:764], mem_q[765:765], mem_q[766:766], mem_q[767:767], mem_q[768:768], mem_q[769:769], mem_q[770:770], mem_q[771:771], mem_q[772:772], mem_q[773:773], mem_q[774:774], mem_q[775:775], mem_q[776:776], mem_q[777:777], mem_q[778:778], mem_q[779:779], mem_q[780:780], mem_q[781:781], mem_q[782:782], mem_q[783:783], mem_q[784:784], mem_q[785:785], mem_q[786:786], mem_q[787:787], mem_q[788:788], mem_q[789:789], mem_q[790:790], mem_q[791:791], mem_q[792:792], mem_q[793:793], mem_q[794:794], mem_q[795:795], mem_q[796:796], mem_q[797:797], mem_q[798:798], mem_q[799:799], mem_q[800:800], mem_q[801:801], mem_q[802:802], mem_q[803:803], mem_q[804:804], mem_q[805:805], mem_q[806:806], mem_q[807:807], mem_q[808:808], mem_q[809:809], mem_q[810:810], mem_q[811:811], mem_q[812:812], mem_q[813:813], mem_q[814:814], mem_q[815:815], mem_q[816:816], mem_q[817:817], mem_q[818:818], mem_q[819:819], mem_q[820:820], mem_q[821:821], mem_q[822:822], mem_q[823:823], mem_q[824:824], mem_q[825:825], mem_q[826:826], mem_q[827:827], mem_q[828:828], mem_q[829:829], mem_q[830:830], mem_q[831:831], mem_q[832:832], mem_q[833:833], mem_q[834:834], mem_q[835:835], mem_q[836:836], mem_q[837:837], mem_q[838:838], mem_q[839:839], mem_q[840:840], mem_q[841:841], mem_q[842:842], mem_q[843:843], mem_q[844:844], mem_q[845:845], mem_q[846:846], mem_q[847:847], mem_q[848:848], mem_q[849:849], mem_q[850:850], mem_q[851:851], mem_q[852:852], mem_q[853:853], mem_q[854:854], mem_q[855:855], mem_q[856:856], mem_q[857:857], mem_q[858:858], mem_q[859:859], mem_q[860:860], mem_q[861:861], mem_q[862:862], mem_q[863:863], mem_q[864:864], mem_q[865:865], mem_q[866:866], mem_q[867:867], mem_q[868:868], mem_q[869:869], mem_q[870:870], mem_q[871:871], mem_q[872:872], mem_q[873:873], mem_q[874:874], mem_q[875:875], mem_q[876:876], mem_q[877:877], mem_q[878:878], mem_q[879:879], mem_q[880:880], mem_q[881:881], mem_q[882:882], mem_q[883:883], mem_q[884:884], mem_q[885:885], mem_q[886:886], mem_q[887:887], mem_q[888:888], mem_q[889:889], mem_q[890:890], mem_q[891:891], mem_q[892:892], mem_q[893:893], mem_q[894:894], mem_q[895:895], mem_q[896:896], mem_q[897:897], mem_q[898:898], mem_q[899:899], mem_q[900:900], mem_q[901:901], mem_q[902:902], mem_q[903:903], mem_q[904:904], mem_q[905:905], mem_q[906:906], mem_q[907:907], mem_q[908:908], mem_q[909:909], mem_q[910:910], mem_q[911:911], mem_q[912:912], mem_q[913:913], mem_q[914:914], mem_q[915:915], mem_q[916:916], mem_q[917:917], mem_q[918:918], mem_q[919:919], mem_q[920:920], mem_q[921:921], mem_q[922:922], mem_q[923:923], mem_q[924:924], mem_q[925:925], mem_q[926:926], mem_q[927:927], mem_q[928:928], mem_q[929:929], mem_q[930:930], mem_q[931:931], mem_q[932:932], mem_q[933:933], mem_q[934:934], mem_q[935:935], mem_q[936:936], mem_q[937:937], mem_q[938:938], mem_q[939:939], mem_q[940:940], mem_q[941:941], mem_q[942:942], mem_q[943:943], mem_q[944:944], mem_q[945:945], mem_q[946:946], mem_q[947:947], mem_q[948:948], mem_q[949:949], mem_q[950:950], mem_q[951:951], mem_q[952:952], mem_q[953:953], mem_q[954:954], mem_q[955:955], mem_q[956:956], mem_q[957:957], mem_q[958:958], mem_q[959:959], mem_q[960:960], mem_q[961:961], mem_q[962:962], mem_q[963:963], mem_q[964:964], mem_q[965:965], mem_q[966:966], mem_q[967:967], mem_q[968:968], mem_q[969:969], mem_q[970:970], mem_q[971:971], mem_q[972:972], mem_q[973:973], mem_q[974:974], mem_q[975:975], mem_q[976:976], mem_q[977:977], mem_q[978:978], mem_q[979:979], mem_q[980:980], mem_q[981:981], mem_q[982:982], mem_q[983:983], mem_q[984:984], mem_q[985:985], mem_q[986:986], mem_q[987:987], mem_q[988:988], mem_q[989:989], mem_q[990:990], mem_q[991:991], mem_q[992:992], mem_q[993:993], mem_q[994:994], mem_q[995:995], mem_q[996:996], mem_q[997:997], mem_q[998:998], mem_q[999:999], mem_q[1000:1000], mem_q[1001:1001], mem_q[1002:1002], mem_q[1003:1003], mem_q[1004:1004], mem_q[1005:1005], mem_q[1006:1006], mem_q[1007:1007], mem_q[1008:1008], mem_q[1009:1009], mem_q[1010:1010], mem_q[1011:1011], mem_q[1012:1012], mem_q[1013:1013], mem_q[1014:1014], mem_q[1015:1015], mem_q[1016:1016], mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020], mem_q[1021:1021], mem_q[1022:1022], mem_q[1023:1023], mem_q[1024:1024], mem_q[1025:1025], mem_q[1026:1026], mem_q[1027:1027], mem_q[1028:1028], mem_q[1029:1029], mem_q[1030:1030], mem_q[1031:1031], mem_q[1032:1032], mem_q[1033:1033], mem_q[1034:1034], mem_q[1035:1035], mem_q[1036:1036], mem_q[1037:1037], mem_q[1038:1038], mem_q[1039:1039], mem_q[1040:1040], mem_q[1041:1041], mem_q[1042:1042], mem_q[1043:1043], mem_q[1044:1044], mem_q[1045:1045], mem_q[1046:1046], mem_q[1047:1047], mem_q[1048:1048], mem_q[1049:1049], mem_q[1050:1050], mem_q[1051:1051], mem_q[1052:1052], mem_q[1053:1053], mem_q[1054:1054], mem_q[1055:1055], mem_q[1056:1056], mem_q[1057:1057], mem_q[1058:1058], mem_q[1059:1059], mem_q[1060:1060], mem_q[1061:1061], mem_q[1062:1062], mem_q[1063:1063], mem_q[1064:1064], mem_q[1065:1065], mem_q[1066:1066], mem_q[1067:1067], mem_q[1068:1068], mem_q[1069:1069], mem_q[1070:1070], mem_q[1071:1071], mem_q[1072:1072], mem_q[1073:1073], mem_q[1074:1074], mem_q[1075:1075], mem_q[1076:1076], mem_q[1077:1077], mem_q[1078:1078], mem_q[1079:1079], mem_q[1080:1080], mem_q[1081:1081], mem_q[1082:1082], mem_q[1083:1083], mem_q[1084:1084], mem_q[1085:1085], mem_q[1086:1086], mem_q[1087:1087], mem_q[1088:1088] } : 1'b0;
  assign N150 = N890;
  assign { N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989 } = (N151)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N1988)? { mem_q[1089:1089], mem_q[1090:1090], mem_q[1091:1091], mem_q[1092:1092], mem_q[1093:1093], mem_q[1094:1094], mem_q[1095:1095], mem_q[1096:1096], mem_q[1097:1097], mem_q[1098:1098], mem_q[1099:1099], mem_q[1100:1100], mem_q[1101:1101], mem_q[1102:1102], mem_q[1103:1103], mem_q[1104:1104], mem_q[1105:1105], mem_q[1106:1106], mem_q[1107:1107], mem_q[1108:1108], mem_q[1109:1109], mem_q[1110:1110], mem_q[1111:1111], mem_q[1112:1112], mem_q[1113:1113], mem_q[1114:1114], mem_q[1115:1115], mem_q[1116:1116], mem_q[1117:1117], mem_q[1118:1118], mem_q[1119:1119], mem_q[1120:1120], mem_q[1121:1121], mem_q[1122:1122], mem_q[1123:1123], mem_q[1124:1124], mem_q[1125:1125], mem_q[1126:1126], mem_q[1127:1127], mem_q[1128:1128], mem_q[1129:1129], mem_q[1130:1130], mem_q[1131:1131], mem_q[1132:1132], mem_q[1133:1133], mem_q[1134:1134], mem_q[1135:1135], mem_q[1136:1136], mem_q[1137:1137], mem_q[1138:1138], mem_q[1139:1139], mem_q[1140:1140], mem_q[1141:1141], mem_q[1142:1142], mem_q[1143:1143], mem_q[1144:1144], mem_q[1145:1145], mem_q[1146:1146], mem_q[1147:1147], mem_q[1148:1148], mem_q[1149:1149], mem_q[1150:1150], mem_q[1151:1151], mem_q[1152:1152], mem_q[1153:1153], mem_q[1154:1154], mem_q[1155:1155], mem_q[1156:1156], mem_q[1157:1157], mem_q[1158:1158], mem_q[1159:1159], mem_q[1160:1160], mem_q[1161:1161], mem_q[1162:1162], mem_q[1163:1163], mem_q[1164:1164], mem_q[1165:1165], mem_q[1166:1166], mem_q[1167:1167], mem_q[1168:1168], mem_q[1169:1169], mem_q[1170:1170], mem_q[1171:1171], mem_q[1172:1172], mem_q[1173:1173], mem_q[1174:1174], mem_q[1175:1175], mem_q[1176:1176], mem_q[1177:1177], mem_q[1178:1178], mem_q[1179:1179], mem_q[1180:1180], mem_q[1181:1181], mem_q[1182:1182], mem_q[1183:1183], mem_q[1184:1184], mem_q[1185:1185], mem_q[1186:1186], mem_q[1187:1187], mem_q[1188:1188], mem_q[1189:1189], mem_q[1190:1190], mem_q[1191:1191], mem_q[1192:1192], mem_q[1193:1193], mem_q[1194:1194], mem_q[1195:1195], mem_q[1196:1196], mem_q[1197:1197], mem_q[1198:1198], mem_q[1199:1199], mem_q[1200:1200], mem_q[1201:1201], mem_q[1202:1202], mem_q[1203:1203], mem_q[1204:1204], mem_q[1205:1205], mem_q[1206:1206], mem_q[1207:1207], mem_q[1208:1208], mem_q[1209:1209], mem_q[1210:1210], mem_q[1211:1211], mem_q[1212:1212], mem_q[1213:1213], mem_q[1214:1214], mem_q[1215:1215], mem_q[1216:1216], mem_q[1217:1217], mem_q[1218:1218], mem_q[1219:1219], mem_q[1220:1220], mem_q[1221:1221], mem_q[1222:1222], mem_q[1223:1223], mem_q[1224:1224], mem_q[1225:1225], mem_q[1226:1226], mem_q[1227:1227], mem_q[1228:1228], mem_q[1229:1229], mem_q[1230:1230], mem_q[1231:1231], mem_q[1232:1232], mem_q[1233:1233], mem_q[1234:1234], mem_q[1235:1235], mem_q[1236:1236], mem_q[1237:1237], mem_q[1238:1238], mem_q[1239:1239], mem_q[1240:1240], mem_q[1241:1241], mem_q[1242:1242], mem_q[1243:1243], mem_q[1244:1244], mem_q[1245:1245], mem_q[1246:1246], mem_q[1247:1247], mem_q[1248:1248], mem_q[1249:1249], mem_q[1250:1250], mem_q[1251:1251], mem_q[1252:1252], mem_q[1253:1253], mem_q[1254:1254], mem_q[1255:1255], mem_q[1256:1256], mem_q[1257:1257], mem_q[1258:1258], mem_q[1259:1259], mem_q[1260:1260], mem_q[1261:1261], mem_q[1262:1262], mem_q[1263:1263], mem_q[1264:1264], mem_q[1265:1265], mem_q[1266:1266], mem_q[1267:1267], mem_q[1268:1268], mem_q[1269:1269], mem_q[1270:1270], mem_q[1271:1271], mem_q[1272:1272], mem_q[1273:1273], mem_q[1274:1274], mem_q[1275:1275], mem_q[1276:1276], mem_q[1277:1277], mem_q[1278:1278], mem_q[1279:1279], mem_q[1280:1280], mem_q[1281:1281], mem_q[1282:1282], mem_q[1283:1283], mem_q[1284:1284], mem_q[1285:1285], mem_q[1286:1286], mem_q[1287:1287], mem_q[1288:1288], mem_q[1289:1289], mem_q[1290:1290], mem_q[1291:1291], mem_q[1292:1292], mem_q[1293:1293], mem_q[1294:1294], mem_q[1295:1295], mem_q[1296:1296], mem_q[1297:1297], mem_q[1298:1298], mem_q[1299:1299], mem_q[1300:1300], mem_q[1301:1301], mem_q[1302:1302], mem_q[1303:1303], mem_q[1304:1304], mem_q[1305:1305], mem_q[1306:1306], mem_q[1307:1307], mem_q[1308:1308], mem_q[1309:1309], mem_q[1310:1310], mem_q[1311:1311], mem_q[1312:1312], mem_q[1313:1313], mem_q[1314:1314], mem_q[1315:1315], mem_q[1316:1316], mem_q[1317:1317], mem_q[1318:1318], mem_q[1319:1319], mem_q[1320:1320], mem_q[1321:1321], mem_q[1322:1322], mem_q[1323:1323], mem_q[1324:1324], mem_q[1325:1325], mem_q[1326:1326], mem_q[1327:1327], mem_q[1328:1328], mem_q[1329:1329], mem_q[1330:1330], mem_q[1331:1331], mem_q[1332:1332], mem_q[1333:1333], mem_q[1334:1334], mem_q[1335:1335], mem_q[1336:1336], mem_q[1337:1337], mem_q[1338:1338], mem_q[1339:1339], mem_q[1340:1340], mem_q[1341:1341], mem_q[1342:1342], mem_q[1343:1343], mem_q[1344:1344], mem_q[1345:1345], mem_q[1346:1346], mem_q[1347:1347], mem_q[1348:1348], mem_q[1349:1349], mem_q[1350:1350], mem_q[1351:1351], mem_q[1352:1352], mem_q[1353:1353], mem_q[1354:1354], mem_q[1355:1355], mem_q[1356:1356], mem_q[1357:1357], mem_q[1358:1358], mem_q[1359:1359], mem_q[1360:1360], mem_q[1361:1361], mem_q[1362:1362], mem_q[1363:1363], mem_q[1364:1364], mem_q[1365:1365], mem_q[1366:1366], mem_q[1367:1367], mem_q[1368:1368], mem_q[1369:1369], mem_q[1370:1370], mem_q[1371:1371], mem_q[1372:1372], mem_q[1373:1373], mem_q[1374:1374], mem_q[1375:1375], mem_q[1376:1376], mem_q[1377:1377], mem_q[1378:1378], mem_q[1379:1379], mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383], mem_q[1384:1384], mem_q[1385:1385], mem_q[1386:1386], mem_q[1387:1387], mem_q[1388:1388], mem_q[1389:1389], mem_q[1390:1390], mem_q[1391:1391], mem_q[1392:1392], mem_q[1393:1393], mem_q[1394:1394], mem_q[1395:1395], mem_q[1396:1396], mem_q[1397:1397], mem_q[1398:1398], mem_q[1399:1399], mem_q[1400:1400], mem_q[1401:1401], mem_q[1402:1402], mem_q[1403:1403], mem_q[1404:1404], mem_q[1405:1405], mem_q[1406:1406], mem_q[1407:1407], mem_q[1408:1408], mem_q[1409:1409], mem_q[1410:1410], mem_q[1411:1411], mem_q[1412:1412], mem_q[1413:1413], mem_q[1414:1414], mem_q[1415:1415], mem_q[1416:1416], mem_q[1417:1417], mem_q[1418:1418], mem_q[1419:1419], mem_q[1420:1420], mem_q[1421:1421], mem_q[1422:1422], mem_q[1423:1423], mem_q[1424:1424], mem_q[1425:1425], mem_q[1426:1426], mem_q[1427:1427], mem_q[1428:1428], mem_q[1429:1429], mem_q[1430:1430], mem_q[1431:1431], mem_q[1432:1432], mem_q[1433:1433], mem_q[1434:1434], mem_q[1435:1435], mem_q[1436:1436], mem_q[1437:1437], mem_q[1438:1438], mem_q[1439:1439], mem_q[1440:1440], mem_q[1441:1441], mem_q[1442:1442], mem_q[1443:1443], mem_q[1444:1444], mem_q[1445:1445], mem_q[1446:1446], mem_q[1447:1447], mem_q[1448:1448], mem_q[1449:1449], mem_q[1450:1450], mem_q[1451:1451] } : 1'b0;
  assign N151 = N891;
  assign { N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353 } = (N152)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N2352)? { mem_q[1452:1452], mem_q[1453:1453], mem_q[1454:1454], mem_q[1455:1455], mem_q[1456:1456], mem_q[1457:1457], mem_q[1458:1458], mem_q[1459:1459], mem_q[1460:1460], mem_q[1461:1461], mem_q[1462:1462], mem_q[1463:1463], mem_q[1464:1464], mem_q[1465:1465], mem_q[1466:1466], mem_q[1467:1467], mem_q[1468:1468], mem_q[1469:1469], mem_q[1470:1470], mem_q[1471:1471], mem_q[1472:1472], mem_q[1473:1473], mem_q[1474:1474], mem_q[1475:1475], mem_q[1476:1476], mem_q[1477:1477], mem_q[1478:1478], mem_q[1479:1479], mem_q[1480:1480], mem_q[1481:1481], mem_q[1482:1482], mem_q[1483:1483], mem_q[1484:1484], mem_q[1485:1485], mem_q[1486:1486], mem_q[1487:1487], mem_q[1488:1488], mem_q[1489:1489], mem_q[1490:1490], mem_q[1491:1491], mem_q[1492:1492], mem_q[1493:1493], mem_q[1494:1494], mem_q[1495:1495], mem_q[1496:1496], mem_q[1497:1497], mem_q[1498:1498], mem_q[1499:1499], mem_q[1500:1500], mem_q[1501:1501], mem_q[1502:1502], mem_q[1503:1503], mem_q[1504:1504], mem_q[1505:1505], mem_q[1506:1506], mem_q[1507:1507], mem_q[1508:1508], mem_q[1509:1509], mem_q[1510:1510], mem_q[1511:1511], mem_q[1512:1512], mem_q[1513:1513], mem_q[1514:1514], mem_q[1515:1515], mem_q[1516:1516], mem_q[1517:1517], mem_q[1518:1518], mem_q[1519:1519], mem_q[1520:1520], mem_q[1521:1521], mem_q[1522:1522], mem_q[1523:1523], mem_q[1524:1524], mem_q[1525:1525], mem_q[1526:1526], mem_q[1527:1527], mem_q[1528:1528], mem_q[1529:1529], mem_q[1530:1530], mem_q[1531:1531], mem_q[1532:1532], mem_q[1533:1533], mem_q[1534:1534], mem_q[1535:1535], mem_q[1536:1536], mem_q[1537:1537], mem_q[1538:1538], mem_q[1539:1539], mem_q[1540:1540], mem_q[1541:1541], mem_q[1542:1542], mem_q[1543:1543], mem_q[1544:1544], mem_q[1545:1545], mem_q[1546:1546], mem_q[1547:1547], mem_q[1548:1548], mem_q[1549:1549], mem_q[1550:1550], mem_q[1551:1551], mem_q[1552:1552], mem_q[1553:1553], mem_q[1554:1554], mem_q[1555:1555], mem_q[1556:1556], mem_q[1557:1557], mem_q[1558:1558], mem_q[1559:1559], mem_q[1560:1560], mem_q[1561:1561], mem_q[1562:1562], mem_q[1563:1563], mem_q[1564:1564], mem_q[1565:1565], mem_q[1566:1566], mem_q[1567:1567], mem_q[1568:1568], mem_q[1569:1569], mem_q[1570:1570], mem_q[1571:1571], mem_q[1572:1572], mem_q[1573:1573], mem_q[1574:1574], mem_q[1575:1575], mem_q[1576:1576], mem_q[1577:1577], mem_q[1578:1578], mem_q[1579:1579], mem_q[1580:1580], mem_q[1581:1581], mem_q[1582:1582], mem_q[1583:1583], mem_q[1584:1584], mem_q[1585:1585], mem_q[1586:1586], mem_q[1587:1587], mem_q[1588:1588], mem_q[1589:1589], mem_q[1590:1590], mem_q[1591:1591], mem_q[1592:1592], mem_q[1593:1593], mem_q[1594:1594], mem_q[1595:1595], mem_q[1596:1596], mem_q[1597:1597], mem_q[1598:1598], mem_q[1599:1599], mem_q[1600:1600], mem_q[1601:1601], mem_q[1602:1602], mem_q[1603:1603], mem_q[1604:1604], mem_q[1605:1605], mem_q[1606:1606], mem_q[1607:1607], mem_q[1608:1608], mem_q[1609:1609], mem_q[1610:1610], mem_q[1611:1611], mem_q[1612:1612], mem_q[1613:1613], mem_q[1614:1614], mem_q[1615:1615], mem_q[1616:1616], mem_q[1617:1617], mem_q[1618:1618], mem_q[1619:1619], mem_q[1620:1620], mem_q[1621:1621], mem_q[1622:1622], mem_q[1623:1623], mem_q[1624:1624], mem_q[1625:1625], mem_q[1626:1626], mem_q[1627:1627], mem_q[1628:1628], mem_q[1629:1629], mem_q[1630:1630], mem_q[1631:1631], mem_q[1632:1632], mem_q[1633:1633], mem_q[1634:1634], mem_q[1635:1635], mem_q[1636:1636], mem_q[1637:1637], mem_q[1638:1638], mem_q[1639:1639], mem_q[1640:1640], mem_q[1641:1641], mem_q[1642:1642], mem_q[1643:1643], mem_q[1644:1644], mem_q[1645:1645], mem_q[1646:1646], mem_q[1647:1647], mem_q[1648:1648], mem_q[1649:1649], mem_q[1650:1650], mem_q[1651:1651], mem_q[1652:1652], mem_q[1653:1653], mem_q[1654:1654], mem_q[1655:1655], mem_q[1656:1656], mem_q[1657:1657], mem_q[1658:1658], mem_q[1659:1659], mem_q[1660:1660], mem_q[1661:1661], mem_q[1662:1662], mem_q[1663:1663], mem_q[1664:1664], mem_q[1665:1665], mem_q[1666:1666], mem_q[1667:1667], mem_q[1668:1668], mem_q[1669:1669], mem_q[1670:1670], mem_q[1671:1671], mem_q[1672:1672], mem_q[1673:1673], mem_q[1674:1674], mem_q[1675:1675], mem_q[1676:1676], mem_q[1677:1677], mem_q[1678:1678], mem_q[1679:1679], mem_q[1680:1680], mem_q[1681:1681], mem_q[1682:1682], mem_q[1683:1683], mem_q[1684:1684], mem_q[1685:1685], mem_q[1686:1686], mem_q[1687:1687], mem_q[1688:1688], mem_q[1689:1689], mem_q[1690:1690], mem_q[1691:1691], mem_q[1692:1692], mem_q[1693:1693], mem_q[1694:1694], mem_q[1695:1695], mem_q[1696:1696], mem_q[1697:1697], mem_q[1698:1698], mem_q[1699:1699], mem_q[1700:1700], mem_q[1701:1701], mem_q[1702:1702], mem_q[1703:1703], mem_q[1704:1704], mem_q[1705:1705], mem_q[1706:1706], mem_q[1707:1707], mem_q[1708:1708], mem_q[1709:1709], mem_q[1710:1710], mem_q[1711:1711], mem_q[1712:1712], mem_q[1713:1713], mem_q[1714:1714], mem_q[1715:1715], mem_q[1716:1716], mem_q[1717:1717], mem_q[1718:1718], mem_q[1719:1719], mem_q[1720:1720], mem_q[1721:1721], mem_q[1722:1722], mem_q[1723:1723], mem_q[1724:1724], mem_q[1725:1725], mem_q[1726:1726], mem_q[1727:1727], mem_q[1728:1728], mem_q[1729:1729], mem_q[1730:1730], mem_q[1731:1731], mem_q[1732:1732], mem_q[1733:1733], mem_q[1734:1734], mem_q[1735:1735], mem_q[1736:1736], mem_q[1737:1737], mem_q[1738:1738], mem_q[1739:1739], mem_q[1740:1740], mem_q[1741:1741], mem_q[1742:1742], mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746], mem_q[1747:1747], mem_q[1748:1748], mem_q[1749:1749], mem_q[1750:1750], mem_q[1751:1751], mem_q[1752:1752], mem_q[1753:1753], mem_q[1754:1754], mem_q[1755:1755], mem_q[1756:1756], mem_q[1757:1757], mem_q[1758:1758], mem_q[1759:1759], mem_q[1760:1760], mem_q[1761:1761], mem_q[1762:1762], mem_q[1763:1763], mem_q[1764:1764], mem_q[1765:1765], mem_q[1766:1766], mem_q[1767:1767], mem_q[1768:1768], mem_q[1769:1769], mem_q[1770:1770], mem_q[1771:1771], mem_q[1772:1772], mem_q[1773:1773], mem_q[1774:1774], mem_q[1775:1775], mem_q[1776:1776], mem_q[1777:1777], mem_q[1778:1778], mem_q[1779:1779], mem_q[1780:1780], mem_q[1781:1781], mem_q[1782:1782], mem_q[1783:1783], mem_q[1784:1784], mem_q[1785:1785], mem_q[1786:1786], mem_q[1787:1787], mem_q[1788:1788], mem_q[1789:1789], mem_q[1790:1790], mem_q[1791:1791], mem_q[1792:1792], mem_q[1793:1793], mem_q[1794:1794], mem_q[1795:1795], mem_q[1796:1796], mem_q[1797:1797], mem_q[1798:1798], mem_q[1799:1799], mem_q[1800:1800], mem_q[1801:1801], mem_q[1802:1802], mem_q[1803:1803], mem_q[1804:1804], mem_q[1805:1805], mem_q[1806:1806], mem_q[1807:1807], mem_q[1808:1808], mem_q[1809:1809], mem_q[1810:1810], mem_q[1811:1811], mem_q[1812:1812], mem_q[1813:1813], mem_q[1814:1814] } : 1'b0;
  assign N152 = N892;
  assign { N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717 } = (N153)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N2716)? { mem_q[1815:1815], mem_q[1816:1816], mem_q[1817:1817], mem_q[1818:1818], mem_q[1819:1819], mem_q[1820:1820], mem_q[1821:1821], mem_q[1822:1822], mem_q[1823:1823], mem_q[1824:1824], mem_q[1825:1825], mem_q[1826:1826], mem_q[1827:1827], mem_q[1828:1828], mem_q[1829:1829], mem_q[1830:1830], mem_q[1831:1831], mem_q[1832:1832], mem_q[1833:1833], mem_q[1834:1834], mem_q[1835:1835], mem_q[1836:1836], mem_q[1837:1837], mem_q[1838:1838], mem_q[1839:1839], mem_q[1840:1840], mem_q[1841:1841], mem_q[1842:1842], mem_q[1843:1843], mem_q[1844:1844], mem_q[1845:1845], mem_q[1846:1846], mem_q[1847:1847], mem_q[1848:1848], mem_q[1849:1849], mem_q[1850:1850], mem_q[1851:1851], mem_q[1852:1852], mem_q[1853:1853], mem_q[1854:1854], mem_q[1855:1855], mem_q[1856:1856], mem_q[1857:1857], mem_q[1858:1858], mem_q[1859:1859], mem_q[1860:1860], mem_q[1861:1861], mem_q[1862:1862], mem_q[1863:1863], mem_q[1864:1864], mem_q[1865:1865], mem_q[1866:1866], mem_q[1867:1867], mem_q[1868:1868], mem_q[1869:1869], mem_q[1870:1870], mem_q[1871:1871], mem_q[1872:1872], mem_q[1873:1873], mem_q[1874:1874], mem_q[1875:1875], mem_q[1876:1876], mem_q[1877:1877], mem_q[1878:1878], mem_q[1879:1879], mem_q[1880:1880], mem_q[1881:1881], mem_q[1882:1882], mem_q[1883:1883], mem_q[1884:1884], mem_q[1885:1885], mem_q[1886:1886], mem_q[1887:1887], mem_q[1888:1888], mem_q[1889:1889], mem_q[1890:1890], mem_q[1891:1891], mem_q[1892:1892], mem_q[1893:1893], mem_q[1894:1894], mem_q[1895:1895], mem_q[1896:1896], mem_q[1897:1897], mem_q[1898:1898], mem_q[1899:1899], mem_q[1900:1900], mem_q[1901:1901], mem_q[1902:1902], mem_q[1903:1903], mem_q[1904:1904], mem_q[1905:1905], mem_q[1906:1906], mem_q[1907:1907], mem_q[1908:1908], mem_q[1909:1909], mem_q[1910:1910], mem_q[1911:1911], mem_q[1912:1912], mem_q[1913:1913], mem_q[1914:1914], mem_q[1915:1915], mem_q[1916:1916], mem_q[1917:1917], mem_q[1918:1918], mem_q[1919:1919], mem_q[1920:1920], mem_q[1921:1921], mem_q[1922:1922], mem_q[1923:1923], mem_q[1924:1924], mem_q[1925:1925], mem_q[1926:1926], mem_q[1927:1927], mem_q[1928:1928], mem_q[1929:1929], mem_q[1930:1930], mem_q[1931:1931], mem_q[1932:1932], mem_q[1933:1933], mem_q[1934:1934], mem_q[1935:1935], mem_q[1936:1936], mem_q[1937:1937], mem_q[1938:1938], mem_q[1939:1939], mem_q[1940:1940], mem_q[1941:1941], mem_q[1942:1942], mem_q[1943:1943], mem_q[1944:1944], mem_q[1945:1945], mem_q[1946:1946], mem_q[1947:1947], mem_q[1948:1948], mem_q[1949:1949], mem_q[1950:1950], mem_q[1951:1951], mem_q[1952:1952], mem_q[1953:1953], mem_q[1954:1954], mem_q[1955:1955], mem_q[1956:1956], mem_q[1957:1957], mem_q[1958:1958], mem_q[1959:1959], mem_q[1960:1960], mem_q[1961:1961], mem_q[1962:1962], mem_q[1963:1963], mem_q[1964:1964], mem_q[1965:1965], mem_q[1966:1966], mem_q[1967:1967], mem_q[1968:1968], mem_q[1969:1969], mem_q[1970:1970], mem_q[1971:1971], mem_q[1972:1972], mem_q[1973:1973], mem_q[1974:1974], mem_q[1975:1975], mem_q[1976:1976], mem_q[1977:1977], mem_q[1978:1978], mem_q[1979:1979], mem_q[1980:1980], mem_q[1981:1981], mem_q[1982:1982], mem_q[1983:1983], mem_q[1984:1984], mem_q[1985:1985], mem_q[1986:1986], mem_q[1987:1987], mem_q[1988:1988], mem_q[1989:1989], mem_q[1990:1990], mem_q[1991:1991], mem_q[1992:1992], mem_q[1993:1993], mem_q[1994:1994], mem_q[1995:1995], mem_q[1996:1996], mem_q[1997:1997], mem_q[1998:1998], mem_q[1999:1999], mem_q[2000:2000], mem_q[2001:2001], mem_q[2002:2002], mem_q[2003:2003], mem_q[2004:2004], mem_q[2005:2005], mem_q[2006:2006], mem_q[2007:2007], mem_q[2008:2008], mem_q[2009:2009], mem_q[2010:2010], mem_q[2011:2011], mem_q[2012:2012], mem_q[2013:2013], mem_q[2014:2014], mem_q[2015:2015], mem_q[2016:2016], mem_q[2017:2017], mem_q[2018:2018], mem_q[2019:2019], mem_q[2020:2020], mem_q[2021:2021], mem_q[2022:2022], mem_q[2023:2023], mem_q[2024:2024], mem_q[2025:2025], mem_q[2026:2026], mem_q[2027:2027], mem_q[2028:2028], mem_q[2029:2029], mem_q[2030:2030], mem_q[2031:2031], mem_q[2032:2032], mem_q[2033:2033], mem_q[2034:2034], mem_q[2035:2035], mem_q[2036:2036], mem_q[2037:2037], mem_q[2038:2038], mem_q[2039:2039], mem_q[2040:2040], mem_q[2041:2041], mem_q[2042:2042], mem_q[2043:2043], mem_q[2044:2044], mem_q[2045:2045], mem_q[2046:2046], mem_q[2047:2047], mem_q[2048:2048], mem_q[2049:2049], mem_q[2050:2050], mem_q[2051:2051], mem_q[2052:2052], mem_q[2053:2053], mem_q[2054:2054], mem_q[2055:2055], mem_q[2056:2056], mem_q[2057:2057], mem_q[2058:2058], mem_q[2059:2059], mem_q[2060:2060], mem_q[2061:2061], mem_q[2062:2062], mem_q[2063:2063], mem_q[2064:2064], mem_q[2065:2065], mem_q[2066:2066], mem_q[2067:2067], mem_q[2068:2068], mem_q[2069:2069], mem_q[2070:2070], mem_q[2071:2071], mem_q[2072:2072], mem_q[2073:2073], mem_q[2074:2074], mem_q[2075:2075], mem_q[2076:2076], mem_q[2077:2077], mem_q[2078:2078], mem_q[2079:2079], mem_q[2080:2080], mem_q[2081:2081], mem_q[2082:2082], mem_q[2083:2083], mem_q[2084:2084], mem_q[2085:2085], mem_q[2086:2086], mem_q[2087:2087], mem_q[2088:2088], mem_q[2089:2089], mem_q[2090:2090], mem_q[2091:2091], mem_q[2092:2092], mem_q[2093:2093], mem_q[2094:2094], mem_q[2095:2095], mem_q[2096:2096], mem_q[2097:2097], mem_q[2098:2098], mem_q[2099:2099], mem_q[2100:2100], mem_q[2101:2101], mem_q[2102:2102], mem_q[2103:2103], mem_q[2104:2104], mem_q[2105:2105], mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109], mem_q[2110:2110], mem_q[2111:2111], mem_q[2112:2112], mem_q[2113:2113], mem_q[2114:2114], mem_q[2115:2115], mem_q[2116:2116], mem_q[2117:2117], mem_q[2118:2118], mem_q[2119:2119], mem_q[2120:2120], mem_q[2121:2121], mem_q[2122:2122], mem_q[2123:2123], mem_q[2124:2124], mem_q[2125:2125], mem_q[2126:2126], mem_q[2127:2127], mem_q[2128:2128], mem_q[2129:2129], mem_q[2130:2130], mem_q[2131:2131], mem_q[2132:2132], mem_q[2133:2133], mem_q[2134:2134], mem_q[2135:2135], mem_q[2136:2136], mem_q[2137:2137], mem_q[2138:2138], mem_q[2139:2139], mem_q[2140:2140], mem_q[2141:2141], mem_q[2142:2142], mem_q[2143:2143], mem_q[2144:2144], mem_q[2145:2145], mem_q[2146:2146], mem_q[2147:2147], mem_q[2148:2148], mem_q[2149:2149], mem_q[2150:2150], mem_q[2151:2151], mem_q[2152:2152], mem_q[2153:2153], mem_q[2154:2154], mem_q[2155:2155], mem_q[2156:2156], mem_q[2157:2157], mem_q[2158:2158], mem_q[2159:2159], mem_q[2160:2160], mem_q[2161:2161], mem_q[2162:2162], mem_q[2163:2163], mem_q[2164:2164], mem_q[2165:2165], mem_q[2166:2166], mem_q[2167:2167], mem_q[2168:2168], mem_q[2169:2169], mem_q[2170:2170], mem_q[2171:2171], mem_q[2172:2172], mem_q[2173:2173], mem_q[2174:2174], mem_q[2175:2175], mem_q[2176:2176], mem_q[2177:2177] } : 1'b0;
  assign N153 = N893;
  assign { N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251, N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N3226, N3225, N3224, N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081 } = (N154)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N3080)? { mem_q[2178:2178], mem_q[2179:2179], mem_q[2180:2180], mem_q[2181:2181], mem_q[2182:2182], mem_q[2183:2183], mem_q[2184:2184], mem_q[2185:2185], mem_q[2186:2186], mem_q[2187:2187], mem_q[2188:2188], mem_q[2189:2189], mem_q[2190:2190], mem_q[2191:2191], mem_q[2192:2192], mem_q[2193:2193], mem_q[2194:2194], mem_q[2195:2195], mem_q[2196:2196], mem_q[2197:2197], mem_q[2198:2198], mem_q[2199:2199], mem_q[2200:2200], mem_q[2201:2201], mem_q[2202:2202], mem_q[2203:2203], mem_q[2204:2204], mem_q[2205:2205], mem_q[2206:2206], mem_q[2207:2207], mem_q[2208:2208], mem_q[2209:2209], mem_q[2210:2210], mem_q[2211:2211], mem_q[2212:2212], mem_q[2213:2213], mem_q[2214:2214], mem_q[2215:2215], mem_q[2216:2216], mem_q[2217:2217], mem_q[2218:2218], mem_q[2219:2219], mem_q[2220:2220], mem_q[2221:2221], mem_q[2222:2222], mem_q[2223:2223], mem_q[2224:2224], mem_q[2225:2225], mem_q[2226:2226], mem_q[2227:2227], mem_q[2228:2228], mem_q[2229:2229], mem_q[2230:2230], mem_q[2231:2231], mem_q[2232:2232], mem_q[2233:2233], mem_q[2234:2234], mem_q[2235:2235], mem_q[2236:2236], mem_q[2237:2237], mem_q[2238:2238], mem_q[2239:2239], mem_q[2240:2240], mem_q[2241:2241], mem_q[2242:2242], mem_q[2243:2243], mem_q[2244:2244], mem_q[2245:2245], mem_q[2246:2246], mem_q[2247:2247], mem_q[2248:2248], mem_q[2249:2249], mem_q[2250:2250], mem_q[2251:2251], mem_q[2252:2252], mem_q[2253:2253], mem_q[2254:2254], mem_q[2255:2255], mem_q[2256:2256], mem_q[2257:2257], mem_q[2258:2258], mem_q[2259:2259], mem_q[2260:2260], mem_q[2261:2261], mem_q[2262:2262], mem_q[2263:2263], mem_q[2264:2264], mem_q[2265:2265], mem_q[2266:2266], mem_q[2267:2267], mem_q[2268:2268], mem_q[2269:2269], mem_q[2270:2270], mem_q[2271:2271], mem_q[2272:2272], mem_q[2273:2273], mem_q[2274:2274], mem_q[2275:2275], mem_q[2276:2276], mem_q[2277:2277], mem_q[2278:2278], mem_q[2279:2279], mem_q[2280:2280], mem_q[2281:2281], mem_q[2282:2282], mem_q[2283:2283], mem_q[2284:2284], mem_q[2285:2285], mem_q[2286:2286], mem_q[2287:2287], mem_q[2288:2288], mem_q[2289:2289], mem_q[2290:2290], mem_q[2291:2291], mem_q[2292:2292], mem_q[2293:2293], mem_q[2294:2294], mem_q[2295:2295], mem_q[2296:2296], mem_q[2297:2297], mem_q[2298:2298], mem_q[2299:2299], mem_q[2300:2300], mem_q[2301:2301], mem_q[2302:2302], mem_q[2303:2303], mem_q[2304:2304], mem_q[2305:2305], mem_q[2306:2306], mem_q[2307:2307], mem_q[2308:2308], mem_q[2309:2309], mem_q[2310:2310], mem_q[2311:2311], mem_q[2312:2312], mem_q[2313:2313], mem_q[2314:2314], mem_q[2315:2315], mem_q[2316:2316], mem_q[2317:2317], mem_q[2318:2318], mem_q[2319:2319], mem_q[2320:2320], mem_q[2321:2321], mem_q[2322:2322], mem_q[2323:2323], mem_q[2324:2324], mem_q[2325:2325], mem_q[2326:2326], mem_q[2327:2327], mem_q[2328:2328], mem_q[2329:2329], mem_q[2330:2330], mem_q[2331:2331], mem_q[2332:2332], mem_q[2333:2333], mem_q[2334:2334], mem_q[2335:2335], mem_q[2336:2336], mem_q[2337:2337], mem_q[2338:2338], mem_q[2339:2339], mem_q[2340:2340], mem_q[2341:2341], mem_q[2342:2342], mem_q[2343:2343], mem_q[2344:2344], mem_q[2345:2345], mem_q[2346:2346], mem_q[2347:2347], mem_q[2348:2348], mem_q[2349:2349], mem_q[2350:2350], mem_q[2351:2351], mem_q[2352:2352], mem_q[2353:2353], mem_q[2354:2354], mem_q[2355:2355], mem_q[2356:2356], mem_q[2357:2357], mem_q[2358:2358], mem_q[2359:2359], mem_q[2360:2360], mem_q[2361:2361], mem_q[2362:2362], mem_q[2363:2363], mem_q[2364:2364], mem_q[2365:2365], mem_q[2366:2366], mem_q[2367:2367], mem_q[2368:2368], mem_q[2369:2369], mem_q[2370:2370], mem_q[2371:2371], mem_q[2372:2372], mem_q[2373:2373], mem_q[2374:2374], mem_q[2375:2375], mem_q[2376:2376], mem_q[2377:2377], mem_q[2378:2378], mem_q[2379:2379], mem_q[2380:2380], mem_q[2381:2381], mem_q[2382:2382], mem_q[2383:2383], mem_q[2384:2384], mem_q[2385:2385], mem_q[2386:2386], mem_q[2387:2387], mem_q[2388:2388], mem_q[2389:2389], mem_q[2390:2390], mem_q[2391:2391], mem_q[2392:2392], mem_q[2393:2393], mem_q[2394:2394], mem_q[2395:2395], mem_q[2396:2396], mem_q[2397:2397], mem_q[2398:2398], mem_q[2399:2399], mem_q[2400:2400], mem_q[2401:2401], mem_q[2402:2402], mem_q[2403:2403], mem_q[2404:2404], mem_q[2405:2405], mem_q[2406:2406], mem_q[2407:2407], mem_q[2408:2408], mem_q[2409:2409], mem_q[2410:2410], mem_q[2411:2411], mem_q[2412:2412], mem_q[2413:2413], mem_q[2414:2414], mem_q[2415:2415], mem_q[2416:2416], mem_q[2417:2417], mem_q[2418:2418], mem_q[2419:2419], mem_q[2420:2420], mem_q[2421:2421], mem_q[2422:2422], mem_q[2423:2423], mem_q[2424:2424], mem_q[2425:2425], mem_q[2426:2426], mem_q[2427:2427], mem_q[2428:2428], mem_q[2429:2429], mem_q[2430:2430], mem_q[2431:2431], mem_q[2432:2432], mem_q[2433:2433], mem_q[2434:2434], mem_q[2435:2435], mem_q[2436:2436], mem_q[2437:2437], mem_q[2438:2438], mem_q[2439:2439], mem_q[2440:2440], mem_q[2441:2441], mem_q[2442:2442], mem_q[2443:2443], mem_q[2444:2444], mem_q[2445:2445], mem_q[2446:2446], mem_q[2447:2447], mem_q[2448:2448], mem_q[2449:2449], mem_q[2450:2450], mem_q[2451:2451], mem_q[2452:2452], mem_q[2453:2453], mem_q[2454:2454], mem_q[2455:2455], mem_q[2456:2456], mem_q[2457:2457], mem_q[2458:2458], mem_q[2459:2459], mem_q[2460:2460], mem_q[2461:2461], mem_q[2462:2462], mem_q[2463:2463], mem_q[2464:2464], mem_q[2465:2465], mem_q[2466:2466], mem_q[2467:2467], mem_q[2468:2468], mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472], mem_q[2473:2473], mem_q[2474:2474], mem_q[2475:2475], mem_q[2476:2476], mem_q[2477:2477], mem_q[2478:2478], mem_q[2479:2479], mem_q[2480:2480], mem_q[2481:2481], mem_q[2482:2482], mem_q[2483:2483], mem_q[2484:2484], mem_q[2485:2485], mem_q[2486:2486], mem_q[2487:2487], mem_q[2488:2488], mem_q[2489:2489], mem_q[2490:2490], mem_q[2491:2491], mem_q[2492:2492], mem_q[2493:2493], mem_q[2494:2494], mem_q[2495:2495], mem_q[2496:2496], mem_q[2497:2497], mem_q[2498:2498], mem_q[2499:2499], mem_q[2500:2500], mem_q[2501:2501], mem_q[2502:2502], mem_q[2503:2503], mem_q[2504:2504], mem_q[2505:2505], mem_q[2506:2506], mem_q[2507:2507], mem_q[2508:2508], mem_q[2509:2509], mem_q[2510:2510], mem_q[2511:2511], mem_q[2512:2512], mem_q[2513:2513], mem_q[2514:2514], mem_q[2515:2515], mem_q[2516:2516], mem_q[2517:2517], mem_q[2518:2518], mem_q[2519:2519], mem_q[2520:2520], mem_q[2521:2521], mem_q[2522:2522], mem_q[2523:2523], mem_q[2524:2524], mem_q[2525:2525], mem_q[2526:2526], mem_q[2527:2527], mem_q[2528:2528], mem_q[2529:2529], mem_q[2530:2530], mem_q[2531:2531], mem_q[2532:2532], mem_q[2533:2533], mem_q[2534:2534], mem_q[2535:2535], mem_q[2536:2536], mem_q[2537:2537], mem_q[2538:2538], mem_q[2539:2539], mem_q[2540:2540] } : 1'b0;
  assign N154 = N894;
  assign { N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445 } = (N155)? { decoded_instr_i[0:0], decoded_instr_i[1:1], decoded_instr_i[2:2], decoded_instr_i[3:3], decoded_instr_i[4:4], decoded_instr_i[5:5], decoded_instr_i[6:6], decoded_instr_i[7:7], decoded_instr_i[8:8], decoded_instr_i[9:9], decoded_instr_i[10:10], decoded_instr_i[11:11], decoded_instr_i[12:12], decoded_instr_i[13:13], decoded_instr_i[14:14], decoded_instr_i[15:15], decoded_instr_i[16:16], decoded_instr_i[17:17], decoded_instr_i[18:18], decoded_instr_i[19:19], decoded_instr_i[20:20], decoded_instr_i[21:21], decoded_instr_i[22:22], decoded_instr_i[23:23], decoded_instr_i[24:24], decoded_instr_i[25:25], decoded_instr_i[26:26], decoded_instr_i[27:27], decoded_instr_i[28:28], decoded_instr_i[29:29], decoded_instr_i[30:30], decoded_instr_i[31:31], decoded_instr_i[32:32], decoded_instr_i[33:33], decoded_instr_i[34:34], decoded_instr_i[35:35], decoded_instr_i[36:36], decoded_instr_i[37:37], decoded_instr_i[38:38], decoded_instr_i[39:39], decoded_instr_i[40:40], decoded_instr_i[41:41], decoded_instr_i[42:42], decoded_instr_i[43:43], decoded_instr_i[44:44], decoded_instr_i[45:45], decoded_instr_i[46:46], decoded_instr_i[47:47], decoded_instr_i[48:48], decoded_instr_i[49:49], decoded_instr_i[50:50], decoded_instr_i[51:51], decoded_instr_i[52:52], decoded_instr_i[53:53], decoded_instr_i[54:54], decoded_instr_i[55:55], decoded_instr_i[56:56], decoded_instr_i[57:57], decoded_instr_i[58:58], decoded_instr_i[59:59], decoded_instr_i[60:60], decoded_instr_i[61:61], decoded_instr_i[62:62], decoded_instr_i[63:63], decoded_instr_i[64:64], decoded_instr_i[65:65], decoded_instr_i[66:66], decoded_instr_i[67:67], decoded_instr_i[68:68], decoded_instr_i[69:69], decoded_instr_i[70:70], decoded_instr_i[71:71], decoded_instr_i[72:72], decoded_instr_i[73:73], decoded_instr_i[74:74], decoded_instr_i[75:75], decoded_instr_i[76:76], decoded_instr_i[77:77], decoded_instr_i[78:78], decoded_instr_i[79:79], decoded_instr_i[80:80], decoded_instr_i[81:81], decoded_instr_i[82:82], decoded_instr_i[83:83], decoded_instr_i[84:84], decoded_instr_i[85:85], decoded_instr_i[86:86], decoded_instr_i[87:87], decoded_instr_i[88:88], decoded_instr_i[89:89], decoded_instr_i[90:90], decoded_instr_i[91:91], decoded_instr_i[92:92], decoded_instr_i[93:93], decoded_instr_i[94:94], decoded_instr_i[95:95], decoded_instr_i[96:96], decoded_instr_i[97:97], decoded_instr_i[98:98], decoded_instr_i[99:99], decoded_instr_i[100:100], decoded_instr_i[101:101], decoded_instr_i[102:102], decoded_instr_i[103:103], decoded_instr_i[104:104], decoded_instr_i[105:105], decoded_instr_i[106:106], decoded_instr_i[107:107], decoded_instr_i[108:108], decoded_instr_i[109:109], decoded_instr_i[110:110], decoded_instr_i[111:111], decoded_instr_i[112:112], decoded_instr_i[113:113], decoded_instr_i[114:114], decoded_instr_i[115:115], decoded_instr_i[116:116], decoded_instr_i[117:117], decoded_instr_i[118:118], decoded_instr_i[119:119], decoded_instr_i[120:120], decoded_instr_i[121:121], decoded_instr_i[122:122], decoded_instr_i[123:123], decoded_instr_i[124:124], decoded_instr_i[125:125], decoded_instr_i[126:126], decoded_instr_i[127:127], decoded_instr_i[128:128], decoded_instr_i[129:129], decoded_instr_i[130:130], decoded_instr_i[131:131], decoded_instr_i[132:132], decoded_instr_i[133:133], decoded_instr_i[134:134], decoded_instr_i[135:135], decoded_instr_i[136:136], decoded_instr_i[137:137], decoded_instr_i[138:138], decoded_instr_i[139:139], decoded_instr_i[140:140], decoded_instr_i[141:141], decoded_instr_i[142:142], decoded_instr_i[143:143], decoded_instr_i[144:144], decoded_instr_i[145:145], decoded_instr_i[146:146], decoded_instr_i[147:147], decoded_instr_i[148:148], decoded_instr_i[149:149], decoded_instr_i[150:150], decoded_instr_i[151:151], decoded_instr_i[152:152], decoded_instr_i[153:153], decoded_instr_i[154:154], decoded_instr_i[155:155], decoded_instr_i[156:156], decoded_instr_i[157:157], decoded_instr_i[158:158], decoded_instr_i[159:159], decoded_instr_i[160:160], decoded_instr_i[161:161], decoded_instr_i[162:162], decoded_instr_i[163:163], decoded_instr_i[164:164], decoded_instr_i[165:165], decoded_instr_i[166:166], decoded_instr_i[167:167], decoded_instr_i[168:168], decoded_instr_i[169:169], decoded_instr_i[170:170], decoded_instr_i[171:171], decoded_instr_i[172:172], decoded_instr_i[173:173], decoded_instr_i[174:174], decoded_instr_i[175:175], decoded_instr_i[176:176], decoded_instr_i[177:177], decoded_instr_i[178:178], decoded_instr_i[179:179], decoded_instr_i[180:180], decoded_instr_i[181:181], decoded_instr_i[182:182], decoded_instr_i[183:183], decoded_instr_i[184:184], decoded_instr_i[185:185], decoded_instr_i[186:186], decoded_instr_i[187:187], decoded_instr_i[188:188], decoded_instr_i[189:189], decoded_instr_i[190:190], decoded_instr_i[191:191], decoded_instr_i[192:192], decoded_instr_i[193:193], decoded_instr_i[194:194], decoded_instr_i[195:195], decoded_instr_i[196:196], decoded_instr_i[197:197], decoded_instr_i[198:198], decoded_instr_i[199:199], decoded_instr_i[200:200], decoded_instr_i[201:201], decoded_instr_i[202:202], decoded_instr_i[203:203], decoded_instr_i[204:204], decoded_instr_i[205:205], decoded_instr_i[206:206], decoded_instr_i[207:207], decoded_instr_i[208:208], decoded_instr_i[209:209], decoded_instr_i[210:210], decoded_instr_i[211:211], decoded_instr_i[212:212], decoded_instr_i[213:213], decoded_instr_i[214:214], decoded_instr_i[215:215], decoded_instr_i[216:216], decoded_instr_i[217:217], decoded_instr_i[218:218], decoded_instr_i[219:219], decoded_instr_i[220:220], decoded_instr_i[221:221], decoded_instr_i[222:222], decoded_instr_i[223:223], decoded_instr_i[224:224], decoded_instr_i[225:225], decoded_instr_i[226:226], decoded_instr_i[227:227], decoded_instr_i[228:228], decoded_instr_i[229:229], decoded_instr_i[230:230], decoded_instr_i[231:231], decoded_instr_i[232:232], decoded_instr_i[233:233], decoded_instr_i[234:234], decoded_instr_i[235:235], decoded_instr_i[236:236], decoded_instr_i[237:237], decoded_instr_i[238:238], decoded_instr_i[239:239], decoded_instr_i[240:240], decoded_instr_i[241:241], decoded_instr_i[242:242], decoded_instr_i[243:243], decoded_instr_i[244:244], decoded_instr_i[245:245], decoded_instr_i[246:246], decoded_instr_i[247:247], decoded_instr_i[248:248], decoded_instr_i[249:249], decoded_instr_i[250:250], decoded_instr_i[251:251], decoded_instr_i[252:252], decoded_instr_i[253:253], decoded_instr_i[254:254], decoded_instr_i[255:255], decoded_instr_i[256:256], decoded_instr_i[257:257], decoded_instr_i[258:258], decoded_instr_i[259:259], decoded_instr_i[260:260], decoded_instr_i[261:261], decoded_instr_i[262:262], decoded_instr_i[263:263], decoded_instr_i[264:264], decoded_instr_i[265:265], decoded_instr_i[266:266], decoded_instr_i[267:267], decoded_instr_i[268:268], decoded_instr_i[269:269], decoded_instr_i[270:270], decoded_instr_i[271:271], decoded_instr_i[272:272], decoded_instr_i[273:273], decoded_instr_i[274:274], decoded_instr_i[275:275], decoded_instr_i[276:276], decoded_instr_i[277:277], decoded_instr_i[278:278], decoded_instr_i[279:279], decoded_instr_i[280:280], decoded_instr_i[281:281], decoded_instr_i[282:282], decoded_instr_i[283:283], decoded_instr_i[284:284], decoded_instr_i[285:285], decoded_instr_i[286:286], decoded_instr_i[287:287], decoded_instr_i[288:288], decoded_instr_i[289:289], decoded_instr_i[290:290], decoded_instr_i[291:291], decoded_instr_i[292:292], decoded_instr_i[293:293], decoded_instr_i[294:294], decoded_instr_i[295:295], decoded_instr_i[296:296], decoded_instr_i[297:297], decoded_instr_i[298:298], decoded_instr_i[299:299], decoded_instr_i[300:300], decoded_instr_i[301:301], decoded_instr_i[302:302], decoded_instr_i[303:303], decoded_instr_i[304:304], decoded_instr_i[305:305], decoded_instr_i[306:306], decoded_instr_i[307:307], decoded_instr_i[308:308], decoded_instr_i[309:309], decoded_instr_i[310:310], decoded_instr_i[311:311], decoded_instr_i[312:312], decoded_instr_i[313:313], decoded_instr_i[314:314], decoded_instr_i[315:315], decoded_instr_i[316:316], decoded_instr_i[317:317], decoded_instr_i[318:318], decoded_instr_i[319:319], decoded_instr_i[320:320], decoded_instr_i[321:321], decoded_instr_i[322:322], decoded_instr_i[323:323], decoded_instr_i[324:324], decoded_instr_i[325:325], decoded_instr_i[326:326], decoded_instr_i[327:327], decoded_instr_i[328:328], decoded_instr_i[329:329], decoded_instr_i[330:330], decoded_instr_i[331:331], decoded_instr_i[332:332], decoded_instr_i[333:333], decoded_instr_i[334:334], decoded_instr_i[335:335], decoded_instr_i[336:336], decoded_instr_i[337:337], decoded_instr_i[338:338], decoded_instr_i[339:339], decoded_instr_i[340:340], decoded_instr_i[341:341], decoded_instr_i[342:342], decoded_instr_i[343:343], decoded_instr_i[344:344], decoded_instr_i[345:345], decoded_instr_i[346:346], decoded_instr_i[347:347], decoded_instr_i[348:348], decoded_instr_i[349:349], decoded_instr_i[350:350], decoded_instr_i[351:351], decoded_instr_i[352:352], decoded_instr_i[353:353], decoded_instr_i[354:354], decoded_instr_i[355:355], decoded_instr_i[356:356], decoded_instr_i[357:357], decoded_instr_i[358:358], decoded_instr_i[359:359], decoded_instr_i[360:360], decoded_instr_i[361:361], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N3444)? { mem_q[2541:2541], mem_q[2542:2542], mem_q[2543:2543], mem_q[2544:2544], mem_q[2545:2545], mem_q[2546:2546], mem_q[2547:2547], mem_q[2548:2548], mem_q[2549:2549], mem_q[2550:2550], mem_q[2551:2551], mem_q[2552:2552], mem_q[2553:2553], mem_q[2554:2554], mem_q[2555:2555], mem_q[2556:2556], mem_q[2557:2557], mem_q[2558:2558], mem_q[2559:2559], mem_q[2560:2560], mem_q[2561:2561], mem_q[2562:2562], mem_q[2563:2563], mem_q[2564:2564], mem_q[2565:2565], mem_q[2566:2566], mem_q[2567:2567], mem_q[2568:2568], mem_q[2569:2569], mem_q[2570:2570], mem_q[2571:2571], mem_q[2572:2572], mem_q[2573:2573], mem_q[2574:2574], mem_q[2575:2575], mem_q[2576:2576], mem_q[2577:2577], mem_q[2578:2578], mem_q[2579:2579], mem_q[2580:2580], mem_q[2581:2581], mem_q[2582:2582], mem_q[2583:2583], mem_q[2584:2584], mem_q[2585:2585], mem_q[2586:2586], mem_q[2587:2587], mem_q[2588:2588], mem_q[2589:2589], mem_q[2590:2590], mem_q[2591:2591], mem_q[2592:2592], mem_q[2593:2593], mem_q[2594:2594], mem_q[2595:2595], mem_q[2596:2596], mem_q[2597:2597], mem_q[2598:2598], mem_q[2599:2599], mem_q[2600:2600], mem_q[2601:2601], mem_q[2602:2602], mem_q[2603:2603], mem_q[2604:2604], mem_q[2605:2605], mem_q[2606:2606], mem_q[2607:2607], mem_q[2608:2608], mem_q[2609:2609], mem_q[2610:2610], mem_q[2611:2611], mem_q[2612:2612], mem_q[2613:2613], mem_q[2614:2614], mem_q[2615:2615], mem_q[2616:2616], mem_q[2617:2617], mem_q[2618:2618], mem_q[2619:2619], mem_q[2620:2620], mem_q[2621:2621], mem_q[2622:2622], mem_q[2623:2623], mem_q[2624:2624], mem_q[2625:2625], mem_q[2626:2626], mem_q[2627:2627], mem_q[2628:2628], mem_q[2629:2629], mem_q[2630:2630], mem_q[2631:2631], mem_q[2632:2632], mem_q[2633:2633], mem_q[2634:2634], mem_q[2635:2635], mem_q[2636:2636], mem_q[2637:2637], mem_q[2638:2638], mem_q[2639:2639], mem_q[2640:2640], mem_q[2641:2641], mem_q[2642:2642], mem_q[2643:2643], mem_q[2644:2644], mem_q[2645:2645], mem_q[2646:2646], mem_q[2647:2647], mem_q[2648:2648], mem_q[2649:2649], mem_q[2650:2650], mem_q[2651:2651], mem_q[2652:2652], mem_q[2653:2653], mem_q[2654:2654], mem_q[2655:2655], mem_q[2656:2656], mem_q[2657:2657], mem_q[2658:2658], mem_q[2659:2659], mem_q[2660:2660], mem_q[2661:2661], mem_q[2662:2662], mem_q[2663:2663], mem_q[2664:2664], mem_q[2665:2665], mem_q[2666:2666], mem_q[2667:2667], mem_q[2668:2668], mem_q[2669:2669], mem_q[2670:2670], mem_q[2671:2671], mem_q[2672:2672], mem_q[2673:2673], mem_q[2674:2674], mem_q[2675:2675], mem_q[2676:2676], mem_q[2677:2677], mem_q[2678:2678], mem_q[2679:2679], mem_q[2680:2680], mem_q[2681:2681], mem_q[2682:2682], mem_q[2683:2683], mem_q[2684:2684], mem_q[2685:2685], mem_q[2686:2686], mem_q[2687:2687], mem_q[2688:2688], mem_q[2689:2689], mem_q[2690:2690], mem_q[2691:2691], mem_q[2692:2692], mem_q[2693:2693], mem_q[2694:2694], mem_q[2695:2695], mem_q[2696:2696], mem_q[2697:2697], mem_q[2698:2698], mem_q[2699:2699], mem_q[2700:2700], mem_q[2701:2701], mem_q[2702:2702], mem_q[2703:2703], mem_q[2704:2704], mem_q[2705:2705], mem_q[2706:2706], mem_q[2707:2707], mem_q[2708:2708], mem_q[2709:2709], mem_q[2710:2710], mem_q[2711:2711], mem_q[2712:2712], mem_q[2713:2713], mem_q[2714:2714], mem_q[2715:2715], mem_q[2716:2716], mem_q[2717:2717], mem_q[2718:2718], mem_q[2719:2719], mem_q[2720:2720], mem_q[2721:2721], mem_q[2722:2722], mem_q[2723:2723], mem_q[2724:2724], mem_q[2725:2725], mem_q[2726:2726], mem_q[2727:2727], mem_q[2728:2728], mem_q[2729:2729], mem_q[2730:2730], mem_q[2731:2731], mem_q[2732:2732], mem_q[2733:2733], mem_q[2734:2734], mem_q[2735:2735], mem_q[2736:2736], mem_q[2737:2737], mem_q[2738:2738], mem_q[2739:2739], mem_q[2740:2740], mem_q[2741:2741], mem_q[2742:2742], mem_q[2743:2743], mem_q[2744:2744], mem_q[2745:2745], mem_q[2746:2746], mem_q[2747:2747], mem_q[2748:2748], mem_q[2749:2749], mem_q[2750:2750], mem_q[2751:2751], mem_q[2752:2752], mem_q[2753:2753], mem_q[2754:2754], mem_q[2755:2755], mem_q[2756:2756], mem_q[2757:2757], mem_q[2758:2758], mem_q[2759:2759], mem_q[2760:2760], mem_q[2761:2761], mem_q[2762:2762], mem_q[2763:2763], mem_q[2764:2764], mem_q[2765:2765], mem_q[2766:2766], mem_q[2767:2767], mem_q[2768:2768], mem_q[2769:2769], mem_q[2770:2770], mem_q[2771:2771], mem_q[2772:2772], mem_q[2773:2773], mem_q[2774:2774], mem_q[2775:2775], mem_q[2776:2776], mem_q[2777:2777], mem_q[2778:2778], mem_q[2779:2779], mem_q[2780:2780], mem_q[2781:2781], mem_q[2782:2782], mem_q[2783:2783], mem_q[2784:2784], mem_q[2785:2785], mem_q[2786:2786], mem_q[2787:2787], mem_q[2788:2788], mem_q[2789:2789], mem_q[2790:2790], mem_q[2791:2791], mem_q[2792:2792], mem_q[2793:2793], mem_q[2794:2794], mem_q[2795:2795], mem_q[2796:2796], mem_q[2797:2797], mem_q[2798:2798], mem_q[2799:2799], mem_q[2800:2800], mem_q[2801:2801], mem_q[2802:2802], mem_q[2803:2803], mem_q[2804:2804], mem_q[2805:2805], mem_q[2806:2806], mem_q[2807:2807], mem_q[2808:2808], mem_q[2809:2809], mem_q[2810:2810], mem_q[2811:2811], mem_q[2812:2812], mem_q[2813:2813], mem_q[2814:2814], mem_q[2815:2815], mem_q[2816:2816], mem_q[2817:2817], mem_q[2818:2818], mem_q[2819:2819], mem_q[2820:2820], mem_q[2821:2821], mem_q[2822:2822], mem_q[2823:2823], mem_q[2824:2824], mem_q[2825:2825], mem_q[2826:2826], mem_q[2827:2827], mem_q[2828:2828], mem_q[2829:2829], mem_q[2830:2830], mem_q[2831:2831], mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835], mem_q[2836:2836], mem_q[2837:2837], mem_q[2838:2838], mem_q[2839:2839], mem_q[2840:2840], mem_q[2841:2841], mem_q[2842:2842], mem_q[2843:2843], mem_q[2844:2844], mem_q[2845:2845], mem_q[2846:2846], mem_q[2847:2847], mem_q[2848:2848], mem_q[2849:2849], mem_q[2850:2850], mem_q[2851:2851], mem_q[2852:2852], mem_q[2853:2853], mem_q[2854:2854], mem_q[2855:2855], mem_q[2856:2856], mem_q[2857:2857], mem_q[2858:2858], mem_q[2859:2859], mem_q[2860:2860], mem_q[2861:2861], mem_q[2862:2862], mem_q[2863:2863], mem_q[2864:2864], mem_q[2865:2865], mem_q[2866:2866], mem_q[2867:2867], mem_q[2868:2868], mem_q[2869:2869], mem_q[2870:2870], mem_q[2871:2871], mem_q[2872:2872], mem_q[2873:2873], mem_q[2874:2874], mem_q[2875:2875], mem_q[2876:2876], mem_q[2877:2877], mem_q[2878:2878], mem_q[2879:2879], mem_q[2880:2880], mem_q[2881:2881], mem_q[2882:2882], mem_q[2883:2883], mem_q[2884:2884], mem_q[2885:2885], mem_q[2886:2886], mem_q[2887:2887], mem_q[2888:2888], mem_q[2889:2889], mem_q[2890:2890], mem_q[2891:2891], mem_q[2892:2892], mem_q[2893:2893], mem_q[2894:2894], mem_q[2895:2895], mem_q[2896:2896], mem_q[2897:2897], mem_q[2898:2898], mem_q[2899:2899], mem_q[2900:2900], mem_q[2901:2901], mem_q[2902:2902], mem_q[2903:2903] } : 1'b0;
  assign N155 = N895;
  assign { N3813, N3812, N3811 } = (N156)? { N887, N886, N885 } : 
                                   (N884)? issue_cnt_q : 1'b0;
  assign N156 = N883;
  assign { N5885, mem_n[2902:2807], N5884, N5883, N5882, N5881, N5880, N5879, N5878, N5877, N5876, N5875, N5874, N5873, N5872, N5871, N5870, N5869, N5868, N5867, N5866, N5865, N5864, N5863, N5862, N5861, N5860, N5859, N5858, N5857, N5856, N5855, N5854, N5853, N5852, N5851, N5850, N5849, N5848, N5847, N5846, N5845, N5844, N5843, N5842, N5841, N5840, N5839, N5838, N5837, N5836, N5835, N5834, N5833, N5832, N5831, N5830, N5829, N5828, N5827, N5826, N5825, N5824, N5823, N5822, N5821, N5820, mem_n[2741:2739], N5819, N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719, N5718, N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691, mem_n[2609:2609], N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654, N5653, N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627, mem_n[2544:2541], N5626, mem_n[2539:2444], N5625, N5624, N5623, N5622, N5621, N5620, N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588, N5587, N5586, N5585, N5584, N5583, N5582, N5581, N5580, N5579, N5578, N5577, N5576, N5575, N5574, N5573, N5572, N5571, N5570, N5569, N5568, N5567, N5566, N5565, N5564, N5563, N5562, N5561, mem_n[2378:2376], N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458, N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432, mem_n[2246:2246], N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, N5418, N5417, N5416, N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, mem_n[2181:2178], N5367, mem_n[2176:2081], N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, mem_n[2015:2013], N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, mem_n[1883:1883], N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, mem_n[1818:1815], N5108, mem_n[1813:1718], N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, mem_n[1652:1650], N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, mem_n[1520:1520], N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, mem_n[1455:1452], N4849, mem_n[1450:1355], N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, mem_n[1289:1287], N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, mem_n[1157:1157], N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, mem_n[1092:1089], N4590, mem_n[1087:992], N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, mem_n[926:924], N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, mem_n[794:794], N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, mem_n[729:726], N4331, mem_n[724:629], N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, mem_n[563:561], N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, mem_n[431:431], N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073, mem_n[366:363], N4072, mem_n[361:266], N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, mem_n[200:198], N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, mem_n[68:68], N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, mem_n[3:0] } = (N156)? { N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3457, N3458, N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3467, N3468, N3469, N3470, N3471, N3472, N3473, N3474, N3475, N3476, N3477, N3478, N3479, N3480, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, N3495, N3496, N3497, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, N3515, N3516, N3517, N3518, N3519, N3520, N3521, N3522, N3523, N3524, N3525, N3526, N3527, N3528, N3529, N3530, N3531, N3532, N3533, N3534, N3535, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545, N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3553, N3554, N3555, N3556, N3557, N3558, N3559, N3560, N3561, N3562, N3563, N3564, N3565, N3566, N3567, N3568, N3569, N3570, N3571, N3572, N3573, N3574, N3575, N3576, N3577, N3578, N3579, N3580, N3581, N3582, N3583, N3584, N3585, N3586, N3587, N3588, N3589, N3590, N3591, N3592, N3593, N3594, N3595, N3596, N3597, N3598, N3599, N3600, N3601, N3602, N3603, N3604, N3605, N3606, N3607, N3608, N3609, N3610, N3611, N3612, N3613, N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3690, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3698, N3699, N3700, N3701, N3702, N3703, N3704, N3705, N3706, N3707, N3708, N3709, N3710, N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734, N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3772, N3773, N3774, N3775, N3776, N3777, N3778, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3790, N3791, N3792, N3793, N3794, N3795, N3796, N3797, N3798, N3799, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174, N3175, N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184, N3185, N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3201, N3202, N3203, N3204, N3205, N3206, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, N3339, N3340, N3341, N3342, N3343, N3344, N3345, N3346, N3347, N3348, N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3417, N3418, N3419, N3420, N3421, N3422, N3423, N3424, N3425, N3426, N3427, N3428, N3429, N3430, N3431, N3432, N3433, N3434, N3435, N3436, N3437, N3438, N3439, N3440, N3441, N3442, N3443, N2717, N2718, N2719, N2720, N2721, N2722, N2723, N2724, N2725, N2726, N2727, N2728, N2729, N2730, N2731, N2732, N2733, N2734, N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756, N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794, N2795, N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804, N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814, N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2369, N2370, N2371, N2372, N2373, N2374, N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394, N2395, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414, N2415, N2416, N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437, N2438, N2439, N2440, N2441, N2442, N2443, N2444, N2445, N2446, N2447, N2448, N2449, N2450, N2451, N2452, N2453, N2454, N2455, N2456, N2457, N2458, N2459, N2460, N2461, N2462, N2463, N2464, N2465, N2466, N2467, N2468, N2469, N2470, N2471, N2472, N2473, N2474, N2475, N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484, N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544, N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2554, N2555, N2556, N2557, N2558, N2559, N2560, N2561, N2562, N2563, N2564, N2565, N2566, N2567, N2568, N2569, N2570, N2571, N2572, N2573, N2574, N2575, N2576, N2577, N2578, N2579, N2580, N2581, N2582, N2583, N2584, N2585, N2586, N2587, N2588, N2589, N2590, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2623, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682, N2683, N2684, N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694, N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2704, N2705, N2706, N2707, N2708, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N1989, N1990, N1991, N1992, N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002, N2003, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053, N2054, N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079, N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089, N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114, N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2123, N2124, N2125, N2126, N2127, N2128, N2129, N2130, N2131, N2132, N2133, N2134, N2135, N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143, N2144, N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154, N2155, N2156, N2157, N2158, N2159, N2160, N2161, N2162, N2163, N2164, N2165, N2166, N2167, N2168, N2169, N2170, N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2179, N2180, N2181, N2182, N2183, N2184, N2185, N2186, N2187, N2188, N2189, N2190, N2191, N2192, N2193, N2194, N2195, N2196, N2197, N2198, N2199, N2200, N2201, N2202, N2203, N2204, N2205, N2206, N2207, N2208, N2209, N2210, N2211, N2212, N2213, N2214, N2215, N2216, N2217, N2218, N2219, N2220, N2221, N2222, N2223, N2224, N2225, N2226, N2227, N2228, N2229, N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260, N2261, N2262, N2263, N2264, N2265, N2266, N2267, N2268, N2269, N2270, N2271, N2272, N2273, N2274, N2275, N2276, N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2288, N2289, N2290, N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2351, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804, N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1832, N1833, N1834, N1835, N1836, N1837, N1838, N1839, N1840, N1841, N1842, N1843, N1844, N1845, N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854, N1855, N1856, N1857, N1858, N1859, N1860, N1861, N1862, N1863, N1864, N1865, N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875, N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1885, N1886, N1887, N1888, N1889, N1890, N1891, N1892, N1893, N1894, N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902, N1903, N1904, N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922, N1923, N1924, N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952, N1953, N1954, N1955, N1956, N1957, N1958, N1959, N1960, N1961, N1962, N1963, N1964, N1965, N1966, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1982, N1983, N1984, N1985, N1986, N1987, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513, N1514, N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         (N884)? mem_q : 1'b0;
  assign N5904 = (N157)? 1'b1 : 
                 (N5920)? N4007 : 1'b0;
  assign N157 = N5912;
  assign N5905 = (N158)? 1'b1 : 
                 (N5985)? N4266 : 1'b0;
  assign N158 = N5913;
  assign N5906 = (N159)? 1'b1 : 
                 (N6050)? N4525 : 1'b0;
  assign N159 = N5914;
  assign N5907 = (N160)? 1'b1 : 
                 (N6115)? N4784 : 1'b0;
  assign N160 = N5915;
  assign N5908 = (N161)? 1'b1 : 
                 (N6180)? N5043 : 1'b0;
  assign N161 = N5916;
  assign N5909 = (N162)? 1'b1 : 
                 (N6245)? N5302 : 1'b0;
  assign N162 = N5917;
  assign N5910 = (N163)? 1'b1 : 
                 (N6310)? N5561 : 1'b0;
  assign N163 = N5918;
  assign N5911 = (N164)? 1'b1 : 
                 (N6375)? N5820 : 1'b0;
  assign N164 = N5919;
  assign { N5984, N5983, N5982, N5981, N5980, N5979, N5978, N5977, N5976, N5975, N5974, N5973, N5972, N5971, N5970, N5969, N5968, N5967, N5966, N5965, N5964, N5963, N5962, N5961, N5960, N5959, N5958, N5957, N5956, N5955, N5954, N5953, N5952, N5951, N5950, N5949, N5948, N5947, N5946, N5945, N5944, N5943, N5942, N5941, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N5932, N5931, N5930, N5929, N5928, N5927, N5926, N5925, N5924, N5923, N5922, N5921 } = (N157)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5920)? { N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008 } : 1'b0;
  assign { N6049, N6048, N6047, N6046, N6045, N6044, N6043, N6042, N6041, N6040, N6039, N6038, N6037, N6036, N6035, N6034, N6033, N6032, N6031, N6030, N6029, N6028, N6027, N6026, N6025, N6024, N6023, N6022, N6021, N6020, N6019, N6018, N6017, N6016, N6015, N6014, N6013, N6012, N6011, N6010, N6009, N6008, N6007, N6006, N6005, N6004, N6003, N6002, N6001, N6000, N5999, N5998, N5997, N5996, N5995, N5994, N5993, N5992, N5991, N5990, N5989, N5988, N5987, N5986 } = (N158)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5985)? { N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267 } : 1'b0;
  assign { N6114, N6113, N6112, N6111, N6110, N6109, N6108, N6107, N6106, N6105, N6104, N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, N6093, N6092, N6091, N6090, N6089, N6088, N6087, N6086, N6085, N6084, N6083, N6082, N6081, N6080, N6079, N6078, N6077, N6076, N6075, N6074, N6073, N6072, N6071, N6070, N6069, N6068, N6067, N6066, N6065, N6064, N6063, N6062, N6061, N6060, N6059, N6058, N6057, N6056, N6055, N6054, N6053, N6052, N6051 } = (N159)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6050)? { N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526 } : 1'b0;
  assign { N6179, N6178, N6177, N6176, N6175, N6174, N6173, N6172, N6171, N6170, N6169, N6168, N6167, N6166, N6165, N6164, N6163, N6162, N6161, N6160, N6159, N6158, N6157, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N6149, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N6141, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N6133, N6132, N6131, N6130, N6129, N6128, N6127, N6126, N6125, N6124, N6123, N6122, N6121, N6120, N6119, N6118, N6117, N6116 } = (N160)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6115)? { N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785 } : 1'b0;
  assign { N6244, N6243, N6242, N6241, N6240, N6239, N6238, N6237, N6236, N6235, N6234, N6233, N6232, N6231, N6230, N6229, N6228, N6227, N6226, N6225, N6224, N6223, N6222, N6221, N6220, N6219, N6218, N6217, N6216, N6215, N6214, N6213, N6212, N6211, N6210, N6209, N6208, N6207, N6206, N6205, N6204, N6203, N6202, N6201, N6200, N6199, N6198, N6197, N6196, N6195, N6194, N6193, N6192, N6191, N6190, N6189, N6188, N6187, N6186, N6185, N6184, N6183, N6182, N6181 } = (N161)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6180)? { N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044 } : 1'b0;
  assign { N6309, N6308, N6307, N6306, N6305, N6304, N6303, N6302, N6301, N6300, N6299, N6298, N6297, N6296, N6295, N6294, N6293, N6292, N6291, N6290, N6289, N6288, N6287, N6286, N6285, N6284, N6283, N6282, N6281, N6280, N6279, N6278, N6277, N6276, N6275, N6274, N6273, N6272, N6271, N6270, N6269, N6268, N6267, N6266, N6265, N6264, N6263, N6262, N6261, N6260, N6259, N6258, N6257, N6256, N6255, N6254, N6253, N6252, N6251, N6250, N6249, N6248, N6247, N6246 } = (N162)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6245)? { N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303 } : 1'b0;
  assign { N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366, N6365, N6364, N6363, N6362, N6361, N6360, N6359, N6358, N6357, N6356, N6355, N6354, N6353, N6352, N6351, N6350, N6349, N6348, N6347, N6346, N6345, N6344, N6343, N6342, N6341, N6340, N6339, N6338, N6337, N6336, N6335, N6334, N6333, N6332, N6331, N6330, N6329, N6328, N6327, N6326, N6325, N6324, N6323, N6322, N6321, N6320, N6319, N6318, N6317, N6316, N6315, N6314, N6313, N6312, N6311 } = (N163)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6310)? { N5625, N5624, N5623, N5622, N5621, N5620, N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588, N5587, N5586, N5585, N5584, N5583, N5582, N5581, N5580, N5579, N5578, N5577, N5576, N5575, N5574, N5573, N5572, N5571, N5570, N5569, N5568, N5567, N5566, N5565, N5564, N5563, N5562 } : 1'b0;
  assign { N6439, N6438, N6437, N6436, N6435, N6434, N6433, N6432, N6431, N6430, N6429, N6428, N6427, N6426, N6425, N6424, N6423, N6422, N6421, N6420, N6419, N6418, N6417, N6416, N6415, N6414, N6413, N6412, N6411, N6410, N6409, N6408, N6407, N6406, N6405, N6404, N6403, N6402, N6401, N6400, N6399, N6398, N6397, N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377, N6376 } = (N164)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6375)? { N5884, N5883, N5882, N5881, N5880, N5879, N5878, N5877, N5876, N5875, N5874, N5873, N5872, N5871, N5870, N5869, N5868, N5867, N5866, N5865, N5864, N5863, N5862, N5861, N5860, N5859, N5858, N5857, N5856, N5855, N5854, N5853, N5852, N5851, N5850, N5849, N5848, N5847, N5846, N5845, N5844, N5843, N5842, N5841, N5840, N5839, N5838, N5837, N5836, N5835, N5834, N5833, N5832, N5831, N5830, N5829, N5828, N5827, N5826, N5825, N5824, N5823, N5822, N5821 } : 1'b0;
  assign { N6503, N6502, N6501, N6500, N6499, N6498, N6497, N6496, N6495, N6494, N6493, N6492, N6491, N6490, N6489, N6488, N6487, N6486, N6485, N6484, N6483, N6482, N6481, N6480, N6479, N6478, N6477, N6476, N6475, N6474, N6473, N6472, N6471, N6470, N6469, N6468, N6467, N6466, N6465, N6464, N6463, N6462, N6461, N6460, N6459, N6458, N6457, N6456, N6455, N6454, N6453, N6452, N6451, N6450, N6449, N6448, N6447, N6446, N6445, N6444, N6443, N6442, N6441, N6440 } = (N157)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5920)? { N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814 } : 1'b0;
  assign { N6567, N6566, N6565, N6564, N6563, N6562, N6561, N6560, N6559, N6558, N6557, N6556, N6555, N6554, N6553, N6552, N6551, N6550, N6549, N6548, N6547, N6546, N6545, N6544, N6543, N6542, N6541, N6540, N6539, N6538, N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530, N6529, N6528, N6527, N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, N6518, N6517, N6516, N6515, N6514, N6513, N6512, N6511, N6510, N6509, N6508, N6507, N6506, N6505, N6504 } = (N158)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5985)? { N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073 } : 1'b0;
  assign { N6631, N6630, N6629, N6628, N6627, N6626, N6625, N6624, N6623, N6622, N6621, N6620, N6619, N6618, N6617, N6616, N6615, N6614, N6613, N6612, N6611, N6610, N6609, N6608, N6607, N6606, N6605, N6604, N6603, N6602, N6601, N6600, N6599, N6598, N6597, N6596, N6595, N6594, N6593, N6592, N6591, N6590, N6589, N6588, N6587, N6586, N6585, N6584, N6583, N6582, N6581, N6580, N6579, N6578, N6577, N6576, N6575, N6574, N6573, N6572, N6571, N6570, N6569, N6568 } = (N159)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6050)? { N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332 } : 1'b0;
  assign { N6695, N6694, N6693, N6692, N6691, N6690, N6689, N6688, N6687, N6686, N6685, N6684, N6683, N6682, N6681, N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667, N6666, N6665, N6664, N6663, N6662, N6661, N6660, N6659, N6658, N6657, N6656, N6655, N6654, N6653, N6652, N6651, N6650, N6649, N6648, N6647, N6646, N6645, N6644, N6643, N6642, N6641, N6640, N6639, N6638, N6637, N6636, N6635, N6634, N6633, N6632 } = (N160)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6115)? { N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591 } : 1'b0;
  assign { N6759, N6758, N6757, N6756, N6755, N6754, N6753, N6752, N6751, N6750, N6749, N6748, N6747, N6746, N6745, N6744, N6743, N6742, N6741, N6740, N6739, N6738, N6737, N6736, N6735, N6734, N6733, N6732, N6731, N6730, N6729, N6728, N6727, N6726, N6725, N6724, N6723, N6722, N6721, N6720, N6719, N6718, N6717, N6716, N6715, N6714, N6713, N6712, N6711, N6710, N6709, N6708, N6707, N6706, N6705, N6704, N6703, N6702, N6701, N6700, N6699, N6698, N6697, N6696 } = (N161)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6180)? { N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850 } : 1'b0;
  assign { N6823, N6822, N6821, N6820, N6819, N6818, N6817, N6816, N6815, N6814, N6813, N6812, N6811, N6810, N6809, N6808, N6807, N6806, N6805, N6804, N6803, N6802, N6801, N6800, N6799, N6798, N6797, N6796, N6795, N6794, N6793, N6792, N6791, N6790, N6789, N6788, N6787, N6786, N6785, N6784, N6783, N6782, N6781, N6780, N6779, N6778, N6777, N6776, N6775, N6774, N6773, N6772, N6771, N6770, N6769, N6768, N6767, N6766, N6765, N6764, N6763, N6762, N6761, N6760 } = (N162)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6245)? { N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109 } : 1'b0;
  assign { N6887, N6886, N6885, N6884, N6883, N6882, N6881, N6880, N6879, N6878, N6877, N6876, N6875, N6874, N6873, N6872, N6871, N6870, N6869, N6868, N6867, N6866, N6865, N6864, N6863, N6862, N6861, N6860, N6859, N6858, N6857, N6856, N6855, N6854, N6853, N6852, N6851, N6850, N6849, N6848, N6847, N6846, N6845, N6844, N6843, N6842, N6841, N6840, N6839, N6838, N6837, N6836, N6835, N6834, N6833, N6832, N6831, N6830, N6829, N6828, N6827, N6826, N6825, N6824 } = (N163)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6310)? { N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, N5418, N5417, N5416, N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368 } : 1'b0;
  assign { N6951, N6950, N6949, N6948, N6947, N6946, N6945, N6944, N6943, N6942, N6941, N6940, N6939, N6938, N6937, N6936, N6935, N6934, N6933, N6932, N6931, N6930, N6929, N6928, N6927, N6926, N6925, N6924, N6923, N6922, N6921, N6920, N6919, N6918, N6917, N6916, N6915, N6914, N6913, N6912, N6911, N6910, N6909, N6908, N6907, N6906, N6905, N6904, N6903, N6902, N6901, N6900, N6899, N6898, N6897, N6896, N6895, N6894, N6893, N6892, N6891, N6890, N6889, N6888 } = (N164)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6375)? { N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654, N5653, N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627 } : 1'b0;
  assign { N7085, N7084, N7083, N7082, N7081, N7080, N7079, N7078, N7077, N7076, N7075, N7074, N7073, N7072, N7071, N7070, N7069, N7068, N7067, N7066, N7065, N7064, N7063, N7062, N7061, N7060, N7059, N7058, N7057, N7056, N7055, N7054, N7053, N7052, N7051, N7050, N7049, N7048, N7047, N7046, N7045, N7044, N7043, N7042, N7041, N7040, N7039, N7038, N7037, N7036, N7035, N7034, N7033, N7032, N7031, N7030, N7029, N7028, N7027, N7026, N7025, N7024, N7023, N7022, N7021, N7020, N7019, N7018, N7017, N7016, N7015, N7014, N7013, N7012, N7011, N7010, N7009, N7008, N7007, N7006, N7005, N7004, N7003, N7002, N7001, N7000, N6999, N6998, N6997, N6996, N6995, N6994, N6993, N6992, N6991, N6990, N6989, N6988, N6987, N6986, N6985, N6984, N6983, N6982, N6981, N6980, N6979, N6978, N6977, N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, N6957 } = (N157)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N5920)? { N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878 } : 1'b0;
  assign { N7214, N7213, N7212, N7211, N7210, N7209, N7208, N7207, N7206, N7205, N7204, N7203, N7202, N7201, N7200, N7199, N7198, N7197, N7196, N7195, N7194, N7193, N7192, N7191, N7190, N7189, N7188, N7187, N7186, N7185, N7184, N7183, N7182, N7181, N7180, N7179, N7178, N7177, N7176, N7175, N7174, N7173, N7172, N7171, N7170, N7169, N7168, N7167, N7166, N7165, N7164, N7163, N7162, N7161, N7160, N7159, N7158, N7157, N7156, N7155, N7154, N7153, N7152, N7151, N7150, N7149, N7148, N7147, N7146, N7145, N7144, N7143, N7142, N7141, N7140, N7139, N7138, N7137, N7136, N7135, N7134, N7133, N7132, N7131, N7130, N7129, N7128, N7127, N7126, N7125, N7124, N7123, N7122, N7121, N7120, N7119, N7118, N7117, N7116, N7115, N7114, N7113, N7112, N7111, N7110, N7109, N7108, N7107, N7106, N7105, N7104, N7103, N7102, N7101, N7100, N7099, N7098, N7097, N7096, N7095, N7094, N7093, N7092, N7091, N7090, N7089, N7088, N7087, N7086 } = (N158)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N5985)? { N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137 } : 1'b0;
  assign { N7343, N7342, N7341, N7340, N7339, N7338, N7337, N7336, N7335, N7334, N7333, N7332, N7331, N7330, N7329, N7328, N7327, N7326, N7325, N7324, N7323, N7322, N7321, N7320, N7319, N7318, N7317, N7316, N7315, N7314, N7313, N7312, N7311, N7310, N7309, N7308, N7307, N7306, N7305, N7304, N7303, N7302, N7301, N7300, N7299, N7298, N7297, N7296, N7295, N7294, N7293, N7292, N7291, N7290, N7289, N7288, N7287, N7286, N7285, N7284, N7283, N7282, N7281, N7280, N7279, N7278, N7277, N7276, N7275, N7274, N7273, N7272, N7271, N7270, N7269, N7268, N7267, N7266, N7265, N7264, N7263, N7262, N7261, N7260, N7259, N7258, N7257, N7256, N7255, N7254, N7253, N7252, N7251, N7250, N7249, N7248, N7247, N7246, N7245, N7244, N7243, N7242, N7241, N7240, N7239, N7238, N7237, N7236, N7235, N7234, N7233, N7232, N7231, N7230, N7229, N7228, N7227, N7226, N7225, N7224, N7223, N7222, N7221, N7220, N7219, N7218, N7217, N7216, N7215 } = (N159)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N6050)? { N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396 } : 1'b0;
  assign { N7472, N7471, N7470, N7469, N7468, N7467, N7466, N7465, N7464, N7463, N7462, N7461, N7460, N7459, N7458, N7457, N7456, N7455, N7454, N7453, N7452, N7451, N7450, N7449, N7448, N7447, N7446, N7445, N7444, N7443, N7442, N7441, N7440, N7439, N7438, N7437, N7436, N7435, N7434, N7433, N7432, N7431, N7430, N7429, N7428, N7427, N7426, N7425, N7424, N7423, N7422, N7421, N7420, N7419, N7418, N7417, N7416, N7415, N7414, N7413, N7412, N7411, N7410, N7409, N7408, N7407, N7406, N7405, N7404, N7403, N7402, N7401, N7400, N7399, N7398, N7397, N7396, N7395, N7394, N7393, N7392, N7391, N7390, N7389, N7388, N7387, N7386, N7385, N7384, N7383, N7382, N7381, N7380, N7379, N7378, N7377, N7376, N7375, N7374, N7373, N7372, N7371, N7370, N7369, N7368, N7367, N7366, N7365, N7364, N7363, N7362, N7361, N7360, N7359, N7358, N7357, N7356, N7355, N7354, N7353, N7352, N7351, N7350, N7349, N7348, N7347, N7346, N7345, N7344 } = (N160)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N6115)? { N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655 } : 1'b0;
  assign { N7601, N7600, N7599, N7598, N7597, N7596, N7595, N7594, N7593, N7592, N7591, N7590, N7589, N7588, N7587, N7586, N7585, N7584, N7583, N7582, N7581, N7580, N7579, N7578, N7577, N7576, N7575, N7574, N7573, N7572, N7571, N7570, N7569, N7568, N7567, N7566, N7565, N7564, N7563, N7562, N7561, N7560, N7559, N7558, N7557, N7556, N7555, N7554, N7553, N7552, N7551, N7550, N7549, N7548, N7547, N7546, N7545, N7544, N7543, N7542, N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534, N7533, N7532, N7531, N7530, N7529, N7528, N7527, N7526, N7525, N7524, N7523, N7522, N7521, N7520, N7519, N7518, N7517, N7516, N7515, N7514, N7513, N7512, N7511, N7510, N7509, N7508, N7507, N7506, N7505, N7504, N7503, N7502, N7501, N7500, N7499, N7498, N7497, N7496, N7495, N7494, N7493, N7492, N7491, N7490, N7489, N7488, N7487, N7486, N7485, N7484, N7483, N7482, N7481, N7480, N7479, N7478, N7477, N7476, N7475, N7474, N7473 } = (N161)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N6180)? { N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914 } : 1'b0;
  assign { N7730, N7729, N7728, N7727, N7726, N7725, N7724, N7723, N7722, N7721, N7720, N7719, N7718, N7717, N7716, N7715, N7714, N7713, N7712, N7711, N7710, N7709, N7708, N7707, N7706, N7705, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696, N7695, N7694, N7693, N7692, N7691, N7690, N7689, N7688, N7687, N7686, N7685, N7684, N7683, N7682, N7681, N7680, N7679, N7678, N7677, N7676, N7675, N7674, N7673, N7672, N7671, N7670, N7669, N7668, N7667, N7666, N7665, N7664, N7663, N7662, N7661, N7660, N7659, N7658, N7657, N7656, N7655, N7654, N7653, N7652, N7651, N7650, N7649, N7648, N7647, N7646, N7645, N7644, N7643, N7642, N7641, N7640, N7639, N7638, N7637, N7636, N7635, N7634, N7633, N7632, N7631, N7630, N7629, N7628, N7627, N7626, N7625, N7624, N7623, N7622, N7621, N7620, N7619, N7618, N7617, N7616, N7615, N7614, N7613, N7612, N7611, N7610, N7609, N7608, N7607, N7606, N7605, N7604, N7603, N7602 } = (N162)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N6245)? { N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173 } : 1'b0;
  assign { N7859, N7858, N7857, N7856, N7855, N7854, N7853, N7852, N7851, N7850, N7849, N7848, N7847, N7846, N7845, N7844, N7843, N7842, N7841, N7840, N7839, N7838, N7837, N7836, N7835, N7834, N7833, N7832, N7831, N7830, N7829, N7828, N7827, N7826, N7825, N7824, N7823, N7822, N7821, N7820, N7819, N7818, N7817, N7816, N7815, N7814, N7813, N7812, N7811, N7810, N7809, N7808, N7807, N7806, N7805, N7804, N7803, N7802, N7801, N7800, N7799, N7798, N7797, N7796, N7795, N7794, N7793, N7792, N7791, N7790, N7789, N7788, N7787, N7786, N7785, N7784, N7783, N7782, N7781, N7780, N7779, N7778, N7777, N7776, N7775, N7774, N7773, N7772, N7771, N7770, N7769, N7768, N7767, N7766, N7765, N7764, N7763, N7762, N7761, N7760, N7759, N7758, N7757, N7756, N7755, N7754, N7753, N7752, N7751, N7750, N7749, N7748, N7747, N7746, N7745, N7744, N7743, N7742, N7741, N7740, N7739, N7738, N7737, N7736, N7735, N7734, N7733, N7732, N7731 } = (N163)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N6310)? { N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458, N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432 } : 1'b0;
  assign { N7988, N7987, N7986, N7985, N7984, N7983, N7982, N7981, N7980, N7979, N7978, N7977, N7976, N7975, N7974, N7973, N7972, N7971, N7970, N7969, N7968, N7967, N7966, N7965, N7964, N7963, N7962, N7961, N7960, N7959, N7958, N7957, N7956, N7955, N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946, N7945, N7944, N7943, N7942, N7941, N7940, N7939, N7938, N7937, N7936, N7935, N7934, N7933, N7932, N7931, N7930, N7929, N7928, N7927, N7926, N7925, N7924, N7923, N7922, N7921, N7920, N7919, N7918, N7917, N7916, N7915, N7914, N7913, N7912, N7911, N7910, N7909, N7908, N7907, N7906, N7905, N7904, N7903, N7902, N7901, N7900, N7899, N7898, N7897, N7896, N7895, N7894, N7893, N7892, N7891, N7890, N7889, N7888, N7887, N7886, N7885, N7884, N7883, N7882, N7881, N7880, N7879, N7878, N7877, N7876, N7875, N7874, N7873, N7872, N7871, N7870, N7869, N7868, N7867, N7866, N7865, N7864, N7863, N7862, N7861, N7860 } = (N164)? ex_i[128:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N6375)? { N5819, N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719, N5718, N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691 } : 1'b0;
  assign { N8064, N8063, N8062, N8061, N8060, N8059, N8058, N8057, N8056, N8055, N8054, N8053, N8052, N8051, N8050, N8049, N8048, N8047, N8046, N8045, N8044, N8043, N8042, N8041, N8040, N8039, N8038, N8037, N8036, N8035, N8034, N8033, N8032, N8031, N8030, N8029, N8028, N8027, N8026, N8025, N8024, N8023, N8022, N8021, N8020, N8019, N8018, N8017, N8016, N8015, N8014, N8013, N8012, N8011, N8010, N8009, N8008, N8007, N8006, N8005, N8004, N8003, N8002, N8001 } = (N157)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5920)? { N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943 } : 1'b0;
  assign { N8128, N8127, N8126, N8125, N8124, N8123, N8122, N8121, N8120, N8119, N8118, N8117, N8116, N8115, N8114, N8113, N8112, N8111, N8110, N8109, N8108, N8107, N8106, N8105, N8104, N8103, N8102, N8101, N8100, N8099, N8098, N8097, N8096, N8095, N8094, N8093, N8092, N8091, N8090, N8089, N8088, N8087, N8086, N8085, N8084, N8083, N8082, N8081, N8080, N8079, N8078, N8077, N8076, N8075, N8074, N8073, N8072, N8071, N8070, N8069, N8068, N8067, N8066, N8065 } = (N158)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5985)? { N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202 } : 1'b0;
  assign { N8192, N8191, N8190, N8189, N8188, N8187, N8186, N8185, N8184, N8183, N8182, N8181, N8180, N8179, N8178, N8177, N8176, N8175, N8174, N8173, N8172, N8171, N8170, N8169, N8168, N8167, N8166, N8165, N8164, N8163, N8162, N8161, N8160, N8159, N8158, N8157, N8156, N8155, N8154, N8153, N8152, N8151, N8150, N8149, N8148, N8147, N8146, N8145, N8144, N8143, N8142, N8141, N8140, N8139, N8138, N8137, N8136, N8135, N8134, N8133, N8132, N8131, N8130, N8129 } = (N159)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6050)? { N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461 } : 1'b0;
  assign { N8256, N8255, N8254, N8253, N8252, N8251, N8250, N8249, N8248, N8247, N8246, N8245, N8244, N8243, N8242, N8241, N8240, N8239, N8238, N8237, N8236, N8235, N8234, N8233, N8232, N8231, N8230, N8229, N8228, N8227, N8226, N8225, N8224, N8223, N8222, N8221, N8220, N8219, N8218, N8217, N8216, N8215, N8214, N8213, N8212, N8211, N8210, N8209, N8208, N8207, N8206, N8205, N8204, N8203, N8202, N8201, N8200, N8199, N8198, N8197, N8196, N8195, N8194, N8193 } = (N160)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6115)? { N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720 } : 1'b0;
  assign { N8320, N8319, N8318, N8317, N8316, N8315, N8314, N8313, N8312, N8311, N8310, N8309, N8308, N8307, N8306, N8305, N8304, N8303, N8302, N8301, N8300, N8299, N8298, N8297, N8296, N8295, N8294, N8293, N8292, N8291, N8290, N8289, N8288, N8287, N8286, N8285, N8284, N8283, N8282, N8281, N8280, N8279, N8278, N8277, N8276, N8275, N8274, N8273, N8272, N8271, N8270, N8269, N8268, N8267, N8266, N8265, N8264, N8263, N8262, N8261, N8260, N8259, N8258, N8257 } = (N161)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6180)? { N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979 } : 1'b0;
  assign { N8384, N8383, N8382, N8381, N8380, N8379, N8378, N8377, N8376, N8375, N8374, N8373, N8372, N8371, N8370, N8369, N8368, N8367, N8366, N8365, N8364, N8363, N8362, N8361, N8360, N8359, N8358, N8357, N8356, N8355, N8354, N8353, N8352, N8351, N8350, N8349, N8348, N8347, N8346, N8345, N8344, N8343, N8342, N8341, N8340, N8339, N8338, N8337, N8336, N8335, N8334, N8333, N8332, N8331, N8330, N8329, N8328, N8327, N8326, N8325, N8324, N8323, N8322, N8321 } = (N162)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6245)? { N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238 } : 1'b0;
  assign { N8448, N8447, N8446, N8445, N8444, N8443, N8442, N8441, N8440, N8439, N8438, N8437, N8436, N8435, N8434, N8433, N8432, N8431, N8430, N8429, N8428, N8427, N8426, N8425, N8424, N8423, N8422, N8421, N8420, N8419, N8418, N8417, N8416, N8415, N8414, N8413, N8412, N8411, N8410, N8409, N8408, N8407, N8406, N8405, N8404, N8403, N8402, N8401, N8400, N8399, N8398, N8397, N8396, N8395, N8394, N8393, N8392, N8391, N8390, N8389, N8388, N8387, N8386, N8385 } = (N163)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6310)? { N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497 } : 1'b0;
  assign { N8512, N8511, N8510, N8509, N8508, N8507, N8506, N8505, N8504, N8503, N8502, N8501, N8500, N8499, N8498, N8497, N8496, N8495, N8494, N8493, N8492, N8491, N8490, N8489, N8488, N8487, N8486, N8485, N8484, N8483, N8482, N8481, N8480, N8479, N8478, N8477, N8476, N8475, N8474, N8473, N8472, N8471, N8470, N8469, N8468, N8467, N8466, N8465, N8464, N8463, N8462, N8461, N8460, N8459, N8458, N8457, N8456, N8455, N8454, N8453, N8452, N8451, N8450, N8449 } = (N164)? ex_i[128:65] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6375)? { N5819, N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756 } : 1'b0;
  assign { N9024, N9023, N9022, N9021, N9020, N9019, N9018, N9017, N9016, N9015, N9014, N9013, N9012, N9011, N9010, N9009, N9008, N9007, N9006, N9005, N9004, N9003, N9002, N9001, N9000, N8999, N8998, N8997, N8996, N8995, N8994, N8993, N8992, N8991, N8990, N8989, N8988, N8987, N8986, N8985, N8984, N8983, N8982, N8981, N8980, N8979, N8978, N8977, N8976, N8975, N8974, N8973, N8972, N8971, N8970, N8969, N8968, N8967, N8966, N8965, N8964, N8963, N8962, N8961, N8960, N8959, N8958, N8957, N8956, N8955, N8954, N8953, N8952, N8951, N8950, N8949, N8948, N8947, N8946, N8945, N8944, N8943, N8942, N8941, N8940, N8939, N8938, N8937, N8936, N8935, N8934, N8933, N8932, N8931, N8930, N8929, N8928, N8927, N8926, N8925, N8924, N8923, N8922, N8921, N8920, N8919, N8918, N8917, N8916, N8915, N8914, N8913, N8912, N8911, N8910, N8909, N8908, N8907, N8906, N8905, N8904, N8903, N8902, N8901, N8900, N8899, N8898, N8897, N8896, N8895, N8894, N8893, N8892, N8891, N8890, N8889, N8888, N8887, N8886, N8885, N8884, N8883, N8882, N8881, N8880, N8879, N8878, N8877, N8876, N8875, N8874, N8873, N8872, N8871, N8870, N8869, N8868, N8867, N8866, N8865, N8864, N8863, N8862, N8861, N8860, N8859, N8858, N8857, N8856, N8855, N8854, N8853, N8852, N8851, N8850, N8849, N8848, N8847, N8846, N8845, N8844, N8843, N8842, N8841, N8840, N8839, N8838, N8837, N8836, N8835, N8834, N8833, N8832, N8831, N8830, N8829, N8828, N8827, N8826, N8825, N8824, N8823, N8822, N8821, N8820, N8819, N8818, N8817, N8816, N8815, N8814, N8813, N8812, N8811, N8810, N8809, N8808, N8807, N8806, N8805, N8804, N8803, N8802, N8801, N8800, N8799, N8798, N8797, N8796, N8795, N8794, N8793, N8792, N8791, N8790, N8789, N8788, N8787, N8786, N8785, N8784, N8783, N8782, N8781, N8780, N8779, N8778, N8777, N8776, N8775, N8774, N8773, N8772, N8771, N8770, N8769, N8768, N8767, N8766, N8765, N8764, N8763, N8762, N8761, N8760, N8759, N8758, N8757, N8756, N8755, N8754, N8753, N8752, N8751, N8750, N8749, N8748, N8747, N8746, N8745, N8744, N8743, N8742, N8741, N8740, N8739, N8738, N8737, N8736, N8735, N8734, N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N8704, N8703, N8702, N8701, N8700, N8699, N8698, N8697, N8696, N8695, N8694, N8693, N8692, N8691, N8690, N8689, N8688, N8687, N8686, N8685, N8684, N8683, N8682, N8681, N8680, N8679, N8678, N8677, N8676, N8675, N8674, N8673, N8672, N8671, N8670, N8669, N8668, N8667, N8666, N8665, N8664, N8663, N8662, N8661, N8660, N8659, N8658, N8657, N8656, N8655, N8654, N8653, N8652, N8651, N8650, N8649, N8648, N8647, N8646, N8645, N8644, N8643, N8642, N8641, N8640, N8639, N8638, N8637, N8636, N8635, N8634, N8633, N8632, N8631, N8630, N8629, N8628, N8627, N8626, N8625, N8624, N8623, N8622, N8621, N8620, N8619, N8618, N8617, N8616, N8615, N8614, N8613, N8612, N8611, N8610, N8609, N8608, N8607, N8606, N8605, N8604, N8603, N8602, N8601, N8600, N8599, N8598, N8597, N8596, N8595, N8594, N8593, N8592, N8591, N8590, N8589, N8588, N8587, N8586, N8585, N8584, N8583, N8582, N8581, N8580, N8579, N8578, N8577, N8576, N8575, N8574, N8573, N8572, N8571, N8570, N8569, N8568, N8567, N8566, N8565, N8564, N8563, N8562, N8561, N8560, N8559, N8558, N8557, N8556, N8555, N8554, N8553, N8552, N8551, N8550, N8549, N8548, N8547, N8546, N8545, N8544, N8543, N8542, N8541, N8540, N8539, N8538, N8537, N8536, N8535, N8534, N8533, N8532, N8531, N8530, N8529, N8528, N8527, N8526, N8525, N8524, N8523, N8522, N8521, N8520, N8519, N8518, N8517, N8516, N8515, N8514, N8513 } = (N165)? { N8512, N8511, N8510, N8509, N8508, N8507, N8506, N8505, N8504, N8503, N8502, N8501, N8500, N8499, N8498, N8497, N8496, N8495, N8494, N8493, N8492, N8491, N8490, N8489, N8488, N8487, N8486, N8485, N8484, N8483, N8482, N8481, N8480, N8479, N8478, N8477, N8476, N8475, N8474, N8473, N8472, N8471, N8470, N8469, N8468, N8467, N8466, N8465, N8464, N8463, N8462, N8461, N8460, N8459, N8458, N8457, N8456, N8455, N8454, N8453, N8452, N8451, N8450, N8449, N8448, N8447, N8446, N8445, N8444, N8443, N8442, N8441, N8440, N8439, N8438, N8437, N8436, N8435, N8434, N8433, N8432, N8431, N8430, N8429, N8428, N8427, N8426, N8425, N8424, N8423, N8422, N8421, N8420, N8419, N8418, N8417, N8416, N8415, N8414, N8413, N8412, N8411, N8410, N8409, N8408, N8407, N8406, N8405, N8404, N8403, N8402, N8401, N8400, N8399, N8398, N8397, N8396, N8395, N8394, N8393, N8392, N8391, N8390, N8389, N8388, N8387, N8386, N8385, N8384, N8383, N8382, N8381, N8380, N8379, N8378, N8377, N8376, N8375, N8374, N8373, N8372, N8371, N8370, N8369, N8368, N8367, N8366, N8365, N8364, N8363, N8362, N8361, N8360, N8359, N8358, N8357, N8356, N8355, N8354, N8353, N8352, N8351, N8350, N8349, N8348, N8347, N8346, N8345, N8344, N8343, N8342, N8341, N8340, N8339, N8338, N8337, N8336, N8335, N8334, N8333, N8332, N8331, N8330, N8329, N8328, N8327, N8326, N8325, N8324, N8323, N8322, N8321, N8320, N8319, N8318, N8317, N8316, N8315, N8314, N8313, N8312, N8311, N8310, N8309, N8308, N8307, N8306, N8305, N8304, N8303, N8302, N8301, N8300, N8299, N8298, N8297, N8296, N8295, N8294, N8293, N8292, N8291, N8290, N8289, N8288, N8287, N8286, N8285, N8284, N8283, N8282, N8281, N8280, N8279, N8278, N8277, N8276, N8275, N8274, N8273, N8272, N8271, N8270, N8269, N8268, N8267, N8266, N8265, N8264, N8263, N8262, N8261, N8260, N8259, N8258, N8257, N8256, N8255, N8254, N8253, N8252, N8251, N8250, N8249, N8248, N8247, N8246, N8245, N8244, N8243, N8242, N8241, N8240, N8239, N8238, N8237, N8236, N8235, N8234, N8233, N8232, N8231, N8230, N8229, N8228, N8227, N8226, N8225, N8224, N8223, N8222, N8221, N8220, N8219, N8218, N8217, N8216, N8215, N8214, N8213, N8212, N8211, N8210, N8209, N8208, N8207, N8206, N8205, N8204, N8203, N8202, N8201, N8200, N8199, N8198, N8197, N8196, N8195, N8194, N8193, N8192, N8191, N8190, N8189, N8188, N8187, N8186, N8185, N8184, N8183, N8182, N8181, N8180, N8179, N8178, N8177, N8176, N8175, N8174, N8173, N8172, N8171, N8170, N8169, N8168, N8167, N8166, N8165, N8164, N8163, N8162, N8161, N8160, N8159, N8158, N8157, N8156, N8155, N8154, N8153, N8152, N8151, N8150, N8149, N8148, N8147, N8146, N8145, N8144, N8143, N8142, N8141, N8140, N8139, N8138, N8137, N8136, N8135, N8134, N8133, N8132, N8131, N8130, N8129, N8128, N8127, N8126, N8125, N8124, N8123, N8122, N8121, N8120, N8119, N8118, N8117, N8116, N8115, N8114, N8113, N8112, N8111, N8110, N8109, N8108, N8107, N8106, N8105, N8104, N8103, N8102, N8101, N8100, N8099, N8098, N8097, N8096, N8095, N8094, N8093, N8092, N8091, N8090, N8089, N8088, N8087, N8086, N8085, N8084, N8083, N8082, N8081, N8080, N8079, N8078, N8077, N8076, N8075, N8074, N8073, N8072, N8071, N8070, N8069, N8068, N8067, N8066, N8065, N8064, N8063, N8062, N8061, N8060, N8059, N8058, N8057, N8056, N8055, N8054, N8053, N8052, N8051, N8050, N8049, N8048, N8047, N8046, N8045, N8044, N8043, N8042, N8041, N8040, N8039, N8038, N8037, N8036, N8035, N8034, N8033, N8032, N8031, N8030, N8029, N8028, N8027, N8026, N8025, N8024, N8023, N8022, N8021, N8020, N8019, N8018, N8017, N8016, N8015, N8014, N8013, N8012, N8011, N8010, N8009, N8008, N8007, N8006, N8005, N8004, N8003, N8002, N8001 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N166)? { N5819, N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943 } : 1'b0;
  assign N165 = N7999;
  assign N166 = N8000;
  assign { N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002, N10001, N10000, N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9967, N9966, N9965, N9964, N9963, N9962, N9961, N9960, N9959, N9958, N9957, N9956, N9955, N9954, N9953, N9952, N9951, N9950, N9949, N9948, N9947, N9946, N9945, N9944, N9943, N9942, N9941, N9940, N9939, N9938, N9937, N9936, N9935, N9934, N9933, N9932, N9931, N9930, N9929, N9928, N9927, N9926, N9925, N9924, N9923, N9922, N9921, N9920, N9919, N9918, N9917, N9916, N9915, N9914, N9913, N9912, N9911, N9910, N9909, N9908, N9907, N9906, N9905, N9904, N9903, N9902, N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838, N9837, N9836, N9835, N9834, N9833, N9832, N9831, N9830, N9829, N9828, N9827, N9826, N9825, N9824, N9823, N9822, N9821, N9820, N9819, N9818, N9817, N9816, N9815, N9814, N9813, N9812, N9811, N9810, N9809, N9808, N9807, N9806, N9805, N9804, N9803, N9802, N9801, N9800, N9799, N9798, N9797, N9796, N9795, N9794, N9793, N9792, N9791, N9790, N9789, N9788, N9787, N9786, N9785, N9784, N9783, N9782, N9781, N9780, N9779, N9778, N9777, N9776, N9775, N9774, N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742, N9741, N9740, N9739, N9738, N9737, N9736, N9735, N9734, N9733, N9732, N9731, N9730, N9729, N9728, N9727, N9726, N9725, N9724, N9723, N9722, N9721, N9720, N9719, N9718, N9717, N9716, N9715, N9714, N9713, N9712, N9711, N9710, N9709, N9708, N9707, N9706, N9705, N9704, N9703, N9702, N9701, N9700, N9699, N9698, N9697, N9696, N9695, N9694, N9693, N9692, N9691, N9690, N9689, N9688, N9687, N9686, N9685, N9684, N9683, N9682, N9681, N9680, N9679, N9678, N9677, N9676, N9675, N9674, N9673, N9672, N9671, N9670, N9669, N9668, N9667, N9666, N9665, N9664, N9663, N9662, N9661, N9660, N9659, N9658, N9657, N9656, N9655, N9654, N9653, N9652, N9651, N9650, N9649, N9648, N9647, N9646, N9645, N9644, N9643, N9642, N9641, N9640, N9639, N9638, N9637, N9636, N9635, N9634, N9633, N9632, N9631, N9630, N9629, N9628, N9627, N9626, N9625, N9624, N9623, N9622, N9621, N9620, N9619, N9618, N9617, N9616, N9615, N9614, N9613, N9612, N9611, N9610, N9609, N9608, N9607, N9606, N9605, N9604, N9603, N9602, N9601, N9600, N9599, N9598, N9597, N9596, N9595, N9594, N9593, N9592, N9591, N9590, N9589, N9588, N9587, N9586, N9585, N9584, N9583, N9582, N9581, N9580, N9579, N9578, N9577, N9576, N9575, N9574, N9573, N9572, N9571, N9570, N9569, N9568, N9567, N9566, N9565, N9564, N9563, N9562, N9561, N9560, N9559, N9558, N9557, N9556, N9555, N9554, N9553, N9552, N9551, N9550, N9549, N9548, N9547, N9546, N9545, N9544, N9543, N9542, N9541, N9540, N9539, N9538, N9537, N9536, N9535, N9534, N9533, N9532, N9531, N9530, N9529, N9528, N9527, N9526, N9525, N9524, N9523, N9522, N9521, N9520, N9519, N9518, N9517, N9516, N9515, N9514, N9513, N9512, N9511, N9510, N9509, N9508, N9507, N9506, N9505, N9504, N9503, N9502, N9501, N9500, N9499, N9498, N9497, N9496, N9495, N9494, N9493, N9492, N9491, N9490, N9489, N9488, N9487, N9486, N9485, N9484, N9483, N9482, N9481, N9480, N9479, N9478, N9477, N9476, N9475, N9474, N9473, N9472, N9471, N9470, N9469, N9468, N9467, N9466, N9465, N9464, N9463, N9462, N9461, N9460, N9459, N9458, N9457, N9456, N9455, N9454, N9453, N9452, N9451, N9450, N9449, N9448, N9447, N9446, N9445, N9444, N9443, N9442, N9441, N9440, N9439, N9438, N9437, N9436, N9435, N9434, N9433, N9432, N9431, N9430, N9429, N9428, N9427, N9426, N9425, N9424, N9423, N9422, N9421, N9420, N9419, N9418, N9417, N9416, N9415, N9414, N9413, N9412, N9411, N9410, N9409, N9408, N9407, N9406, N9405, N9404, N9403, N9402, N9401, N9400, N9399, N9398, N9397, N9396, N9395, N9394, N9393, N9392, N9391, N9390, N9389, N9388, N9387, N9386, N9385, N9384, N9383, N9382, N9381, N9380, N9379, N9378, N9377, N9376, N9375, N9374, N9373, N9372, N9371, N9370, N9369, N9368, N9367, N9366, N9365, N9364, N9363, N9362, N9361, N9360, N9359, N9358, N9357, N9356, N9355, N9354, N9353, N9352, N9351, N9350, N9349, N9348, N9347, N9346, N9345, N9344, N9343, N9342, N9341, N9340, N9339, N9338, N9337, N9336, N9335, N9334, N9333, N9332, N9331, N9330, N9329, N9328, N9327, N9326, N9325, N9324, N9323, N9322, N9321, N9320, N9319, N9318, N9317, N9316, N9315, N9314, N9313, N9312, N9311, N9310, N9309, N9308, N9307, N9306, N9305, N9304, N9303, N9302, N9301, N9300, N9299, N9298, N9297, N9296, N9295, N9294, N9293, N9292, N9291, N9290, N9289, N9288, N9287, N9286, N9285, N9284, N9283, N9282, N9281, N9280, N9279, N9278, N9277, N9276, N9275, N9274, N9273, N9272, N9271, N9270, N9269, N9268, N9267, N9266, N9265, N9264, N9263, N9262, N9261, N9260, N9259, N9258, N9257, N9256, N9255, N9254, N9253, N9252, N9251, N9250, N9249, N9248, N9247, N9246, N9245, N9244, N9243, N9242, N9241, N9240, N9239, N9238, N9237, N9236, N9235, N9234, N9233, N9232, N9231, N9230, N9229, N9228, N9227, N9226, N9225, N9224, N9223, N9222, N9221, N9220, N9219, N9218, N9217, N9216, N9215, N9214, N9213, N9212, N9211, N9210, N9209, N9208, N9207, N9206, N9205, N9204, N9203, N9202, N9201, N9200, N9199, N9198, N9197, N9196, N9195, N9194, N9193, N9192, N9191, N9190, N9189, N9188, N9187, N9186, N9185, N9184, N9183, N9182, N9181, N9180, N9179, N9178, N9177, N9176, N9175, N9174, N9173, N9172, N9171, N9170, N9169, N9168, N9167, N9166, N9165, N9164, N9163, N9162, N9161, N9160, N9159, N9158, N9157, N9156, N9155, N9154, N9153, N9152, N9151, N9150, N9149, N9148, N9147, N9146, N9145, N9144, N9143, N9142, N9141, N9140, N9139, N9138, N9137, N9136, N9135, N9134, N9133, N9132, N9131, N9130, N9129, N9128, N9127, N9126, N9125, N9124, N9123, N9122, N9121, N9120, N9119, N9118, N9117, N9116, N9115, N9114, N9113, N9112, N9111, N9110, N9109, N9108, N9107, N9106, N9105, N9104, N9103, N9102, N9101, N9100, N9099, N9098, N9097, N9096, N9095, N9094, N9093, N9092, N9091, N9090, N9089, N9088, N9087, N9086, N9085, N9084, N9083, N9082, N9081, N9080, N9079, N9078, N9077, N9076, N9075, N9074, N9073, N9072, N9071, N9070, N9069, N9068, N9067, N9066, N9065, N9064, N9063, N9062, N9061, N9060, N9059, N9058, N9057, N9056, N9055, N9054, N9053, N9052, N9051, N9050, N9049, N9048, N9047, N9046, N9045, N9044, N9043, N9042, N9041, N9040, N9039, N9038, N9037, N9036, N9035, N9034, N9033, N9032, N9031, N9030, N9029, N9028, N9027, N9026, N9025 } = (N167)? { N7988, N7987, N7986, N7985, N7984, N7983, N7982, N7981, N7980, N7979, N7978, N7977, N7976, N7975, N7974, N7973, N7972, N7971, N7970, N7969, N7968, N7967, N7966, N7965, N7964, N7963, N7962, N7961, N7960, N7959, N7958, N7957, N7956, N7955, N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946, N7945, N7944, N7943, N7942, N7941, N7940, N7939, N7938, N7937, N7936, N7935, N7934, N7933, N7932, N7931, N7930, N7929, N7928, N7927, N7926, N7925, N7924, N7923, N7922, N7921, N7920, N7919, N7918, N7917, N7916, N7915, N7914, N7913, N7912, N7911, N7910, N7909, N7908, N7907, N7906, N7905, N7904, N7903, N7902, N7901, N7900, N7899, N7898, N7897, N7896, N7895, N7894, N7893, N7892, N7891, N7890, N7889, N7888, N7887, N7886, N7885, N7884, N7883, N7882, N7881, N7880, N7879, N7878, N7877, N7876, N7875, N7874, N7873, N7872, N7871, N7870, N7869, N7868, N7867, N7866, N7865, N7864, N7863, N7862, N7861, N7860, N7859, N7858, N7857, N7856, N7855, N7854, N7853, N7852, N7851, N7850, N7849, N7848, N7847, N7846, N7845, N7844, N7843, N7842, N7841, N7840, N7839, N7838, N7837, N7836, N7835, N7834, N7833, N7832, N7831, N7830, N7829, N7828, N7827, N7826, N7825, N7824, N7823, N7822, N7821, N7820, N7819, N7818, N7817, N7816, N7815, N7814, N7813, N7812, N7811, N7810, N7809, N7808, N7807, N7806, N7805, N7804, N7803, N7802, N7801, N7800, N7799, N7798, N7797, N7796, N7795, N7794, N7793, N7792, N7791, N7790, N7789, N7788, N7787, N7786, N7785, N7784, N7783, N7782, N7781, N7780, N7779, N7778, N7777, N7776, N7775, N7774, N7773, N7772, N7771, N7770, N7769, N7768, N7767, N7766, N7765, N7764, N7763, N7762, N7761, N7760, N7759, N7758, N7757, N7756, N7755, N7754, N7753, N7752, N7751, N7750, N7749, N7748, N7747, N7746, N7745, N7744, N7743, N7742, N7741, N7740, N7739, N7738, N7737, N7736, N7735, N7734, N7733, N7732, N7731, N7730, N7729, N7728, N7727, N7726, N7725, N7724, N7723, N7722, N7721, N7720, N7719, N7718, N7717, N7716, N7715, N7714, N7713, N7712, N7711, N7710, N7709, N7708, N7707, N7706, N7705, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696, N7695, N7694, N7693, N7692, N7691, N7690, N7689, N7688, N7687, N7686, N7685, N7684, N7683, N7682, N7681, N7680, N7679, N7678, N7677, N7676, N7675, N7674, N7673, N7672, N7671, N7670, N7669, N7668, N7667, N7666, N7665, N7664, N7663, N7662, N7661, N7660, N7659, N7658, N7657, N7656, N7655, N7654, N7653, N7652, N7651, N7650, N7649, N7648, N7647, N7646, N7645, N7644, N7643, N7642, N7641, N7640, N7639, N7638, N7637, N7636, N7635, N7634, N7633, N7632, N7631, N7630, N7629, N7628, N7627, N7626, N7625, N7624, N7623, N7622, N7621, N7620, N7619, N7618, N7617, N7616, N7615, N7614, N7613, N7612, N7611, N7610, N7609, N7608, N7607, N7606, N7605, N7604, N7603, N7602, N7601, N7600, N7599, N7598, N7597, N7596, N7595, N7594, N7593, N7592, N7591, N7590, N7589, N7588, N7587, N7586, N7585, N7584, N7583, N7582, N7581, N7580, N7579, N7578, N7577, N7576, N7575, N7574, N7573, N7572, N7571, N7570, N7569, N7568, N7567, N7566, N7565, N7564, N7563, N7562, N7561, N7560, N7559, N7558, N7557, N7556, N7555, N7554, N7553, N7552, N7551, N7550, N7549, N7548, N7547, N7546, N7545, N7544, N7543, N7542, N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534, N7533, N7532, N7531, N7530, N7529, N7528, N7527, N7526, N7525, N7524, N7523, N7522, N7521, N7520, N7519, N7518, N7517, N7516, N7515, N7514, N7513, N7512, N7511, N7510, N7509, N7508, N7507, N7506, N7505, N7504, N7503, N7502, N7501, N7500, N7499, N7498, N7497, N7496, N7495, N7494, N7493, N7492, N7491, N7490, N7489, N7488, N7487, N7486, N7485, N7484, N7483, N7482, N7481, N7480, N7479, N7478, N7477, N7476, N7475, N7474, N7473, N7472, N7471, N7470, N7469, N7468, N7467, N7466, N7465, N7464, N7463, N7462, N7461, N7460, N7459, N7458, N7457, N7456, N7455, N7454, N7453, N7452, N7451, N7450, N7449, N7448, N7447, N7446, N7445, N7444, N7443, N7442, N7441, N7440, N7439, N7438, N7437, N7436, N7435, N7434, N7433, N7432, N7431, N7430, N7429, N7428, N7427, N7426, N7425, N7424, N7423, N7422, N7421, N7420, N7419, N7418, N7417, N7416, N7415, N7414, N7413, N7412, N7411, N7410, N7409, N7408, N7407, N7406, N7405, N7404, N7403, N7402, N7401, N7400, N7399, N7398, N7397, N7396, N7395, N7394, N7393, N7392, N7391, N7390, N7389, N7388, N7387, N7386, N7385, N7384, N7383, N7382, N7381, N7380, N7379, N7378, N7377, N7376, N7375, N7374, N7373, N7372, N7371, N7370, N7369, N7368, N7367, N7366, N7365, N7364, N7363, N7362, N7361, N7360, N7359, N7358, N7357, N7356, N7355, N7354, N7353, N7352, N7351, N7350, N7349, N7348, N7347, N7346, N7345, N7344, N7343, N7342, N7341, N7340, N7339, N7338, N7337, N7336, N7335, N7334, N7333, N7332, N7331, N7330, N7329, N7328, N7327, N7326, N7325, N7324, N7323, N7322, N7321, N7320, N7319, N7318, N7317, N7316, N7315, N7314, N7313, N7312, N7311, N7310, N7309, N7308, N7307, N7306, N7305, N7304, N7303, N7302, N7301, N7300, N7299, N7298, N7297, N7296, N7295, N7294, N7293, N7292, N7291, N7290, N7289, N7288, N7287, N7286, N7285, N7284, N7283, N7282, N7281, N7280, N7279, N7278, N7277, N7276, N7275, N7274, N7273, N7272, N7271, N7270, N7269, N7268, N7267, N7266, N7265, N7264, N7263, N7262, N7261, N7260, N7259, N7258, N7257, N7256, N7255, N7254, N7253, N7252, N7251, N7250, N7249, N7248, N7247, N7246, N7245, N7244, N7243, N7242, N7241, N7240, N7239, N7238, N7237, N7236, N7235, N7234, N7233, N7232, N7231, N7230, N7229, N7228, N7227, N7226, N7225, N7224, N7223, N7222, N7221, N7220, N7219, N7218, N7217, N7216, N7215, N7214, N7213, N7212, N7211, N7210, N7209, N7208, N7207, N7206, N7205, N7204, N7203, N7202, N7201, N7200, N7199, N7198, N7197, N7196, N7195, N7194, N7193, N7192, N7191, N7190, N7189, N7188, N7187, N7186, N7185, N7184, N7183, N7182, N7181, N7180, N7179, N7178, N7177, N7176, N7175, N7174, N7173, N7172, N7171, N7170, N7169, N7168, N7167, N7166, N7165, N7164, N7163, N7162, N7161, N7160, N7159, N7158, N7157, N7156, N7155, N7154, N7153, N7152, N7151, N7150, N7149, N7148, N7147, N7146, N7145, N7144, N7143, N7142, N7141, N7140, N7139, N7138, N7137, N7136, N7135, N7134, N7133, N7132, N7131, N7130, N7129, N7128, N7127, N7126, N7125, N7124, N7123, N7122, N7121, N7120, N7119, N7118, N7117, N7116, N7115, N7114, N7113, N7112, N7111, N7110, N7109, N7108, N7107, N7106, N7105, N7104, N7103, N7102, N7101, N7100, N7099, N7098, N7097, N7096, N7095, N7094, N7093, N7092, N7091, N7090, N7089, N7088, N7087, N7086, N7085, N7084, N7083, N7082, N7081, N7080, N7079, N7078, N7077, N7076, N7075, N7074, N7073, N7072, N7071, N7070, N7069, N7068, N7067, N7066, N7065, N7064, N7063, N7062, N7061, N7060, N7059, N7058, N7057, N7056, N7055, N7054, N7053, N7052, N7051, N7050, N7049, N7048, N7047, N7046, N7045, N7044, N7043, N7042, N7041, N7040, N7039, N7038, N7037, N7036, N7035, N7034, N7033, N7032, N7031, N7030, N7029, N7028, N7027, N7026, N7025, N7024, N7023, N7022, N7021, N7020, N7019, N7018, N7017, N7016, N7015, N7014, N7013, N7012, N7011, N7010, N7009, N7008, N7007, N7006, N7005, N7004, N7003, N7002, N7001, N7000, N6999, N6998, N6997, N6996, N6995, N6994, N6993, N6992, N6991, N6990, N6989, N6988, N6987, N6986, N6985, N6984, N6983, N6982, N6981, N6980, N6979, N6978, N6977, N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, N6957 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               (N6956)? { N9024, N9023, N9022, N9021, N9020, N9019, N9018, N9017, N9016, N9015, N9014, N9013, N9012, N9011, N9010, N9009, N9008, N9007, N9006, N9005, N9004, N9003, N9002, N9001, N9000, N8999, N8998, N8997, N8996, N8995, N8994, N8993, N8992, N8991, N8990, N8989, N8988, N8987, N8986, N8985, N8984, N8983, N8982, N8981, N8980, N8979, N8978, N8977, N8976, N8975, N8974, N8973, N8972, N8971, N8970, N8969, N8968, N8967, N8966, N8965, N8964, N8963, N8962, N8961, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719, N5718, N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691, N8960, N8959, N8958, N8957, N8956, N8955, N8954, N8953, N8952, N8951, N8950, N8949, N8948, N8947, N8946, N8945, N8944, N8943, N8942, N8941, N8940, N8939, N8938, N8937, N8936, N8935, N8934, N8933, N8932, N8931, N8930, N8929, N8928, N8927, N8926, N8925, N8924, N8923, N8922, N8921, N8920, N8919, N8918, N8917, N8916, N8915, N8914, N8913, N8912, N8911, N8910, N8909, N8908, N8907, N8906, N8905, N8904, N8903, N8902, N8901, N8900, N8899, N8898, N8897, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458, N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432, N8896, N8895, N8894, N8893, N8892, N8891, N8890, N8889, N8888, N8887, N8886, N8885, N8884, N8883, N8882, N8881, N8880, N8879, N8878, N8877, N8876, N8875, N8874, N8873, N8872, N8871, N8870, N8869, N8868, N8867, N8866, N8865, N8864, N8863, N8862, N8861, N8860, N8859, N8858, N8857, N8856, N8855, N8854, N8853, N8852, N8851, N8850, N8849, N8848, N8847, N8846, N8845, N8844, N8843, N8842, N8841, N8840, N8839, N8838, N8837, N8836, N8835, N8834, N8833, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N8832, N8831, N8830, N8829, N8828, N8827, N8826, N8825, N8824, N8823, N8822, N8821, N8820, N8819, N8818, N8817, N8816, N8815, N8814, N8813, N8812, N8811, N8810, N8809, N8808, N8807, N8806, N8805, N8804, N8803, N8802, N8801, N8800, N8799, N8798, N8797, N8796, N8795, N8794, N8793, N8792, N8791, N8790, N8789, N8788, N8787, N8786, N8785, N8784, N8783, N8782, N8781, N8780, N8779, N8778, N8777, N8776, N8775, N8774, N8773, N8772, N8771, N8770, N8769, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N8768, N8767, N8766, N8765, N8764, N8763, N8762, N8761, N8760, N8759, N8758, N8757, N8756, N8755, N8754, N8753, N8752, N8751, N8750, N8749, N8748, N8747, N8746, N8745, N8744, N8743, N8742, N8741, N8740, N8739, N8738, N8737, N8736, N8735, N8734, N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N8704, N8703, N8702, N8701, N8700, N8699, N8698, N8697, N8696, N8695, N8694, N8693, N8692, N8691, N8690, N8689, N8688, N8687, N8686, N8685, N8684, N8683, N8682, N8681, N8680, N8679, N8678, N8677, N8676, N8675, N8674, N8673, N8672, N8671, N8670, N8669, N8668, N8667, N8666, N8665, N8664, N8663, N8662, N8661, N8660, N8659, N8658, N8657, N8656, N8655, N8654, N8653, N8652, N8651, N8650, N8649, N8648, N8647, N8646, N8645, N8644, N8643, N8642, N8641, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N8640, N8639, N8638, N8637, N8636, N8635, N8634, N8633, N8632, N8631, N8630, N8629, N8628, N8627, N8626, N8625, N8624, N8623, N8622, N8621, N8620, N8619, N8618, N8617, N8616, N8615, N8614, N8613, N8612, N8611, N8610, N8609, N8608, N8607, N8606, N8605, N8604, N8603, N8602, N8601, N8600, N8599, N8598, N8597, N8596, N8595, N8594, N8593, N8592, N8591, N8590, N8589, N8588, N8587, N8586, N8585, N8584, N8583, N8582, N8581, N8580, N8579, N8578, N8577, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N8576, N8575, N8574, N8573, N8572, N8571, N8570, N8569, N8568, N8567, N8566, N8565, N8564, N8563, N8562, N8561, N8560, N8559, N8558, N8557, N8556, N8555, N8554, N8553, N8552, N8551, N8550, N8549, N8548, N8547, N8546, N8545, N8544, N8543, N8542, N8541, N8540, N8539, N8538, N8537, N8536, N8535, N8534, N8533, N8532, N8531, N8530, N8529, N8528, N8527, N8526, N8525, N8524, N8523, N8522, N8521, N8520, N8519, N8518, N8517, N8516, N8515, N8514, N8513, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878 } : 1'b0;
  assign N167 = ex_i[0];
  assign { N12120, N12119, N12118, N12117, N12116, N12115, N12114, N12113, N12112, N12111, N12110, N12109, N12108, N12107, N12106, N12105, N12104, N12103, N12102, N12101, N12100, N12099, N12098, N12097, N12096, N12095, N12094, N12093, N12092, N12091, N12090, N12089, N12088, N12087, N12086, N12085, N12084, N12083, N12082, N12081, N12080, N12079, N12078, N12077, N12076, N12075, N12074, N12073, N12072, N12071, N12070, N12069, N12068, N12067, N12066, N12065, N12064, N12063, N12062, N12061, N12060, N12059, N12058, N12057, N12056, N12055, N12054, N12053, N12052, N12051, N12050, N12049, N12048, N12047, N12046, N12045, N12044, N12043, N12042, N12041, N12040, N12039, N12038, N12037, N12036, N12035, N12034, N12033, N12032, N12031, N12030, N12029, N12028, N12027, N12026, N12025, N12024, N12023, N12022, N12021, N12020, N12019, N12018, N12017, N12016, N12015, N12014, N12013, N12012, N12011, N12010, N12009, N12008, N12007, N12006, N12005, N12004, N12003, N12002, N12001, N12000, N11999, N11998, N11997, N11996, N11995, N11994, N11993, N11992, N11991, N11990, N11989, N11988, N11987, N11986, N11985, N11984, N11983, N11982, N11981, N11980, N11979, N11978, N11977, N11976, N11975, N11974, N11973, N11972, N11971, N11970, N11969, N11968, N11967, N11966, N11965, N11964, N11963, N11962, N11961, N11960, N11959, N11958, N11957, N11956, N11955, N11954, N11953, N11952, N11951, N11950, N11949, N11948, N11947, N11946, N11945, N11944, N11943, N11942, N11941, N11940, N11939, N11938, N11937, N11936, N11935, N11934, N11933, N11932, N11931, N11930, N11929, N11928, N11927, N11926, N11925, N11924, N11923, N11922, N11921, N11920, N11919, N11918, N11917, N11916, N11915, N11914, N11913, N11912, N11911, N11910, N11909, N11908, N11907, N11906, N11905, N11904, N11903, N11902, N11901, N11900, N11899, N11898, N11897, N11896, N11895, N11894, N11893, N11892, N11891, N11890, N11889, N11888, N11887, N11886, N11885, N11884, N11883, N11882, N11881, N11880, N11879, N11878, N11877, N11876, N11875, N11874, N11873, N11872, N11871, N11870, N11869, N11868, N11867, N11866, N11865, N11864, N11863, N11862, N11861, N11860, N11859, N11858, N11857, N11856, N11855, N11854, N11853, N11852, N11851, N11850, N11849, N11848, N11847, N11846, N11845, N11844, N11843, N11842, N11841, N11840, N11839, N11838, N11837, N11836, N11835, N11834, N11833, N11832, N11831, N11830, N11829, N11828, N11827, N11826, N11825, N11824, N11823, N11822, N11821, N11820, N11819, N11818, N11817, N11816, N11815, N11814, N11813, N11812, N11811, N11810, N11809, N11808, N11807, N11806, N11805, N11804, N11803, N11802, N11801, N11800, N11799, N11798, N11797, N11796, N11795, N11794, N11793, N11792, N11791, N11790, N11789, N11788, N11787, N11786, N11785, N11784, N11783, N11782, N11781, N11780, N11779, N11778, N11777, N11776, N11775, N11774, N11773, N11772, N11771, N11770, N11769, N11768, N11767, N11766, N11765, N11764, N11763, N11762, N11761, N11760, N11759, N11758, N11757, N11756, N11755, N11754, N11753, N11752, N11751, N11750, N11749, N11748, N11747, N11746, N11745, N11744, N11743, N11742, N11741, N11740, N11739, N11738, N11737, N11736, N11735, N11734, N11733, N11732, N11731, N11730, N11729, N11728, N11727, N11726, N11725, N11724, N11723, N11722, N11721, N11720, N11719, N11718, N11717, N11716, N11715, N11714, N11713, N11712, N11711, N11710, N11709, N11708, N11707, N11706, N11705, N11704, N11703, N11702, N11701, N11700, N11699, N11698, N11697, N11696, N11695, N11694, N11693, N11692, N11691, N11690, N11689, N11688, N11687, N11686, N11685, N11684, N11683, N11682, N11681, N11680, N11679, N11678, N11677, N11676, N11675, N11674, N11673, N11672, N11671, N11670, N11669, N11668, N11667, N11666, N11665, N11664, N11663, N11662, N11661, N11660, N11659, N11658, N11657, N11656, N11655, N11654, N11653, N11652, N11651, N11650, N11649, N11648, N11647, N11646, N11645, N11644, N11643, N11642, N11641, N11640, N11639, N11638, N11637, N11636, N11635, N11634, N11633, N11632, N11631, N11630, N11629, N11628, N11627, N11626, N11625, N11624, N11623, N11622, N11621, N11620, N11619, N11618, N11617, N11616, N11615, N11614, N11613, N11612, N11611, N11610, N11609, N11608, N11607, N11606, N11605, N11604, N11603, N11602, N11601, N11600, N11599, N11598, N11597, N11596, N11595, N11594, N11593, N11592, N11591, N11590, N11589, N11588, N11587, N11586, N11585, N11584, N11583, N11582, N11581, N11580, N11579, N11578, N11577, N11576, N11575, N11574, N11573, N11572, N11571, N11570, N11569, N11568, N11567, N11566, N11565, N11564, N11563, N11562, N11561, N11560, N11559, N11558, N11557, N11556, N11555, N11554, N11553, N11552, N11551, N11550, N11549, N11548, N11547, N11546, N11545, N11544, N11543, N11542, N11541, N11540, N11539, N11538, N11537, N11536, N11535, N11534, N11533, N11532, N11531, N11530, N11529, N11528, N11527, N11526, N11525, N11524, N11523, N11522, N11521, N11520, N11519, N11518, N11517, N11516, N11515, N11514, N11513, N11512, N11511, N11510, N11509, N11508, N11507, N11506, N11505, N11504, N11503, N11502, N11501, N11500, N11499, N11498, N11497, N11496, N11495, N11494, N11493, N11492, N11491, N11490, N11489, N11488, N11487, N11486, N11485, N11484, N11483, N11482, N11481, N11480, N11479, N11478, N11477, N11476, N11475, N11474, N11473, N11472, N11471, N11470, N11469, N11468, N11467, N11466, N11465, N11464, N11463, N11462, N11461, N11460, N11459, N11458, N11457, N11456, N11455, N11454, N11453, N11452, N11451, N11450, N11449, N11448, N11447, N11446, N11445, N11444, N11443, N11442, N11441, N11440, N11439, N11438, N11437, N11436, N11435, N11434, N11433, N11432, N11431, N11430, N11429, N11428, N11427, N11426, N11425, N11424, N11423, N11422, N11421, N11420, N11419, N11418, N11417, N11416, N11415, N11414, N11413, N11412, N11411, N11410, N11409, N11408, N11407, N11406, N11405, N11404, N11403, N11402, N11401, N11400, N11399, N11398, N11397, N11396, N11395, N11394, N11393, N11392, N11391, N11390, N11389, N11388, N11387, N11386, N11385, N11384, N11383, N11382, N11381, N11380, N11379, N11378, N11377, N11376, N11375, N11374, N11373, N11372, N11371, N11370, N11369, N11368, N11367, N11366, N11365, N11364, N11363, N11362, N11361, N11360, N11359, N11358, N11357, N11356, N11355, N11354, N11353, N11352, N11351, N11350, N11349, N11348, N11347, N11346, N11345, N11344, N11343, N11342, N11341, N11340, N11339, N11338, N11337, N11336, N11335, N11334, N11333, N11332, N11331, N11330, N11329, N11328, N11327, N11326, N11325, N11324, N11323, N11322, N11321, N11320, N11319, N11318, N11317, N11316, N11315, N11314, N11313, N11312, N11311, N11310, N11309, N11308, N11307, N11306, N11305, N11304, N11303, N11302, N11301, N11300, N11299, N11298, N11297, N11296, N11295, N11294, N11293, N11292, N11291, N11290, N11289, N11288, N11287, N11286, N11285, N11284, N11283, N11282, N11281, N11280, N11279, N11278, N11277, N11276, N11275, N11274, N11273, N11272, N11271, N11270, N11269, N11268, N11267, N11266, N11265, N11264, N11263, N11262, N11261, N11260, N11259, N11258, N11257, N11256, N11255, N11254, N11253, N11252, N11251, N11250, N11249, N11248, N11247, N11246, N11245, N11244, N11243, N11242, N11241, N11240, N11239, N11238, N11237, N11236, N11235, N11234, N11233, N11232, N11231, N11230, N11229, N11228, N11227, N11226, N11225, N11224, N11223, N11222, N11221, N11220, N11219, N11218, N11217, N11216, N11215, N11214, N11213, N11212, N11211, N11210, N11209, N11208, N11207, N11206, N11205, N11204, N11203, N11202, N11201, N11200, N11199, N11198, N11197, N11196, N11195, N11194, N11193, N11192, N11191, N11190, N11189, N11188, N11187, N11186, N11185, N11184, N11183, N11182, N11181, N11180, N11179, N11178, N11177, N11176, N11175, N11174, N11173, N11172, N11171, N11170, N11169, N11168, N11167, N11166, N11165, N11164, N11163, N11162, N11161, N11160, N11159, N11158, N11157, N11156, N11155, N11154, N11153, N11152, N11151, N11150, N11149, N11148, N11147, N11146, N11145, N11144, N11143, N11142, N11141, N11140, N11139, N11138, N11137, N11136, N11135, N11134, N11133, N11132, N11131, N11130, N11129, N11128, N11127, N11126, N11125, N11124, N11123, N11122, N11121, N11120, N11119, N11118, N11117, N11116, N11115, N11114, N11113, N11112, N11111, N11110, N11109, N11108, N11107, N11106, N11105, N11104, N11103, N11102, N11101, N11100, N11099, N11098, N11097, N11096, N11095, N11094, N11093, N11092, N11091, N11090, N11089, N11088, N11087, N11086, N11085, N11084, N11083, N11082, N11081, N11080, N11079, N11078, N11077, N11076, N11075, N11074, N11073, N11072, N11071, N11070, N11069, N11068, N11067, N11066, N11065, N11064, N11063, N11062, N11061, N11060, N11059, N11058, N11057, N11056, N11055, N11054, N11053, N11052, N11051, N11050, N11049, N11048, N11047, N11046, N11045, N11044, N11043, N11042, N11041, N11040, N11039, N11038, N11037, N11036, N11035, N11034, N11033, N11032, N11031, N11030, N11029, N11028, N11027, N11026, N11025, N11024, N11023, N11022, N11021, N11020, N11019, N11018, N11017, N11016, N11015, N11014, N11013, N11012, N11011, N11010, N11009, N11008, N11007, N11006, N11005, N11004, N11003, N11002, N11001, N11000, N10999, N10998, N10997, N10996, N10995, N10994, N10993, N10992, N10991, N10990, N10989, N10988, N10987, N10986, N10985, N10984, N10983, N10982, N10981, N10980, N10979, N10978, N10977, N10976, N10975, N10974, N10973, N10972, N10971, N10970, N10969, N10968, N10967, N10966, N10965, N10964, N10963, N10962, N10961, N10960, N10959, N10958, N10957, N10956, N10955, N10954, N10953, N10952, N10951, N10950, N10949, N10948, N10947, N10946, N10945, N10944, N10943, N10942, N10941, N10940, N10939, N10938, N10937, N10936, N10935, N10934, N10933, N10932, N10931, N10930, N10929, N10928, N10927, N10926, N10925, N10924, N10923, N10922, N10921, N10920, N10919, N10918, N10917, N10916, N10915, N10914, N10913, N10912, N10911, N10910, N10909, N10908, N10907, N10906, N10905, N10904, N10903, N10902, N10901, N10900, N10899, N10898, N10897, N10896, N10895, N10894, N10893, N10892, N10891, N10890, N10889, N10888, N10887, N10886, N10885, N10884, N10883, N10882, N10881, N10880, N10879, N10878, N10877, N10876, N10875, N10874, N10873, N10872, N10871, N10870, N10869, N10868, N10867, N10866, N10865, N10864, N10863, N10862, N10861, N10860, N10859, N10858, N10857, N10856, N10855, N10854, N10853, N10852, N10851, N10850, N10849, N10848, N10847, N10846, N10845, N10844, N10843, N10842, N10841, N10840, N10839, N10838, N10837, N10836, N10835, N10834, N10833, N10832, N10831, N10830, N10829, N10828, N10827, N10826, N10825, N10824, N10823, N10822, N10821, N10820, N10819, N10818, N10817, N10816, N10815, N10814, N10813, N10812, N10811, N10810, N10809, N10808, N10807, N10806, N10805, N10804, N10803, N10802, N10801, N10800, N10799, N10798, N10797, N10796, N10795, N10794, N10793, N10792, N10791, N10790, N10789, N10788, N10787, N10786, N10785, N10784, N10783, N10782, N10781, N10780, N10779, N10778, N10777, N10776, N10775, N10774, N10773, N10772, N10771, N10770, N10769, N10768, N10767, N10766, N10765, N10764, N10763, N10762, N10761, N10760, N10759, N10758, N10757, N10756, N10755, N10754, N10753, N10752, N10751, N10750, N10749, N10748, N10747, N10746, N10745, N10744, N10743, N10742, N10741, N10740, N10739, N10738, N10737, N10736, N10735, N10734, N10733, N10732, N10731, N10730, N10729, N10728, N10727, N10726, N10725, N10724, N10723, N10722, N10721, N10720, N10719, N10718, N10717, N10716, N10715, N10714, N10713, N10712, N10711, N10710, N10709, N10708, N10707, N10706, N10705, N10704, N10703, N10702, N10701, N10700, N10699, N10698, N10697, N10696, N10695, N10694, N10693, N10692, N10691, N10690, N10689, N10688, N10687, N10686, N10685, N10684, N10683, N10682, N10681, N10680, N10679, N10678, N10677, N10676, N10675, N10674, N10673, N10672, N10671, N10670, N10669, N10668, N10667, N10666, N10665, N10664, N10663, N10662, N10661, N10660, N10659, N10658, N10657, N10656, N10655, N10654, N10653, N10652, N10651, N10650, N10649, N10648, N10647, N10646, N10645, N10644, N10643, N10642, N10641, N10640, N10639, N10638, N10637, N10636, N10635, N10634, N10633, N10632, N10631, N10630, N10629, N10628, N10627, N10626, N10625, N10624, N10623, N10622, N10621, N10620, N10619, N10618, N10617, N10616, N10615, N10614, N10613, N10612, N10611, N10610, N10609, N10608, N10607, N10606, N10605, N10604, N10603, N10602, N10601, N10600, N10599, N10598, N10597, N10596, N10595, N10594, N10593, N10592, N10591, N10590, N10589, N10588, N10587, N10586, N10585, N10584, N10583, N10582, N10581, N10580, N10579, N10578, N10577, N10576, N10575, N10574, N10573, N10572, N10571, N10570, N10569, N10568, N10567, N10566, N10565, N10564, N10563, N10562, N10561, N10560, N10559, N10558, N10557, N10556, N10555, N10554, N10553, N10552, N10551, N10550, N10549, N10548, N10547, N10546, N10545, N10544, N10543, N10542, N10541, N10540, N10539, N10538, N10537, N10536, N10535, N10534, N10533, N10532, N10531, N10530, N10529, N10528, N10527, N10526, N10525, N10524, N10523, N10522, N10521, N10520, N10519, N10518, N10517, N10516, N10515, N10514, N10513, N10512, N10511, N10510, N10509, N10508, N10507, N10506, N10505, N10504, N10503, N10502, N10501, N10500, N10499, N10498, N10497, N10496, N10495, N10494, N10493, N10492, N10491, N10490, N10489, N10488, N10487, N10486, N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422, N10421, N10420, N10419, N10418, N10417, N10416, N10415, N10414, N10413, N10412, N10411, N10410, N10409, N10408, N10407, N10406, N10405, N10404, N10403, N10402, N10401, N10400, N10399, N10398, N10397, N10396, N10395, N10394, N10393, N10392, N10391, N10390, N10389, N10388, N10387, N10386, N10385, N10384, N10383, N10382, N10381, N10380, N10379, N10378, N10377, N10376, N10375, N10374, N10373, N10372, N10371, N10370, N10369, N10368, N10367, N10366, N10365, N10364, N10363, N10362, N10361, N10360, N10359, N10358, N10357, N10356, N10355, N10354, N10353, N10352, N10351, N10350, N10349, N10348, N10347, N10346, N10345, N10344, N10343, N10342, N10341, N10340, N10339, N10338, N10337, N10336, N10335, N10334, N10333, N10332, N10331, N10330, N10329, N10328, N10327, N10326, N10325, N10324, N10323, N10322, N10321, N10320, N10319, N10318, N10317, N10316, N10315, N10314, N10313, N10312, N10311, N10310, N10309, N10308, N10307, N10306, N10305, N10304, N10303, N10302, N10301, N10300, N10299, N10298, N10297, N10296, N10295, N10294, N10293, N10292, N10291, N10290, N10289, N10288, N10287, N10286, N10285, N10284, N10283, N10282, N10281, N10280, N10279, N10278, N10277, N10276, N10275, N10274, N10273, N10272, N10271, N10270, N10269, N10268, N10267, N10266, N10265, N10264, N10263, N10262, N10261, N10260, N10259, N10258, N10257, N10256, N10255, N10254, N10253, N10252, N10251, N10250, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057 } = (N168)? { N6439, N6438, N6437, N6436, N6435, N6434, N6433, N6432, N6431, N6430, N6429, N6428, N6427, N6426, N6425, N6424, N6423, N6422, N6421, N6420, N6419, N6418, N6417, N6416, N6415, N6414, N6413, N6412, N6411, N6410, N6409, N6408, N6407, N6406, N6405, N6404, N6403, N6402, N6401, N6400, N6399, N6398, N6397, N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377, N6376, N5911, N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002, N10001, N10000, N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9967, N9966, N9965, N9964, N9963, N9962, N9961, N9960, N9959, N9958, N9957, N9956, N9955, N9954, N9953, N9952, N9951, N9950, N9949, N9948, N9947, N9946, N9945, N9944, N9943, N9942, N9941, N9940, N9939, N9938, N9937, N9936, N9935, N9934, N9933, N9932, N9931, N9930, N9929, N9928, N6951, N6950, N6949, N6948, N6947, N6946, N6945, N6944, N6943, N6942, N6941, N6940, N6939, N6938, N6937, N6936, N6935, N6934, N6933, N6932, N6931, N6930, N6929, N6928, N6927, N6926, N6925, N6924, N6923, N6922, N6921, N6920, N6919, N6918, N6917, N6916, N6915, N6914, N6913, N6912, N6911, N6910, N6909, N6908, N6907, N6906, N6905, N6904, N6903, N6902, N6901, N6900, N6899, N6898, N6897, N6896, N6895, N6894, N6893, N6892, N6891, N6890, N6889, N6888, N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366, N6365, N6364, N6363, N6362, N6361, N6360, N6359, N6358, N6357, N6356, N6355, N6354, N6353, N6352, N6351, N6350, N6349, N6348, N6347, N6346, N6345, N6344, N6343, N6342, N6341, N6340, N6339, N6338, N6337, N6336, N6335, N6334, N6333, N6332, N6331, N6330, N6329, N6328, N6327, N6326, N6325, N6324, N6323, N6322, N6321, N6320, N6319, N6318, N6317, N6316, N6315, N6314, N6313, N6312, N6311, N5910, N9927, N9926, N9925, N9924, N9923, N9922, N9921, N9920, N9919, N9918, N9917, N9916, N9915, N9914, N9913, N9912, N9911, N9910, N9909, N9908, N9907, N9906, N9905, N9904, N9903, N9902, N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838, N9837, N9836, N9835, N9834, N9833, N9832, N9831, N9830, N9829, N9828, N9827, N9826, N9825, N9824, N9823, N9822, N9821, N9820, N9819, N9818, N9817, N9816, N9815, N9814, N9813, N9812, N9811, N9810, N9809, N9808, N9807, N9806, N9805, N9804, N9803, N9802, N9801, N9800, N9799, N6887, N6886, N6885, N6884, N6883, N6882, N6881, N6880, N6879, N6878, N6877, N6876, N6875, N6874, N6873, N6872, N6871, N6870, N6869, N6868, N6867, N6866, N6865, N6864, N6863, N6862, N6861, N6860, N6859, N6858, N6857, N6856, N6855, N6854, N6853, N6852, N6851, N6850, N6849, N6848, N6847, N6846, N6845, N6844, N6843, N6842, N6841, N6840, N6839, N6838, N6837, N6836, N6835, N6834, N6833, N6832, N6831, N6830, N6829, N6828, N6827, N6826, N6825, N6824, N6309, N6308, N6307, N6306, N6305, N6304, N6303, N6302, N6301, N6300, N6299, N6298, N6297, N6296, N6295, N6294, N6293, N6292, N6291, N6290, N6289, N6288, N6287, N6286, N6285, N6284, N6283, N6282, N6281, N6280, N6279, N6278, N6277, N6276, N6275, N6274, N6273, N6272, N6271, N6270, N6269, N6268, N6267, N6266, N6265, N6264, N6263, N6262, N6261, N6260, N6259, N6258, N6257, N6256, N6255, N6254, N6253, N6252, N6251, N6250, N6249, N6248, N6247, N6246, N5909, N9798, N9797, N9796, N9795, N9794, N9793, N9792, N9791, N9790, N9789, N9788, N9787, N9786, N9785, N9784, N9783, N9782, N9781, N9780, N9779, N9778, N9777, N9776, N9775, N9774, N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742, N9741, N9740, N9739, N9738, N9737, N9736, N9735, N9734, N9733, N9732, N9731, N9730, N9729, N9728, N9727, N9726, N9725, N9724, N9723, N9722, N9721, N9720, N9719, N9718, N9717, N9716, N9715, N9714, N9713, N9712, N9711, N9710, N9709, N9708, N9707, N9706, N9705, N9704, N9703, N9702, N9701, N9700, N9699, N9698, N9697, N9696, N9695, N9694, N9693, N9692, N9691, N9690, N9689, N9688, N9687, N9686, N9685, N9684, N9683, N9682, N9681, N9680, N9679, N9678, N9677, N9676, N9675, N9674, N9673, N9672, N9671, N9670, N6823, N6822, N6821, N6820, N6819, N6818, N6817, N6816, N6815, N6814, N6813, N6812, N6811, N6810, N6809, N6808, N6807, N6806, N6805, N6804, N6803, N6802, N6801, N6800, N6799, N6798, N6797, N6796, N6795, N6794, N6793, N6792, N6791, N6790, N6789, N6788, N6787, N6786, N6785, N6784, N6783, N6782, N6781, N6780, N6779, N6778, N6777, N6776, N6775, N6774, N6773, N6772, N6771, N6770, N6769, N6768, N6767, N6766, N6765, N6764, N6763, N6762, N6761, N6760, N6244, N6243, N6242, N6241, N6240, N6239, N6238, N6237, N6236, N6235, N6234, N6233, N6232, N6231, N6230, N6229, N6228, N6227, N6226, N6225, N6224, N6223, N6222, N6221, N6220, N6219, N6218, N6217, N6216, N6215, N6214, N6213, N6212, N6211, N6210, N6209, N6208, N6207, N6206, N6205, N6204, N6203, N6202, N6201, N6200, N6199, N6198, N6197, N6196, N6195, N6194, N6193, N6192, N6191, N6190, N6189, N6188, N6187, N6186, N6185, N6184, N6183, N6182, N6181, N5908, N9669, N9668, N9667, N9666, N9665, N9664, N9663, N9662, N9661, N9660, N9659, N9658, N9657, N9656, N9655, N9654, N9653, N9652, N9651, N9650, N9649, N9648, N9647, N9646, N9645, N9644, N9643, N9642, N9641, N9640, N9639, N9638, N9637, N9636, N9635, N9634, N9633, N9632, N9631, N9630, N9629, N9628, N9627, N9626, N9625, N9624, N9623, N9622, N9621, N9620, N9619, N9618, N9617, N9616, N9615, N9614, N9613, N9612, N9611, N9610, N9609, N9608, N9607, N9606, N9605, N9604, N9603, N9602, N9601, N9600, N9599, N9598, N9597, N9596, N9595, N9594, N9593, N9592, N9591, N9590, N9589, N9588, N9587, N9586, N9585, N9584, N9583, N9582, N9581, N9580, N9579, N9578, N9577, N9576, N9575, N9574, N9573, N9572, N9571, N9570, N9569, N9568, N9567, N9566, N9565, N9564, N9563, N9562, N9561, N9560, N9559, N9558, N9557, N9556, N9555, N9554, N9553, N9552, N9551, N9550, N9549, N9548, N9547, N9546, N9545, N9544, N9543, N9542, N9541, N6759, N6758, N6757, N6756, N6755, N6754, N6753, N6752, N6751, N6750, N6749, N6748, N6747, N6746, N6745, N6744, N6743, N6742, N6741, N6740, N6739, N6738, N6737, N6736, N6735, N6734, N6733, N6732, N6731, N6730, N6729, N6728, N6727, N6726, N6725, N6724, N6723, N6722, N6721, N6720, N6719, N6718, N6717, N6716, N6715, N6714, N6713, N6712, N6711, N6710, N6709, N6708, N6707, N6706, N6705, N6704, N6703, N6702, N6701, N6700, N6699, N6698, N6697, N6696, N6179, N6178, N6177, N6176, N6175, N6174, N6173, N6172, N6171, N6170, N6169, N6168, N6167, N6166, N6165, N6164, N6163, N6162, N6161, N6160, N6159, N6158, N6157, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N6149, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N6141, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N6133, N6132, N6131, N6130, N6129, N6128, N6127, N6126, N6125, N6124, N6123, N6122, N6121, N6120, N6119, N6118, N6117, N6116, N5907, N9540, N9539, N9538, N9537, N9536, N9535, N9534, N9533, N9532, N9531, N9530, N9529, N9528, N9527, N9526, N9525, N9524, N9523, N9522, N9521, N9520, N9519, N9518, N9517, N9516, N9515, N9514, N9513, N9512, N9511, N9510, N9509, N9508, N9507, N9506, N9505, N9504, N9503, N9502, N9501, N9500, N9499, N9498, N9497, N9496, N9495, N9494, N9493, N9492, N9491, N9490, N9489, N9488, N9487, N9486, N9485, N9484, N9483, N9482, N9481, N9480, N9479, N9478, N9477, N9476, N9475, N9474, N9473, N9472, N9471, N9470, N9469, N9468, N9467, N9466, N9465, N9464, N9463, N9462, N9461, N9460, N9459, N9458, N9457, N9456, N9455, N9454, N9453, N9452, N9451, N9450, N9449, N9448, N9447, N9446, N9445, N9444, N9443, N9442, N9441, N9440, N9439, N9438, N9437, N9436, N9435, N9434, N9433, N9432, N9431, N9430, N9429, N9428, N9427, N9426, N9425, N9424, N9423, N9422, N9421, N9420, N9419, N9418, N9417, N9416, N9415, N9414, N9413, N9412, N6695, N6694, N6693, N6692, N6691, N6690, N6689, N6688, N6687, N6686, N6685, N6684, N6683, N6682, N6681, N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667, N6666, N6665, N6664, N6663, N6662, N6661, N6660, N6659, N6658, N6657, N6656, N6655, N6654, N6653, N6652, N6651, N6650, N6649, N6648, N6647, N6646, N6645, N6644, N6643, N6642, N6641, N6640, N6639, N6638, N6637, N6636, N6635, N6634, N6633, N6632, N6114, N6113, N6112, N6111, N6110, N6109, N6108, N6107, N6106, N6105, N6104, N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, N6093, N6092, N6091, N6090, N6089, N6088, N6087, N6086, N6085, N6084, N6083, N6082, N6081, N6080, N6079, N6078, N6077, N6076, N6075, N6074, N6073, N6072, N6071, N6070, N6069, N6068, N6067, N6066, N6065, N6064, N6063, N6062, N6061, N6060, N6059, N6058, N6057, N6056, N6055, N6054, N6053, N6052, N6051, N5906, N9411, N9410, N9409, N9408, N9407, N9406, N9405, N9404, N9403, N9402, N9401, N9400, N9399, N9398, N9397, N9396, N9395, N9394, N9393, N9392, N9391, N9390, N9389, N9388, N9387, N9386, N9385, N9384, N9383, N9382, N9381, N9380, N9379, N9378, N9377, N9376, N9375, N9374, N9373, N9372, N9371, N9370, N9369, N9368, N9367, N9366, N9365, N9364, N9363, N9362, N9361, N9360, N9359, N9358, N9357, N9356, N9355, N9354, N9353, N9352, N9351, N9350, N9349, N9348, N9347, N9346, N9345, N9344, N9343, N9342, N9341, N9340, N9339, N9338, N9337, N9336, N9335, N9334, N9333, N9332, N9331, N9330, N9329, N9328, N9327, N9326, N9325, N9324, N9323, N9322, N9321, N9320, N9319, N9318, N9317, N9316, N9315, N9314, N9313, N9312, N9311, N9310, N9309, N9308, N9307, N9306, N9305, N9304, N9303, N9302, N9301, N9300, N9299, N9298, N9297, N9296, N9295, N9294, N9293, N9292, N9291, N9290, N9289, N9288, N9287, N9286, N9285, N9284, N9283, N6631, N6630, N6629, N6628, N6627, N6626, N6625, N6624, N6623, N6622, N6621, N6620, N6619, N6618, N6617, N6616, N6615, N6614, N6613, N6612, N6611, N6610, N6609, N6608, N6607, N6606, N6605, N6604, N6603, N6602, N6601, N6600, N6599, N6598, N6597, N6596, N6595, N6594, N6593, N6592, N6591, N6590, N6589, N6588, N6587, N6586, N6585, N6584, N6583, N6582, N6581, N6580, N6579, N6578, N6577, N6576, N6575, N6574, N6573, N6572, N6571, N6570, N6569, N6568, N6049, N6048, N6047, N6046, N6045, N6044, N6043, N6042, N6041, N6040, N6039, N6038, N6037, N6036, N6035, N6034, N6033, N6032, N6031, N6030, N6029, N6028, N6027, N6026, N6025, N6024, N6023, N6022, N6021, N6020, N6019, N6018, N6017, N6016, N6015, N6014, N6013, N6012, N6011, N6010, N6009, N6008, N6007, N6006, N6005, N6004, N6003, N6002, N6001, N6000, N5999, N5998, N5997, N5996, N5995, N5994, N5993, N5992, N5991, N5990, N5989, N5988, N5987, N5986, N5905, N9282, N9281, N9280, N9279, N9278, N9277, N9276, N9275, N9274, N9273, N9272, N9271, N9270, N9269, N9268, N9267, N9266, N9265, N9264, N9263, N9262, N9261, N9260, N9259, N9258, N9257, N9256, N9255, N9254, N9253, N9252, N9251, N9250, N9249, N9248, N9247, N9246, N9245, N9244, N9243, N9242, N9241, N9240, N9239, N9238, N9237, N9236, N9235, N9234, N9233, N9232, N9231, N9230, N9229, N9228, N9227, N9226, N9225, N9224, N9223, N9222, N9221, N9220, N9219, N9218, N9217, N9216, N9215, N9214, N9213, N9212, N9211, N9210, N9209, N9208, N9207, N9206, N9205, N9204, N9203, N9202, N9201, N9200, N9199, N9198, N9197, N9196, N9195, N9194, N9193, N9192, N9191, N9190, N9189, N9188, N9187, N9186, N9185, N9184, N9183, N9182, N9181, N9180, N9179, N9178, N9177, N9176, N9175, N9174, N9173, N9172, N9171, N9170, N9169, N9168, N9167, N9166, N9165, N9164, N9163, N9162, N9161, N9160, N9159, N9158, N9157, N9156, N9155, N9154, N6567, N6566, N6565, N6564, N6563, N6562, N6561, N6560, N6559, N6558, N6557, N6556, N6555, N6554, N6553, N6552, N6551, N6550, N6549, N6548, N6547, N6546, N6545, N6544, N6543, N6542, N6541, N6540, N6539, N6538, N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530, N6529, N6528, N6527, N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, N6518, N6517, N6516, N6515, N6514, N6513, N6512, N6511, N6510, N6509, N6508, N6507, N6506, N6505, N6504, N5984, N5983, N5982, N5981, N5980, N5979, N5978, N5977, N5976, N5975, N5974, N5973, N5972, N5971, N5970, N5969, N5968, N5967, N5966, N5965, N5964, N5963, N5962, N5961, N5960, N5959, N5958, N5957, N5956, N5955, N5954, N5953, N5952, N5951, N5950, N5949, N5948, N5947, N5946, N5945, N5944, N5943, N5942, N5941, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N5932, N5931, N5930, N5929, N5928, N5927, N5926, N5925, N5924, N5923, N5922, N5921, N5904, N9153, N9152, N9151, N9150, N9149, N9148, N9147, N9146, N9145, N9144, N9143, N9142, N9141, N9140, N9139, N9138, N9137, N9136, N9135, N9134, N9133, N9132, N9131, N9130, N9129, N9128, N9127, N9126, N9125, N9124, N9123, N9122, N9121, N9120, N9119, N9118, N9117, N9116, N9115, N9114, N9113, N9112, N9111, N9110, N9109, N9108, N9107, N9106, N9105, N9104, N9103, N9102, N9101, N9100, N9099, N9098, N9097, N9096, N9095, N9094, N9093, N9092, N9091, N9090, N9089, N9088, N9087, N9086, N9085, N9084, N9083, N9082, N9081, N9080, N9079, N9078, N9077, N9076, N9075, N9074, N9073, N9072, N9071, N9070, N9069, N9068, N9067, N9066, N9065, N9064, N9063, N9062, N9061, N9060, N9059, N9058, N9057, N9056, N9055, N9054, N9053, N9052, N9051, N9050, N9049, N9048, N9047, N9046, N9045, N9044, N9043, N9042, N9041, N9040, N9039, N9038, N9037, N9036, N9035, N9034, N9033, N9032, N9031, N9030, N9029, N9028, N9027, N9026, N9025, N6503, N6502, N6501, N6500, N6499, N6498, N6497, N6496, N6495, N6494, N6493, N6492, N6491, N6490, N6489, N6488, N6487, N6486, N6485, N6484, N6483, N6482, N6481, N6480, N6479, N6478, N6477, N6476, N6475, N6474, N6473, N6472, N6471, N6470, N6469, N6468, N6467, N6466, N6465, N6464, N6463, N6462, N6461, N6460, N6459, N6458, N6457, N6456, N6455, N6454, N6453, N6452, N6451, N6450, N6449, N6448, N6447, N6446, N6445, N6444, N6443, N6442, N6441, N6440 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5903)? { N5884, N5883, N5882, N5881, N5880, N5879, N5878, N5877, N5876, N5875, N5874, N5873, N5872, N5871, N5870, N5869, N5868, N5867, N5866, N5865, N5864, N5863, N5862, N5861, N5860, N5859, N5858, N5857, N5856, N5855, N5854, N5853, N5852, N5851, N5850, N5849, N5848, N5847, N5846, N5845, N5844, N5843, N5842, N5841, N5840, N5839, N5838, N5837, N5836, N5835, N5834, N5833, N5832, N5831, N5830, N5829, N5828, N5827, N5826, N5825, N5824, N5823, N5822, N5821, N5820, N5819, N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719, N5718, N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691, N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654, N5653, N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627, N5625, N5624, N5623, N5622, N5621, N5620, N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588, N5587, N5586, N5585, N5584, N5583, N5582, N5581, N5580, N5579, N5578, N5577, N5576, N5575, N5574, N5573, N5572, N5571, N5570, N5569, N5568, N5567, N5566, N5565, N5564, N5563, N5562, N5561, N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458, N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, N5418, N5417, N5416, N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073, N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814 } : 1'b0;
  assign N168 = N5902;
  assign N12139 = (N169)? 1'b1 : 
                  (N12155)? N10250 : 1'b0;
  assign N169 = N12147;
  assign N12140 = (N170)? 1'b1 : 
                  (N12220)? N10508 : 1'b0;
  assign N170 = N12148;
  assign N12141 = (N171)? 1'b1 : 
                  (N12285)? N10766 : 1'b0;
  assign N171 = N12149;
  assign N12142 = (N172)? 1'b1 : 
                  (N12350)? N11024 : 1'b0;
  assign N172 = N12150;
  assign N12143 = (N173)? 1'b1 : 
                  (N12415)? N11282 : 1'b0;
  assign N173 = N12151;
  assign N12144 = (N174)? 1'b1 : 
                  (N12480)? N11540 : 1'b0;
  assign N174 = N12152;
  assign N12145 = (N175)? 1'b1 : 
                  (N12545)? N11798 : 1'b0;
  assign N175 = N12153;
  assign N12146 = (N176)? 1'b1 : 
                  (N12610)? N12056 : 1'b0;
  assign N176 = N12154;
  assign { N12219, N12218, N12217, N12216, N12215, N12214, N12213, N12212, N12211, N12210, N12209, N12208, N12207, N12206, N12205, N12204, N12203, N12202, N12201, N12200, N12199, N12198, N12197, N12196, N12195, N12194, N12193, N12192, N12191, N12190, N12189, N12188, N12187, N12186, N12185, N12184, N12183, N12182, N12181, N12180, N12179, N12178, N12177, N12176, N12175, N12174, N12173, N12172, N12171, N12170, N12169, N12168, N12167, N12166, N12165, N12164, N12163, N12162, N12161, N12160, N12159, N12158, N12157, N12156 } = (N169)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12155)? { N10314, N10313, N10312, N10311, N10310, N10309, N10308, N10307, N10306, N10305, N10304, N10303, N10302, N10301, N10300, N10299, N10298, N10297, N10296, N10295, N10294, N10293, N10292, N10291, N10290, N10289, N10288, N10287, N10286, N10285, N10284, N10283, N10282, N10281, N10280, N10279, N10278, N10277, N10276, N10275, N10274, N10273, N10272, N10271, N10270, N10269, N10268, N10267, N10266, N10265, N10264, N10263, N10262, N10261, N10260, N10259, N10258, N10257, N10256, N10255, N10254, N10253, N10252, N10251 } : 1'b0;
  assign { N12284, N12283, N12282, N12281, N12280, N12279, N12278, N12277, N12276, N12275, N12274, N12273, N12272, N12271, N12270, N12269, N12268, N12267, N12266, N12265, N12264, N12263, N12262, N12261, N12260, N12259, N12258, N12257, N12256, N12255, N12254, N12253, N12252, N12251, N12250, N12249, N12248, N12247, N12246, N12245, N12244, N12243, N12242, N12241, N12240, N12239, N12238, N12237, N12236, N12235, N12234, N12233, N12232, N12231, N12230, N12229, N12228, N12227, N12226, N12225, N12224, N12223, N12222, N12221 } = (N170)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12220)? { N10572, N10571, N10570, N10569, N10568, N10567, N10566, N10565, N10564, N10563, N10562, N10561, N10560, N10559, N10558, N10557, N10556, N10555, N10554, N10553, N10552, N10551, N10550, N10549, N10548, N10547, N10546, N10545, N10544, N10543, N10542, N10541, N10540, N10539, N10538, N10537, N10536, N10535, N10534, N10533, N10532, N10531, N10530, N10529, N10528, N10527, N10526, N10525, N10524, N10523, N10522, N10521, N10520, N10519, N10518, N10517, N10516, N10515, N10514, N10513, N10512, N10511, N10510, N10509 } : 1'b0;
  assign { N12349, N12348, N12347, N12346, N12345, N12344, N12343, N12342, N12341, N12340, N12339, N12338, N12337, N12336, N12335, N12334, N12333, N12332, N12331, N12330, N12329, N12328, N12327, N12326, N12325, N12324, N12323, N12322, N12321, N12320, N12319, N12318, N12317, N12316, N12315, N12314, N12313, N12312, N12311, N12310, N12309, N12308, N12307, N12306, N12305, N12304, N12303, N12302, N12301, N12300, N12299, N12298, N12297, N12296, N12295, N12294, N12293, N12292, N12291, N12290, N12289, N12288, N12287, N12286 } = (N171)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12285)? { N10830, N10829, N10828, N10827, N10826, N10825, N10824, N10823, N10822, N10821, N10820, N10819, N10818, N10817, N10816, N10815, N10814, N10813, N10812, N10811, N10810, N10809, N10808, N10807, N10806, N10805, N10804, N10803, N10802, N10801, N10800, N10799, N10798, N10797, N10796, N10795, N10794, N10793, N10792, N10791, N10790, N10789, N10788, N10787, N10786, N10785, N10784, N10783, N10782, N10781, N10780, N10779, N10778, N10777, N10776, N10775, N10774, N10773, N10772, N10771, N10770, N10769, N10768, N10767 } : 1'b0;
  assign { N12414, N12413, N12412, N12411, N12410, N12409, N12408, N12407, N12406, N12405, N12404, N12403, N12402, N12401, N12400, N12399, N12398, N12397, N12396, N12395, N12394, N12393, N12392, N12391, N12390, N12389, N12388, N12387, N12386, N12385, N12384, N12383, N12382, N12381, N12380, N12379, N12378, N12377, N12376, N12375, N12374, N12373, N12372, N12371, N12370, N12369, N12368, N12367, N12366, N12365, N12364, N12363, N12362, N12361, N12360, N12359, N12358, N12357, N12356, N12355, N12354, N12353, N12352, N12351 } = (N172)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12350)? { N11088, N11087, N11086, N11085, N11084, N11083, N11082, N11081, N11080, N11079, N11078, N11077, N11076, N11075, N11074, N11073, N11072, N11071, N11070, N11069, N11068, N11067, N11066, N11065, N11064, N11063, N11062, N11061, N11060, N11059, N11058, N11057, N11056, N11055, N11054, N11053, N11052, N11051, N11050, N11049, N11048, N11047, N11046, N11045, N11044, N11043, N11042, N11041, N11040, N11039, N11038, N11037, N11036, N11035, N11034, N11033, N11032, N11031, N11030, N11029, N11028, N11027, N11026, N11025 } : 1'b0;
  assign { N12479, N12478, N12477, N12476, N12475, N12474, N12473, N12472, N12471, N12470, N12469, N12468, N12467, N12466, N12465, N12464, N12463, N12462, N12461, N12460, N12459, N12458, N12457, N12456, N12455, N12454, N12453, N12452, N12451, N12450, N12449, N12448, N12447, N12446, N12445, N12444, N12443, N12442, N12441, N12440, N12439, N12438, N12437, N12436, N12435, N12434, N12433, N12432, N12431, N12430, N12429, N12428, N12427, N12426, N12425, N12424, N12423, N12422, N12421, N12420, N12419, N12418, N12417, N12416 } = (N173)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12415)? { N11346, N11345, N11344, N11343, N11342, N11341, N11340, N11339, N11338, N11337, N11336, N11335, N11334, N11333, N11332, N11331, N11330, N11329, N11328, N11327, N11326, N11325, N11324, N11323, N11322, N11321, N11320, N11319, N11318, N11317, N11316, N11315, N11314, N11313, N11312, N11311, N11310, N11309, N11308, N11307, N11306, N11305, N11304, N11303, N11302, N11301, N11300, N11299, N11298, N11297, N11296, N11295, N11294, N11293, N11292, N11291, N11290, N11289, N11288, N11287, N11286, N11285, N11284, N11283 } : 1'b0;
  assign { N12544, N12543, N12542, N12541, N12540, N12539, N12538, N12537, N12536, N12535, N12534, N12533, N12532, N12531, N12530, N12529, N12528, N12527, N12526, N12525, N12524, N12523, N12522, N12521, N12520, N12519, N12518, N12517, N12516, N12515, N12514, N12513, N12512, N12511, N12510, N12509, N12508, N12507, N12506, N12505, N12504, N12503, N12502, N12501, N12500, N12499, N12498, N12497, N12496, N12495, N12494, N12493, N12492, N12491, N12490, N12489, N12488, N12487, N12486, N12485, N12484, N12483, N12482, N12481 } = (N174)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12480)? { N11604, N11603, N11602, N11601, N11600, N11599, N11598, N11597, N11596, N11595, N11594, N11593, N11592, N11591, N11590, N11589, N11588, N11587, N11586, N11585, N11584, N11583, N11582, N11581, N11580, N11579, N11578, N11577, N11576, N11575, N11574, N11573, N11572, N11571, N11570, N11569, N11568, N11567, N11566, N11565, N11564, N11563, N11562, N11561, N11560, N11559, N11558, N11557, N11556, N11555, N11554, N11553, N11552, N11551, N11550, N11549, N11548, N11547, N11546, N11545, N11544, N11543, N11542, N11541 } : 1'b0;
  assign { N12609, N12608, N12607, N12606, N12605, N12604, N12603, N12602, N12601, N12600, N12599, N12598, N12597, N12596, N12595, N12594, N12593, N12592, N12591, N12590, N12589, N12588, N12587, N12586, N12585, N12584, N12583, N12582, N12581, N12580, N12579, N12578, N12577, N12576, N12575, N12574, N12573, N12572, N12571, N12570, N12569, N12568, N12567, N12566, N12565, N12564, N12563, N12562, N12561, N12560, N12559, N12558, N12557, N12556, N12555, N12554, N12553, N12552, N12551, N12550, N12549, N12548, N12547, N12546 } = (N175)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12545)? { N11862, N11861, N11860, N11859, N11858, N11857, N11856, N11855, N11854, N11853, N11852, N11851, N11850, N11849, N11848, N11847, N11846, N11845, N11844, N11843, N11842, N11841, N11840, N11839, N11838, N11837, N11836, N11835, N11834, N11833, N11832, N11831, N11830, N11829, N11828, N11827, N11826, N11825, N11824, N11823, N11822, N11821, N11820, N11819, N11818, N11817, N11816, N11815, N11814, N11813, N11812, N11811, N11810, N11809, N11808, N11807, N11806, N11805, N11804, N11803, N11802, N11801, N11800, N11799 } : 1'b0;
  assign { N12674, N12673, N12672, N12671, N12670, N12669, N12668, N12667, N12666, N12665, N12664, N12663, N12662, N12661, N12660, N12659, N12658, N12657, N12656, N12655, N12654, N12653, N12652, N12651, N12650, N12649, N12648, N12647, N12646, N12645, N12644, N12643, N12642, N12641, N12640, N12639, N12638, N12637, N12636, N12635, N12634, N12633, N12632, N12631, N12630, N12629, N12628, N12627, N12626, N12625, N12624, N12623, N12622, N12621, N12620, N12619, N12618, N12617, N12616, N12615, N12614, N12613, N12612, N12611 } = (N176)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12610)? { N12120, N12119, N12118, N12117, N12116, N12115, N12114, N12113, N12112, N12111, N12110, N12109, N12108, N12107, N12106, N12105, N12104, N12103, N12102, N12101, N12100, N12099, N12098, N12097, N12096, N12095, N12094, N12093, N12092, N12091, N12090, N12089, N12088, N12087, N12086, N12085, N12084, N12083, N12082, N12081, N12080, N12079, N12078, N12077, N12076, N12075, N12074, N12073, N12072, N12071, N12070, N12069, N12068, N12067, N12066, N12065, N12064, N12063, N12062, N12061, N12060, N12059, N12058, N12057 } : 1'b0;
  assign { N12738, N12737, N12736, N12735, N12734, N12733, N12732, N12731, N12730, N12729, N12728, N12727, N12726, N12725, N12724, N12723, N12722, N12721, N12720, N12719, N12718, N12717, N12716, N12715, N12714, N12713, N12712, N12711, N12710, N12709, N12708, N12707, N12706, N12705, N12704, N12703, N12702, N12701, N12700, N12699, N12698, N12697, N12696, N12695, N12694, N12693, N12692, N12691, N12690, N12689, N12688, N12687, N12686, N12685, N12684, N12683, N12682, N12681, N12680, N12679, N12678, N12677, N12676, N12675 } = (N169)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12155)? { N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057 } : 1'b0;
  assign { N12802, N12801, N12800, N12799, N12798, N12797, N12796, N12795, N12794, N12793, N12792, N12791, N12790, N12789, N12788, N12787, N12786, N12785, N12784, N12783, N12782, N12781, N12780, N12779, N12778, N12777, N12776, N12775, N12774, N12773, N12772, N12771, N12770, N12769, N12768, N12767, N12766, N12765, N12764, N12763, N12762, N12761, N12760, N12759, N12758, N12757, N12756, N12755, N12754, N12753, N12752, N12751, N12750, N12749, N12748, N12747, N12746, N12745, N12744, N12743, N12742, N12741, N12740, N12739 } = (N170)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12220)? { N10378, N10377, N10376, N10375, N10374, N10373, N10372, N10371, N10370, N10369, N10368, N10367, N10366, N10365, N10364, N10363, N10362, N10361, N10360, N10359, N10358, N10357, N10356, N10355, N10354, N10353, N10352, N10351, N10350, N10349, N10348, N10347, N10346, N10345, N10344, N10343, N10342, N10341, N10340, N10339, N10338, N10337, N10336, N10335, N10334, N10333, N10332, N10331, N10330, N10329, N10328, N10327, N10326, N10325, N10324, N10323, N10322, N10321, N10320, N10319, N10318, N10317, N10316, N10315 } : 1'b0;
  assign { N12866, N12865, N12864, N12863, N12862, N12861, N12860, N12859, N12858, N12857, N12856, N12855, N12854, N12853, N12852, N12851, N12850, N12849, N12848, N12847, N12846, N12845, N12844, N12843, N12842, N12841, N12840, N12839, N12838, N12837, N12836, N12835, N12834, N12833, N12832, N12831, N12830, N12829, N12828, N12827, N12826, N12825, N12824, N12823, N12822, N12821, N12820, N12819, N12818, N12817, N12816, N12815, N12814, N12813, N12812, N12811, N12810, N12809, N12808, N12807, N12806, N12805, N12804, N12803 } = (N171)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12285)? { N10636, N10635, N10634, N10633, N10632, N10631, N10630, N10629, N10628, N10627, N10626, N10625, N10624, N10623, N10622, N10621, N10620, N10619, N10618, N10617, N10616, N10615, N10614, N10613, N10612, N10611, N10610, N10609, N10608, N10607, N10606, N10605, N10604, N10603, N10602, N10601, N10600, N10599, N10598, N10597, N10596, N10595, N10594, N10593, N10592, N10591, N10590, N10589, N10588, N10587, N10586, N10585, N10584, N10583, N10582, N10581, N10580, N10579, N10578, N10577, N10576, N10575, N10574, N10573 } : 1'b0;
  assign { N12930, N12929, N12928, N12927, N12926, N12925, N12924, N12923, N12922, N12921, N12920, N12919, N12918, N12917, N12916, N12915, N12914, N12913, N12912, N12911, N12910, N12909, N12908, N12907, N12906, N12905, N12904, N12903, N12902, N12901, N12900, N12899, N12898, N12897, N12896, N12895, N12894, N12893, N12892, N12891, N12890, N12889, N12888, N12887, N12886, N12885, N12884, N12883, N12882, N12881, N12880, N12879, N12878, N12877, N12876, N12875, N12874, N12873, N12872, N12871, N12870, N12869, N12868, N12867 } = (N172)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12350)? { N10894, N10893, N10892, N10891, N10890, N10889, N10888, N10887, N10886, N10885, N10884, N10883, N10882, N10881, N10880, N10879, N10878, N10877, N10876, N10875, N10874, N10873, N10872, N10871, N10870, N10869, N10868, N10867, N10866, N10865, N10864, N10863, N10862, N10861, N10860, N10859, N10858, N10857, N10856, N10855, N10854, N10853, N10852, N10851, N10850, N10849, N10848, N10847, N10846, N10845, N10844, N10843, N10842, N10841, N10840, N10839, N10838, N10837, N10836, N10835, N10834, N10833, N10832, N10831 } : 1'b0;
  assign { N12994, N12993, N12992, N12991, N12990, N12989, N12988, N12987, N12986, N12985, N12984, N12983, N12982, N12981, N12980, N12979, N12978, N12977, N12976, N12975, N12974, N12973, N12972, N12971, N12970, N12969, N12968, N12967, N12966, N12965, N12964, N12963, N12962, N12961, N12960, N12959, N12958, N12957, N12956, N12955, N12954, N12953, N12952, N12951, N12950, N12949, N12948, N12947, N12946, N12945, N12944, N12943, N12942, N12941, N12940, N12939, N12938, N12937, N12936, N12935, N12934, N12933, N12932, N12931 } = (N173)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12415)? { N11152, N11151, N11150, N11149, N11148, N11147, N11146, N11145, N11144, N11143, N11142, N11141, N11140, N11139, N11138, N11137, N11136, N11135, N11134, N11133, N11132, N11131, N11130, N11129, N11128, N11127, N11126, N11125, N11124, N11123, N11122, N11121, N11120, N11119, N11118, N11117, N11116, N11115, N11114, N11113, N11112, N11111, N11110, N11109, N11108, N11107, N11106, N11105, N11104, N11103, N11102, N11101, N11100, N11099, N11098, N11097, N11096, N11095, N11094, N11093, N11092, N11091, N11090, N11089 } : 1'b0;
  assign { N13058, N13057, N13056, N13055, N13054, N13053, N13052, N13051, N13050, N13049, N13048, N13047, N13046, N13045, N13044, N13043, N13042, N13041, N13040, N13039, N13038, N13037, N13036, N13035, N13034, N13033, N13032, N13031, N13030, N13029, N13028, N13027, N13026, N13025, N13024, N13023, N13022, N13021, N13020, N13019, N13018, N13017, N13016, N13015, N13014, N13013, N13012, N13011, N13010, N13009, N13008, N13007, N13006, N13005, N13004, N13003, N13002, N13001, N13000, N12999, N12998, N12997, N12996, N12995 } = (N174)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12480)? { N11410, N11409, N11408, N11407, N11406, N11405, N11404, N11403, N11402, N11401, N11400, N11399, N11398, N11397, N11396, N11395, N11394, N11393, N11392, N11391, N11390, N11389, N11388, N11387, N11386, N11385, N11384, N11383, N11382, N11381, N11380, N11379, N11378, N11377, N11376, N11375, N11374, N11373, N11372, N11371, N11370, N11369, N11368, N11367, N11366, N11365, N11364, N11363, N11362, N11361, N11360, N11359, N11358, N11357, N11356, N11355, N11354, N11353, N11352, N11351, N11350, N11349, N11348, N11347 } : 1'b0;
  assign { N13122, N13121, N13120, N13119, N13118, N13117, N13116, N13115, N13114, N13113, N13112, N13111, N13110, N13109, N13108, N13107, N13106, N13105, N13104, N13103, N13102, N13101, N13100, N13099, N13098, N13097, N13096, N13095, N13094, N13093, N13092, N13091, N13090, N13089, N13088, N13087, N13086, N13085, N13084, N13083, N13082, N13081, N13080, N13079, N13078, N13077, N13076, N13075, N13074, N13073, N13072, N13071, N13070, N13069, N13068, N13067, N13066, N13065, N13064, N13063, N13062, N13061, N13060, N13059 } = (N175)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12545)? { N11668, N11667, N11666, N11665, N11664, N11663, N11662, N11661, N11660, N11659, N11658, N11657, N11656, N11655, N11654, N11653, N11652, N11651, N11650, N11649, N11648, N11647, N11646, N11645, N11644, N11643, N11642, N11641, N11640, N11639, N11638, N11637, N11636, N11635, N11634, N11633, N11632, N11631, N11630, N11629, N11628, N11627, N11626, N11625, N11624, N11623, N11622, N11621, N11620, N11619, N11618, N11617, N11616, N11615, N11614, N11613, N11612, N11611, N11610, N11609, N11608, N11607, N11606, N11605 } : 1'b0;
  assign { N13186, N13185, N13184, N13183, N13182, N13181, N13180, N13179, N13178, N13177, N13176, N13175, N13174, N13173, N13172, N13171, N13170, N13169, N13168, N13167, N13166, N13165, N13164, N13163, N13162, N13161, N13160, N13159, N13158, N13157, N13156, N13155, N13154, N13153, N13152, N13151, N13150, N13149, N13148, N13147, N13146, N13145, N13144, N13143, N13142, N13141, N13140, N13139, N13138, N13137, N13136, N13135, N13134, N13133, N13132, N13131, N13130, N13129, N13128, N13127, N13126, N13125, N13124, N13123 } = (N176)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12610)? { N11926, N11925, N11924, N11923, N11922, N11921, N11920, N11919, N11918, N11917, N11916, N11915, N11914, N11913, N11912, N11911, N11910, N11909, N11908, N11907, N11906, N11905, N11904, N11903, N11902, N11901, N11900, N11899, N11898, N11897, N11896, N11895, N11894, N11893, N11892, N11891, N11890, N11889, N11888, N11887, N11886, N11885, N11884, N11883, N11882, N11881, N11880, N11879, N11878, N11877, N11876, N11875, N11874, N11873, N11872, N11871, N11870, N11869, N11868, N11867, N11866, N11865, N11864, N11863 } : 1'b0;
  assign { N13320, N13319, N13318, N13317, N13316, N13315, N13314, N13313, N13312, N13311, N13310, N13309, N13308, N13307, N13306, N13305, N13304, N13303, N13302, N13301, N13300, N13299, N13298, N13297, N13296, N13295, N13294, N13293, N13292, N13291, N13290, N13289, N13288, N13287, N13286, N13285, N13284, N13283, N13282, N13281, N13280, N13279, N13278, N13277, N13276, N13275, N13274, N13273, N13272, N13271, N13270, N13269, N13268, N13267, N13266, N13265, N13264, N13263, N13262, N13261, N13260, N13259, N13258, N13257, N13256, N13255, N13254, N13253, N13252, N13251, N13250, N13249, N13248, N13247, N13246, N13245, N13244, N13243, N13242, N13241, N13240, N13239, N13238, N13237, N13236, N13235, N13234, N13233, N13232, N13231, N13230, N13229, N13228, N13227, N13226, N13225, N13224, N13223, N13222, N13221, N13220, N13219, N13218, N13217, N13216, N13215, N13214, N13213, N13212, N13211, N13210, N13209, N13208, N13207, N13206, N13205, N13204, N13203, N13202, N13201, N13200, N13199, N13198, N13197, N13196, N13195, N13194, N13193, N13192 } = (N169)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12155)? { N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121 } : 1'b0;
  assign { N13449, N13448, N13447, N13446, N13445, N13444, N13443, N13442, N13441, N13440, N13439, N13438, N13437, N13436, N13435, N13434, N13433, N13432, N13431, N13430, N13429, N13428, N13427, N13426, N13425, N13424, N13423, N13422, N13421, N13420, N13419, N13418, N13417, N13416, N13415, N13414, N13413, N13412, N13411, N13410, N13409, N13408, N13407, N13406, N13405, N13404, N13403, N13402, N13401, N13400, N13399, N13398, N13397, N13396, N13395, N13394, N13393, N13392, N13391, N13390, N13389, N13388, N13387, N13386, N13385, N13384, N13383, N13382, N13381, N13380, N13379, N13378, N13377, N13376, N13375, N13374, N13373, N13372, N13371, N13370, N13369, N13368, N13367, N13366, N13365, N13364, N13363, N13362, N13361, N13360, N13359, N13358, N13357, N13356, N13355, N13354, N13353, N13352, N13351, N13350, N13349, N13348, N13347, N13346, N13345, N13344, N13343, N13342, N13341, N13340, N13339, N13338, N13337, N13336, N13335, N13334, N13333, N13332, N13331, N13330, N13329, N13328, N13327, N13326, N13325, N13324, N13323, N13322, N13321 } = (N170)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12220)? { N10507, N10506, N10505, N10504, N10503, N10502, N10501, N10500, N10499, N10498, N10497, N10496, N10495, N10494, N10493, N10492, N10491, N10490, N10489, N10488, N10487, N10486, N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422, N10421, N10420, N10419, N10418, N10417, N10416, N10415, N10414, N10413, N10412, N10411, N10410, N10409, N10408, N10407, N10406, N10405, N10404, N10403, N10402, N10401, N10400, N10399, N10398, N10397, N10396, N10395, N10394, N10393, N10392, N10391, N10390, N10389, N10388, N10387, N10386, N10385, N10384, N10383, N10382, N10381, N10380, N10379 } : 1'b0;
  assign { N13578, N13577, N13576, N13575, N13574, N13573, N13572, N13571, N13570, N13569, N13568, N13567, N13566, N13565, N13564, N13563, N13562, N13561, N13560, N13559, N13558, N13557, N13556, N13555, N13554, N13553, N13552, N13551, N13550, N13549, N13548, N13547, N13546, N13545, N13544, N13543, N13542, N13541, N13540, N13539, N13538, N13537, N13536, N13535, N13534, N13533, N13532, N13531, N13530, N13529, N13528, N13527, N13526, N13525, N13524, N13523, N13522, N13521, N13520, N13519, N13518, N13517, N13516, N13515, N13514, N13513, N13512, N13511, N13510, N13509, N13508, N13507, N13506, N13505, N13504, N13503, N13502, N13501, N13500, N13499, N13498, N13497, N13496, N13495, N13494, N13493, N13492, N13491, N13490, N13489, N13488, N13487, N13486, N13485, N13484, N13483, N13482, N13481, N13480, N13479, N13478, N13477, N13476, N13475, N13474, N13473, N13472, N13471, N13470, N13469, N13468, N13467, N13466, N13465, N13464, N13463, N13462, N13461, N13460, N13459, N13458, N13457, N13456, N13455, N13454, N13453, N13452, N13451, N13450 } = (N171)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12285)? { N10765, N10764, N10763, N10762, N10761, N10760, N10759, N10758, N10757, N10756, N10755, N10754, N10753, N10752, N10751, N10750, N10749, N10748, N10747, N10746, N10745, N10744, N10743, N10742, N10741, N10740, N10739, N10738, N10737, N10736, N10735, N10734, N10733, N10732, N10731, N10730, N10729, N10728, N10727, N10726, N10725, N10724, N10723, N10722, N10721, N10720, N10719, N10718, N10717, N10716, N10715, N10714, N10713, N10712, N10711, N10710, N10709, N10708, N10707, N10706, N10705, N10704, N10703, N10702, N10701, N10700, N10699, N10698, N10697, N10696, N10695, N10694, N10693, N10692, N10691, N10690, N10689, N10688, N10687, N10686, N10685, N10684, N10683, N10682, N10681, N10680, N10679, N10678, N10677, N10676, N10675, N10674, N10673, N10672, N10671, N10670, N10669, N10668, N10667, N10666, N10665, N10664, N10663, N10662, N10661, N10660, N10659, N10658, N10657, N10656, N10655, N10654, N10653, N10652, N10651, N10650, N10649, N10648, N10647, N10646, N10645, N10644, N10643, N10642, N10641, N10640, N10639, N10638, N10637 } : 1'b0;
  assign { N13707, N13706, N13705, N13704, N13703, N13702, N13701, N13700, N13699, N13698, N13697, N13696, N13695, N13694, N13693, N13692, N13691, N13690, N13689, N13688, N13687, N13686, N13685, N13684, N13683, N13682, N13681, N13680, N13679, N13678, N13677, N13676, N13675, N13674, N13673, N13672, N13671, N13670, N13669, N13668, N13667, N13666, N13665, N13664, N13663, N13662, N13661, N13660, N13659, N13658, N13657, N13656, N13655, N13654, N13653, N13652, N13651, N13650, N13649, N13648, N13647, N13646, N13645, N13644, N13643, N13642, N13641, N13640, N13639, N13638, N13637, N13636, N13635, N13634, N13633, N13632, N13631, N13630, N13629, N13628, N13627, N13626, N13625, N13624, N13623, N13622, N13621, N13620, N13619, N13618, N13617, N13616, N13615, N13614, N13613, N13612, N13611, N13610, N13609, N13608, N13607, N13606, N13605, N13604, N13603, N13602, N13601, N13600, N13599, N13598, N13597, N13596, N13595, N13594, N13593, N13592, N13591, N13590, N13589, N13588, N13587, N13586, N13585, N13584, N13583, N13582, N13581, N13580, N13579 } = (N172)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12350)? { N11023, N11022, N11021, N11020, N11019, N11018, N11017, N11016, N11015, N11014, N11013, N11012, N11011, N11010, N11009, N11008, N11007, N11006, N11005, N11004, N11003, N11002, N11001, N11000, N10999, N10998, N10997, N10996, N10995, N10994, N10993, N10992, N10991, N10990, N10989, N10988, N10987, N10986, N10985, N10984, N10983, N10982, N10981, N10980, N10979, N10978, N10977, N10976, N10975, N10974, N10973, N10972, N10971, N10970, N10969, N10968, N10967, N10966, N10965, N10964, N10963, N10962, N10961, N10960, N10959, N10958, N10957, N10956, N10955, N10954, N10953, N10952, N10951, N10950, N10949, N10948, N10947, N10946, N10945, N10944, N10943, N10942, N10941, N10940, N10939, N10938, N10937, N10936, N10935, N10934, N10933, N10932, N10931, N10930, N10929, N10928, N10927, N10926, N10925, N10924, N10923, N10922, N10921, N10920, N10919, N10918, N10917, N10916, N10915, N10914, N10913, N10912, N10911, N10910, N10909, N10908, N10907, N10906, N10905, N10904, N10903, N10902, N10901, N10900, N10899, N10898, N10897, N10896, N10895 } : 1'b0;
  assign { N13836, N13835, N13834, N13833, N13832, N13831, N13830, N13829, N13828, N13827, N13826, N13825, N13824, N13823, N13822, N13821, N13820, N13819, N13818, N13817, N13816, N13815, N13814, N13813, N13812, N13811, N13810, N13809, N13808, N13807, N13806, N13805, N13804, N13803, N13802, N13801, N13800, N13799, N13798, N13797, N13796, N13795, N13794, N13793, N13792, N13791, N13790, N13789, N13788, N13787, N13786, N13785, N13784, N13783, N13782, N13781, N13780, N13779, N13778, N13777, N13776, N13775, N13774, N13773, N13772, N13771, N13770, N13769, N13768, N13767, N13766, N13765, N13764, N13763, N13762, N13761, N13760, N13759, N13758, N13757, N13756, N13755, N13754, N13753, N13752, N13751, N13750, N13749, N13748, N13747, N13746, N13745, N13744, N13743, N13742, N13741, N13740, N13739, N13738, N13737, N13736, N13735, N13734, N13733, N13732, N13731, N13730, N13729, N13728, N13727, N13726, N13725, N13724, N13723, N13722, N13721, N13720, N13719, N13718, N13717, N13716, N13715, N13714, N13713, N13712, N13711, N13710, N13709, N13708 } = (N173)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12415)? { N11281, N11280, N11279, N11278, N11277, N11276, N11275, N11274, N11273, N11272, N11271, N11270, N11269, N11268, N11267, N11266, N11265, N11264, N11263, N11262, N11261, N11260, N11259, N11258, N11257, N11256, N11255, N11254, N11253, N11252, N11251, N11250, N11249, N11248, N11247, N11246, N11245, N11244, N11243, N11242, N11241, N11240, N11239, N11238, N11237, N11236, N11235, N11234, N11233, N11232, N11231, N11230, N11229, N11228, N11227, N11226, N11225, N11224, N11223, N11222, N11221, N11220, N11219, N11218, N11217, N11216, N11215, N11214, N11213, N11212, N11211, N11210, N11209, N11208, N11207, N11206, N11205, N11204, N11203, N11202, N11201, N11200, N11199, N11198, N11197, N11196, N11195, N11194, N11193, N11192, N11191, N11190, N11189, N11188, N11187, N11186, N11185, N11184, N11183, N11182, N11181, N11180, N11179, N11178, N11177, N11176, N11175, N11174, N11173, N11172, N11171, N11170, N11169, N11168, N11167, N11166, N11165, N11164, N11163, N11162, N11161, N11160, N11159, N11158, N11157, N11156, N11155, N11154, N11153 } : 1'b0;
  assign { N13965, N13964, N13963, N13962, N13961, N13960, N13959, N13958, N13957, N13956, N13955, N13954, N13953, N13952, N13951, N13950, N13949, N13948, N13947, N13946, N13945, N13944, N13943, N13942, N13941, N13940, N13939, N13938, N13937, N13936, N13935, N13934, N13933, N13932, N13931, N13930, N13929, N13928, N13927, N13926, N13925, N13924, N13923, N13922, N13921, N13920, N13919, N13918, N13917, N13916, N13915, N13914, N13913, N13912, N13911, N13910, N13909, N13908, N13907, N13906, N13905, N13904, N13903, N13902, N13901, N13900, N13899, N13898, N13897, N13896, N13895, N13894, N13893, N13892, N13891, N13890, N13889, N13888, N13887, N13886, N13885, N13884, N13883, N13882, N13881, N13880, N13879, N13878, N13877, N13876, N13875, N13874, N13873, N13872, N13871, N13870, N13869, N13868, N13867, N13866, N13865, N13864, N13863, N13862, N13861, N13860, N13859, N13858, N13857, N13856, N13855, N13854, N13853, N13852, N13851, N13850, N13849, N13848, N13847, N13846, N13845, N13844, N13843, N13842, N13841, N13840, N13839, N13838, N13837 } = (N174)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12480)? { N11539, N11538, N11537, N11536, N11535, N11534, N11533, N11532, N11531, N11530, N11529, N11528, N11527, N11526, N11525, N11524, N11523, N11522, N11521, N11520, N11519, N11518, N11517, N11516, N11515, N11514, N11513, N11512, N11511, N11510, N11509, N11508, N11507, N11506, N11505, N11504, N11503, N11502, N11501, N11500, N11499, N11498, N11497, N11496, N11495, N11494, N11493, N11492, N11491, N11490, N11489, N11488, N11487, N11486, N11485, N11484, N11483, N11482, N11481, N11480, N11479, N11478, N11477, N11476, N11475, N11474, N11473, N11472, N11471, N11470, N11469, N11468, N11467, N11466, N11465, N11464, N11463, N11462, N11461, N11460, N11459, N11458, N11457, N11456, N11455, N11454, N11453, N11452, N11451, N11450, N11449, N11448, N11447, N11446, N11445, N11444, N11443, N11442, N11441, N11440, N11439, N11438, N11437, N11436, N11435, N11434, N11433, N11432, N11431, N11430, N11429, N11428, N11427, N11426, N11425, N11424, N11423, N11422, N11421, N11420, N11419, N11418, N11417, N11416, N11415, N11414, N11413, N11412, N11411 } : 1'b0;
  assign { N14094, N14093, N14092, N14091, N14090, N14089, N14088, N14087, N14086, N14085, N14084, N14083, N14082, N14081, N14080, N14079, N14078, N14077, N14076, N14075, N14074, N14073, N14072, N14071, N14070, N14069, N14068, N14067, N14066, N14065, N14064, N14063, N14062, N14061, N14060, N14059, N14058, N14057, N14056, N14055, N14054, N14053, N14052, N14051, N14050, N14049, N14048, N14047, N14046, N14045, N14044, N14043, N14042, N14041, N14040, N14039, N14038, N14037, N14036, N14035, N14034, N14033, N14032, N14031, N14030, N14029, N14028, N14027, N14026, N14025, N14024, N14023, N14022, N14021, N14020, N14019, N14018, N14017, N14016, N14015, N14014, N14013, N14012, N14011, N14010, N14009, N14008, N14007, N14006, N14005, N14004, N14003, N14002, N14001, N14000, N13999, N13998, N13997, N13996, N13995, N13994, N13993, N13992, N13991, N13990, N13989, N13988, N13987, N13986, N13985, N13984, N13983, N13982, N13981, N13980, N13979, N13978, N13977, N13976, N13975, N13974, N13973, N13972, N13971, N13970, N13969, N13968, N13967, N13966 } = (N175)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12545)? { N11797, N11796, N11795, N11794, N11793, N11792, N11791, N11790, N11789, N11788, N11787, N11786, N11785, N11784, N11783, N11782, N11781, N11780, N11779, N11778, N11777, N11776, N11775, N11774, N11773, N11772, N11771, N11770, N11769, N11768, N11767, N11766, N11765, N11764, N11763, N11762, N11761, N11760, N11759, N11758, N11757, N11756, N11755, N11754, N11753, N11752, N11751, N11750, N11749, N11748, N11747, N11746, N11745, N11744, N11743, N11742, N11741, N11740, N11739, N11738, N11737, N11736, N11735, N11734, N11733, N11732, N11731, N11730, N11729, N11728, N11727, N11726, N11725, N11724, N11723, N11722, N11721, N11720, N11719, N11718, N11717, N11716, N11715, N11714, N11713, N11712, N11711, N11710, N11709, N11708, N11707, N11706, N11705, N11704, N11703, N11702, N11701, N11700, N11699, N11698, N11697, N11696, N11695, N11694, N11693, N11692, N11691, N11690, N11689, N11688, N11687, N11686, N11685, N11684, N11683, N11682, N11681, N11680, N11679, N11678, N11677, N11676, N11675, N11674, N11673, N11672, N11671, N11670, N11669 } : 1'b0;
  assign { N14223, N14222, N14221, N14220, N14219, N14218, N14217, N14216, N14215, N14214, N14213, N14212, N14211, N14210, N14209, N14208, N14207, N14206, N14205, N14204, N14203, N14202, N14201, N14200, N14199, N14198, N14197, N14196, N14195, N14194, N14193, N14192, N14191, N14190, N14189, N14188, N14187, N14186, N14185, N14184, N14183, N14182, N14181, N14180, N14179, N14178, N14177, N14176, N14175, N14174, N14173, N14172, N14171, N14170, N14169, N14168, N14167, N14166, N14165, N14164, N14163, N14162, N14161, N14160, N14159, N14158, N14157, N14156, N14155, N14154, N14153, N14152, N14151, N14150, N14149, N14148, N14147, N14146, N14145, N14144, N14143, N14142, N14141, N14140, N14139, N14138, N14137, N14136, N14135, N14134, N14133, N14132, N14131, N14130, N14129, N14128, N14127, N14126, N14125, N14124, N14123, N14122, N14121, N14120, N14119, N14118, N14117, N14116, N14115, N14114, N14113, N14112, N14111, N14110, N14109, N14108, N14107, N14106, N14105, N14104, N14103, N14102, N14101, N14100, N14099, N14098, N14097, N14096, N14095 } = (N176)? ex_i[257:129] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N12610)? { N12055, N12054, N12053, N12052, N12051, N12050, N12049, N12048, N12047, N12046, N12045, N12044, N12043, N12042, N12041, N12040, N12039, N12038, N12037, N12036, N12035, N12034, N12033, N12032, N12031, N12030, N12029, N12028, N12027, N12026, N12025, N12024, N12023, N12022, N12021, N12020, N12019, N12018, N12017, N12016, N12015, N12014, N12013, N12012, N12011, N12010, N12009, N12008, N12007, N12006, N12005, N12004, N12003, N12002, N12001, N12000, N11999, N11998, N11997, N11996, N11995, N11994, N11993, N11992, N11991, N11990, N11989, N11988, N11987, N11986, N11985, N11984, N11983, N11982, N11981, N11980, N11979, N11978, N11977, N11976, N11975, N11974, N11973, N11972, N11971, N11970, N11969, N11968, N11967, N11966, N11965, N11964, N11963, N11962, N11961, N11960, N11959, N11958, N11957, N11956, N11955, N11954, N11953, N11952, N11951, N11950, N11949, N11948, N11947, N11946, N11945, N11944, N11943, N11942, N11941, N11940, N11939, N11938, N11937, N11936, N11935, N11934, N11933, N11932, N11931, N11930, N11929, N11928, N11927 } : 1'b0;
  assign { N14299, N14298, N14297, N14296, N14295, N14294, N14293, N14292, N14291, N14290, N14289, N14288, N14287, N14286, N14285, N14284, N14283, N14282, N14281, N14280, N14279, N14278, N14277, N14276, N14275, N14274, N14273, N14272, N14271, N14270, N14269, N14268, N14267, N14266, N14265, N14264, N14263, N14262, N14261, N14260, N14259, N14258, N14257, N14256, N14255, N14254, N14253, N14252, N14251, N14250, N14249, N14248, N14247, N14246, N14245, N14244, N14243, N14242, N14241, N14240, N14239, N14238, N14237, N14236 } = (N169)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12155)? { N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186 } : 1'b0;
  assign { N14363, N14362, N14361, N14360, N14359, N14358, N14357, N14356, N14355, N14354, N14353, N14352, N14351, N14350, N14349, N14348, N14347, N14346, N14345, N14344, N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336, N14335, N14334, N14333, N14332, N14331, N14330, N14329, N14328, N14327, N14326, N14325, N14324, N14323, N14322, N14321, N14320, N14319, N14318, N14317, N14316, N14315, N14314, N14313, N14312, N14311, N14310, N14309, N14308, N14307, N14306, N14305, N14304, N14303, N14302, N14301, N14300 } = (N170)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12220)? { N10507, N10506, N10505, N10504, N10503, N10502, N10501, N10500, N10499, N10498, N10497, N10496, N10495, N10494, N10493, N10492, N10491, N10490, N10489, N10488, N10487, N10486, N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444 } : 1'b0;
  assign { N14427, N14426, N14425, N14424, N14423, N14422, N14421, N14420, N14419, N14418, N14417, N14416, N14415, N14414, N14413, N14412, N14411, N14410, N14409, N14408, N14407, N14406, N14405, N14404, N14403, N14402, N14401, N14400, N14399, N14398, N14397, N14396, N14395, N14394, N14393, N14392, N14391, N14390, N14389, N14388, N14387, N14386, N14385, N14384, N14383, N14382, N14381, N14380, N14379, N14378, N14377, N14376, N14375, N14374, N14373, N14372, N14371, N14370, N14369, N14368, N14367, N14366, N14365, N14364 } = (N171)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12285)? { N10765, N10764, N10763, N10762, N10761, N10760, N10759, N10758, N10757, N10756, N10755, N10754, N10753, N10752, N10751, N10750, N10749, N10748, N10747, N10746, N10745, N10744, N10743, N10742, N10741, N10740, N10739, N10738, N10737, N10736, N10735, N10734, N10733, N10732, N10731, N10730, N10729, N10728, N10727, N10726, N10725, N10724, N10723, N10722, N10721, N10720, N10719, N10718, N10717, N10716, N10715, N10714, N10713, N10712, N10711, N10710, N10709, N10708, N10707, N10706, N10705, N10704, N10703, N10702 } : 1'b0;
  assign { N14491, N14490, N14489, N14488, N14487, N14486, N14485, N14484, N14483, N14482, N14481, N14480, N14479, N14478, N14477, N14476, N14475, N14474, N14473, N14472, N14471, N14470, N14469, N14468, N14467, N14466, N14465, N14464, N14463, N14462, N14461, N14460, N14459, N14458, N14457, N14456, N14455, N14454, N14453, N14452, N14451, N14450, N14449, N14448, N14447, N14446, N14445, N14444, N14443, N14442, N14441, N14440, N14439, N14438, N14437, N14436, N14435, N14434, N14433, N14432, N14431, N14430, N14429, N14428 } = (N172)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12350)? { N11023, N11022, N11021, N11020, N11019, N11018, N11017, N11016, N11015, N11014, N11013, N11012, N11011, N11010, N11009, N11008, N11007, N11006, N11005, N11004, N11003, N11002, N11001, N11000, N10999, N10998, N10997, N10996, N10995, N10994, N10993, N10992, N10991, N10990, N10989, N10988, N10987, N10986, N10985, N10984, N10983, N10982, N10981, N10980, N10979, N10978, N10977, N10976, N10975, N10974, N10973, N10972, N10971, N10970, N10969, N10968, N10967, N10966, N10965, N10964, N10963, N10962, N10961, N10960 } : 1'b0;
  assign { N14555, N14554, N14553, N14552, N14551, N14550, N14549, N14548, N14547, N14546, N14545, N14544, N14543, N14542, N14541, N14540, N14539, N14538, N14537, N14536, N14535, N14534, N14533, N14532, N14531, N14530, N14529, N14528, N14527, N14526, N14525, N14524, N14523, N14522, N14521, N14520, N14519, N14518, N14517, N14516, N14515, N14514, N14513, N14512, N14511, N14510, N14509, N14508, N14507, N14506, N14505, N14504, N14503, N14502, N14501, N14500, N14499, N14498, N14497, N14496, N14495, N14494, N14493, N14492 } = (N173)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12415)? { N11281, N11280, N11279, N11278, N11277, N11276, N11275, N11274, N11273, N11272, N11271, N11270, N11269, N11268, N11267, N11266, N11265, N11264, N11263, N11262, N11261, N11260, N11259, N11258, N11257, N11256, N11255, N11254, N11253, N11252, N11251, N11250, N11249, N11248, N11247, N11246, N11245, N11244, N11243, N11242, N11241, N11240, N11239, N11238, N11237, N11236, N11235, N11234, N11233, N11232, N11231, N11230, N11229, N11228, N11227, N11226, N11225, N11224, N11223, N11222, N11221, N11220, N11219, N11218 } : 1'b0;
  assign { N14619, N14618, N14617, N14616, N14615, N14614, N14613, N14612, N14611, N14610, N14609, N14608, N14607, N14606, N14605, N14604, N14603, N14602, N14601, N14600, N14599, N14598, N14597, N14596, N14595, N14594, N14593, N14592, N14591, N14590, N14589, N14588, N14587, N14586, N14585, N14584, N14583, N14582, N14581, N14580, N14579, N14578, N14577, N14576, N14575, N14574, N14573, N14572, N14571, N14570, N14569, N14568, N14567, N14566, N14565, N14564, N14563, N14562, N14561, N14560, N14559, N14558, N14557, N14556 } = (N174)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12480)? { N11539, N11538, N11537, N11536, N11535, N11534, N11533, N11532, N11531, N11530, N11529, N11528, N11527, N11526, N11525, N11524, N11523, N11522, N11521, N11520, N11519, N11518, N11517, N11516, N11515, N11514, N11513, N11512, N11511, N11510, N11509, N11508, N11507, N11506, N11505, N11504, N11503, N11502, N11501, N11500, N11499, N11498, N11497, N11496, N11495, N11494, N11493, N11492, N11491, N11490, N11489, N11488, N11487, N11486, N11485, N11484, N11483, N11482, N11481, N11480, N11479, N11478, N11477, N11476 } : 1'b0;
  assign { N14683, N14682, N14681, N14680, N14679, N14678, N14677, N14676, N14675, N14674, N14673, N14672, N14671, N14670, N14669, N14668, N14667, N14666, N14665, N14664, N14663, N14662, N14661, N14660, N14659, N14658, N14657, N14656, N14655, N14654, N14653, N14652, N14651, N14650, N14649, N14648, N14647, N14646, N14645, N14644, N14643, N14642, N14641, N14640, N14639, N14638, N14637, N14636, N14635, N14634, N14633, N14632, N14631, N14630, N14629, N14628, N14627, N14626, N14625, N14624, N14623, N14622, N14621, N14620 } = (N175)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12545)? { N11797, N11796, N11795, N11794, N11793, N11792, N11791, N11790, N11789, N11788, N11787, N11786, N11785, N11784, N11783, N11782, N11781, N11780, N11779, N11778, N11777, N11776, N11775, N11774, N11773, N11772, N11771, N11770, N11769, N11768, N11767, N11766, N11765, N11764, N11763, N11762, N11761, N11760, N11759, N11758, N11757, N11756, N11755, N11754, N11753, N11752, N11751, N11750, N11749, N11748, N11747, N11746, N11745, N11744, N11743, N11742, N11741, N11740, N11739, N11738, N11737, N11736, N11735, N11734 } : 1'b0;
  assign { N14747, N14746, N14745, N14744, N14743, N14742, N14741, N14740, N14739, N14738, N14737, N14736, N14735, N14734, N14733, N14732, N14731, N14730, N14729, N14728, N14727, N14726, N14725, N14724, N14723, N14722, N14721, N14720, N14719, N14718, N14717, N14716, N14715, N14714, N14713, N14712, N14711, N14710, N14709, N14708, N14707, N14706, N14705, N14704, N14703, N14702, N14701, N14700, N14699, N14698, N14697, N14696, N14695, N14694, N14693, N14692, N14691, N14690, N14689, N14688, N14687, N14686, N14685, N14684 } = (N176)? ex_i[257:194] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12610)? { N12055, N12054, N12053, N12052, N12051, N12050, N12049, N12048, N12047, N12046, N12045, N12044, N12043, N12042, N12041, N12040, N12039, N12038, N12037, N12036, N12035, N12034, N12033, N12032, N12031, N12030, N12029, N12028, N12027, N12026, N12025, N12024, N12023, N12022, N12021, N12020, N12019, N12018, N12017, N12016, N12015, N12014, N12013, N12012, N12011, N12010, N12009, N12008, N12007, N12006, N12005, N12004, N12003, N12002, N12001, N12000, N11999, N11998, N11997, N11996, N11995, N11994, N11993, N11992 } : 1'b0;
  assign { N15259, N15258, N15257, N15256, N15255, N15254, N15253, N15252, N15251, N15250, N15249, N15248, N15247, N15246, N15245, N15244, N15243, N15242, N15241, N15240, N15239, N15238, N15237, N15236, N15235, N15234, N15233, N15232, N15231, N15230, N15229, N15228, N15227, N15226, N15225, N15224, N15223, N15222, N15221, N15220, N15219, N15218, N15217, N15216, N15215, N15214, N15213, N15212, N15211, N15210, N15209, N15208, N15207, N15206, N15205, N15204, N15203, N15202, N15201, N15200, N15199, N15198, N15197, N15196, N15195, N15194, N15193, N15192, N15191, N15190, N15189, N15188, N15187, N15186, N15185, N15184, N15183, N15182, N15181, N15180, N15179, N15178, N15177, N15176, N15175, N15174, N15173, N15172, N15171, N15170, N15169, N15168, N15167, N15166, N15165, N15164, N15163, N15162, N15161, N15160, N15159, N15158, N15157, N15156, N15155, N15154, N15153, N15152, N15151, N15150, N15149, N15148, N15147, N15146, N15145, N15144, N15143, N15142, N15141, N15140, N15139, N15138, N15137, N15136, N15135, N15134, N15133, N15132, N15131, N15130, N15129, N15128, N15127, N15126, N15125, N15124, N15123, N15122, N15121, N15120, N15119, N15118, N15117, N15116, N15115, N15114, N15113, N15112, N15111, N15110, N15109, N15108, N15107, N15106, N15105, N15104, N15103, N15102, N15101, N15100, N15099, N15098, N15097, N15096, N15095, N15094, N15093, N15092, N15091, N15090, N15089, N15088, N15087, N15086, N15085, N15084, N15083, N15082, N15081, N15080, N15079, N15078, N15077, N15076, N15075, N15074, N15073, N15072, N15071, N15070, N15069, N15068, N15067, N15066, N15065, N15064, N15063, N15062, N15061, N15060, N15059, N15058, N15057, N15056, N15055, N15054, N15053, N15052, N15051, N15050, N15049, N15048, N15047, N15046, N15045, N15044, N15043, N15042, N15041, N15040, N15039, N15038, N15037, N15036, N15035, N15034, N15033, N15032, N15031, N15030, N15029, N15028, N15027, N15026, N15025, N15024, N15023, N15022, N15021, N15020, N15019, N15018, N15017, N15016, N15015, N15014, N15013, N15012, N15011, N15010, N15009, N15008, N15007, N15006, N15005, N15004, N15003, N15002, N15001, N15000, N14999, N14998, N14997, N14996, N14995, N14994, N14993, N14992, N14991, N14990, N14989, N14988, N14987, N14986, N14985, N14984, N14983, N14982, N14981, N14980, N14979, N14978, N14977, N14976, N14975, N14974, N14973, N14972, N14971, N14970, N14969, N14968, N14967, N14966, N14965, N14964, N14963, N14962, N14961, N14960, N14959, N14958, N14957, N14956, N14955, N14954, N14953, N14952, N14951, N14950, N14949, N14948, N14947, N14946, N14945, N14944, N14943, N14942, N14941, N14940, N14939, N14938, N14937, N14936, N14935, N14934, N14933, N14932, N14931, N14930, N14929, N14928, N14927, N14926, N14925, N14924, N14923, N14922, N14921, N14920, N14919, N14918, N14917, N14916, N14915, N14914, N14913, N14912, N14911, N14910, N14909, N14908, N14907, N14906, N14905, N14904, N14903, N14902, N14901, N14900, N14899, N14898, N14897, N14896, N14895, N14894, N14893, N14892, N14891, N14890, N14889, N14888, N14887, N14886, N14885, N14884, N14883, N14882, N14881, N14880, N14879, N14878, N14877, N14876, N14875, N14874, N14873, N14872, N14871, N14870, N14869, N14868, N14867, N14866, N14865, N14864, N14863, N14862, N14861, N14860, N14859, N14858, N14857, N14856, N14855, N14854, N14853, N14852, N14851, N14850, N14849, N14848, N14847, N14846, N14845, N14844, N14843, N14842, N14841, N14840, N14839, N14838, N14837, N14836, N14835, N14834, N14833, N14832, N14831, N14830, N14829, N14828, N14827, N14826, N14825, N14824, N14823, N14822, N14821, N14820, N14819, N14818, N14817, N14816, N14815, N14814, N14813, N14812, N14811, N14810, N14809, N14808, N14807, N14806, N14805, N14804, N14803, N14802, N14801, N14800, N14799, N14798, N14797, N14796, N14795, N14794, N14793, N14792, N14791, N14790, N14789, N14788, N14787, N14786, N14785, N14784, N14783, N14782, N14781, N14780, N14779, N14778, N14777, N14776, N14775, N14774, N14773, N14772, N14771, N14770, N14769, N14768, N14767, N14766, N14765, N14764, N14763, N14762, N14761, N14760, N14759, N14758, N14757, N14756, N14755, N14754, N14753, N14752, N14751, N14750, N14749, N14748 } = (N177)? { N14747, N14746, N14745, N14744, N14743, N14742, N14741, N14740, N14739, N14738, N14737, N14736, N14735, N14734, N14733, N14732, N14731, N14730, N14729, N14728, N14727, N14726, N14725, N14724, N14723, N14722, N14721, N14720, N14719, N14718, N14717, N14716, N14715, N14714, N14713, N14712, N14711, N14710, N14709, N14708, N14707, N14706, N14705, N14704, N14703, N14702, N14701, N14700, N14699, N14698, N14697, N14696, N14695, N14694, N14693, N14692, N14691, N14690, N14689, N14688, N14687, N14686, N14685, N14684, N14683, N14682, N14681, N14680, N14679, N14678, N14677, N14676, N14675, N14674, N14673, N14672, N14671, N14670, N14669, N14668, N14667, N14666, N14665, N14664, N14663, N14662, N14661, N14660, N14659, N14658, N14657, N14656, N14655, N14654, N14653, N14652, N14651, N14650, N14649, N14648, N14647, N14646, N14645, N14644, N14643, N14642, N14641, N14640, N14639, N14638, N14637, N14636, N14635, N14634, N14633, N14632, N14631, N14630, N14629, N14628, N14627, N14626, N14625, N14624, N14623, N14622, N14621, N14620, N14619, N14618, N14617, N14616, N14615, N14614, N14613, N14612, N14611, N14610, N14609, N14608, N14607, N14606, N14605, N14604, N14603, N14602, N14601, N14600, N14599, N14598, N14597, N14596, N14595, N14594, N14593, N14592, N14591, N14590, N14589, N14588, N14587, N14586, N14585, N14584, N14583, N14582, N14581, N14580, N14579, N14578, N14577, N14576, N14575, N14574, N14573, N14572, N14571, N14570, N14569, N14568, N14567, N14566, N14565, N14564, N14563, N14562, N14561, N14560, N14559, N14558, N14557, N14556, N14555, N14554, N14553, N14552, N14551, N14550, N14549, N14548, N14547, N14546, N14545, N14544, N14543, N14542, N14541, N14540, N14539, N14538, N14537, N14536, N14535, N14534, N14533, N14532, N14531, N14530, N14529, N14528, N14527, N14526, N14525, N14524, N14523, N14522, N14521, N14520, N14519, N14518, N14517, N14516, N14515, N14514, N14513, N14512, N14511, N14510, N14509, N14508, N14507, N14506, N14505, N14504, N14503, N14502, N14501, N14500, N14499, N14498, N14497, N14496, N14495, N14494, N14493, N14492, N14491, N14490, N14489, N14488, N14487, N14486, N14485, N14484, N14483, N14482, N14481, N14480, N14479, N14478, N14477, N14476, N14475, N14474, N14473, N14472, N14471, N14470, N14469, N14468, N14467, N14466, N14465, N14464, N14463, N14462, N14461, N14460, N14459, N14458, N14457, N14456, N14455, N14454, N14453, N14452, N14451, N14450, N14449, N14448, N14447, N14446, N14445, N14444, N14443, N14442, N14441, N14440, N14439, N14438, N14437, N14436, N14435, N14434, N14433, N14432, N14431, N14430, N14429, N14428, N14427, N14426, N14425, N14424, N14423, N14422, N14421, N14420, N14419, N14418, N14417, N14416, N14415, N14414, N14413, N14412, N14411, N14410, N14409, N14408, N14407, N14406, N14405, N14404, N14403, N14402, N14401, N14400, N14399, N14398, N14397, N14396, N14395, N14394, N14393, N14392, N14391, N14390, N14389, N14388, N14387, N14386, N14385, N14384, N14383, N14382, N14381, N14380, N14379, N14378, N14377, N14376, N14375, N14374, N14373, N14372, N14371, N14370, N14369, N14368, N14367, N14366, N14365, N14364, N14363, N14362, N14361, N14360, N14359, N14358, N14357, N14356, N14355, N14354, N14353, N14352, N14351, N14350, N14349, N14348, N14347, N14346, N14345, N14344, N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336, N14335, N14334, N14333, N14332, N14331, N14330, N14329, N14328, N14327, N14326, N14325, N14324, N14323, N14322, N14321, N14320, N14319, N14318, N14317, N14316, N14315, N14314, N14313, N14312, N14311, N14310, N14309, N14308, N14307, N14306, N14305, N14304, N14303, N14302, N14301, N14300, N14299, N14298, N14297, N14296, N14295, N14294, N14293, N14292, N14291, N14290, N14289, N14288, N14287, N14286, N14285, N14284, N14283, N14282, N14281, N14280, N14279, N14278, N14277, N14276, N14275, N14274, N14273, N14272, N14271, N14270, N14269, N14268, N14267, N14266, N14265, N14264, N14263, N14262, N14261, N14260, N14259, N14258, N14257, N14256, N14255, N14254, N14253, N14252, N14251, N14250, N14249, N14248, N14247, N14246, N14245, N14244, N14243, N14242, N14241, N14240, N14239, N14238, N14237, N14236 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N178)? { N12055, N12054, N12053, N12052, N12051, N12050, N12049, N12048, N12047, N12046, N12045, N12044, N12043, N12042, N12041, N12040, N12039, N12038, N12037, N12036, N12035, N12034, N12033, N12032, N12031, N12030, N12029, N12028, N12027, N12026, N12025, N12024, N12023, N12022, N12021, N12020, N12019, N12018, N12017, N12016, N12015, N12014, N12013, N12012, N12011, N12010, N12009, N12008, N12007, N12006, N12005, N12004, N12003, N12002, N12001, N12000, N11999, N11998, N11997, N11996, N11995, N11994, N11993, N11992, N11797, N11796, N11795, N11794, N11793, N11792, N11791, N11790, N11789, N11788, N11787, N11786, N11785, N11784, N11783, N11782, N11781, N11780, N11779, N11778, N11777, N11776, N11775, N11774, N11773, N11772, N11771, N11770, N11769, N11768, N11767, N11766, N11765, N11764, N11763, N11762, N11761, N11760, N11759, N11758, N11757, N11756, N11755, N11754, N11753, N11752, N11751, N11750, N11749, N11748, N11747, N11746, N11745, N11744, N11743, N11742, N11741, N11740, N11739, N11738, N11737, N11736, N11735, N11734, N11539, N11538, N11537, N11536, N11535, N11534, N11533, N11532, N11531, N11530, N11529, N11528, N11527, N11526, N11525, N11524, N11523, N11522, N11521, N11520, N11519, N11518, N11517, N11516, N11515, N11514, N11513, N11512, N11511, N11510, N11509, N11508, N11507, N11506, N11505, N11504, N11503, N11502, N11501, N11500, N11499, N11498, N11497, N11496, N11495, N11494, N11493, N11492, N11491, N11490, N11489, N11488, N11487, N11486, N11485, N11484, N11483, N11482, N11481, N11480, N11479, N11478, N11477, N11476, N11281, N11280, N11279, N11278, N11277, N11276, N11275, N11274, N11273, N11272, N11271, N11270, N11269, N11268, N11267, N11266, N11265, N11264, N11263, N11262, N11261, N11260, N11259, N11258, N11257, N11256, N11255, N11254, N11253, N11252, N11251, N11250, N11249, N11248, N11247, N11246, N11245, N11244, N11243, N11242, N11241, N11240, N11239, N11238, N11237, N11236, N11235, N11234, N11233, N11232, N11231, N11230, N11229, N11228, N11227, N11226, N11225, N11224, N11223, N11222, N11221, N11220, N11219, N11218, N11023, N11022, N11021, N11020, N11019, N11018, N11017, N11016, N11015, N11014, N11013, N11012, N11011, N11010, N11009, N11008, N11007, N11006, N11005, N11004, N11003, N11002, N11001, N11000, N10999, N10998, N10997, N10996, N10995, N10994, N10993, N10992, N10991, N10990, N10989, N10988, N10987, N10986, N10985, N10984, N10983, N10982, N10981, N10980, N10979, N10978, N10977, N10976, N10975, N10974, N10973, N10972, N10971, N10970, N10969, N10968, N10967, N10966, N10965, N10964, N10963, N10962, N10961, N10960, N10765, N10764, N10763, N10762, N10761, N10760, N10759, N10758, N10757, N10756, N10755, N10754, N10753, N10752, N10751, N10750, N10749, N10748, N10747, N10746, N10745, N10744, N10743, N10742, N10741, N10740, N10739, N10738, N10737, N10736, N10735, N10734, N10733, N10732, N10731, N10730, N10729, N10728, N10727, N10726, N10725, N10724, N10723, N10722, N10721, N10720, N10719, N10718, N10717, N10716, N10715, N10714, N10713, N10712, N10711, N10710, N10709, N10708, N10707, N10706, N10705, N10704, N10703, N10702, N10507, N10506, N10505, N10504, N10503, N10502, N10501, N10500, N10499, N10498, N10497, N10496, N10495, N10494, N10493, N10492, N10491, N10490, N10489, N10488, N10487, N10486, N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186 } : 1'b0;
  assign N177 = N14234;
  assign N178 = N14235;
  assign { N16291, N16290, N16289, N16288, N16287, N16286, N16285, N16284, N16283, N16282, N16281, N16280, N16279, N16278, N16277, N16276, N16275, N16274, N16273, N16272, N16271, N16270, N16269, N16268, N16267, N16266, N16265, N16264, N16263, N16262, N16261, N16260, N16259, N16258, N16257, N16256, N16255, N16254, N16253, N16252, N16251, N16250, N16249, N16248, N16247, N16246, N16245, N16244, N16243, N16242, N16241, N16240, N16239, N16238, N16237, N16236, N16235, N16234, N16233, N16232, N16231, N16230, N16229, N16228, N16227, N16226, N16225, N16224, N16223, N16222, N16221, N16220, N16219, N16218, N16217, N16216, N16215, N16214, N16213, N16212, N16211, N16210, N16209, N16208, N16207, N16206, N16205, N16204, N16203, N16202, N16201, N16200, N16199, N16198, N16197, N16196, N16195, N16194, N16193, N16192, N16191, N16190, N16189, N16188, N16187, N16186, N16185, N16184, N16183, N16182, N16181, N16180, N16179, N16178, N16177, N16176, N16175, N16174, N16173, N16172, N16171, N16170, N16169, N16168, N16167, N16166, N16165, N16164, N16163, N16162, N16161, N16160, N16159, N16158, N16157, N16156, N16155, N16154, N16153, N16152, N16151, N16150, N16149, N16148, N16147, N16146, N16145, N16144, N16143, N16142, N16141, N16140, N16139, N16138, N16137, N16136, N16135, N16134, N16133, N16132, N16131, N16130, N16129, N16128, N16127, N16126, N16125, N16124, N16123, N16122, N16121, N16120, N16119, N16118, N16117, N16116, N16115, N16114, N16113, N16112, N16111, N16110, N16109, N16108, N16107, N16106, N16105, N16104, N16103, N16102, N16101, N16100, N16099, N16098, N16097, N16096, N16095, N16094, N16093, N16092, N16091, N16090, N16089, N16088, N16087, N16086, N16085, N16084, N16083, N16082, N16081, N16080, N16079, N16078, N16077, N16076, N16075, N16074, N16073, N16072, N16071, N16070, N16069, N16068, N16067, N16066, N16065, N16064, N16063, N16062, N16061, N16060, N16059, N16058, N16057, N16056, N16055, N16054, N16053, N16052, N16051, N16050, N16049, N16048, N16047, N16046, N16045, N16044, N16043, N16042, N16041, N16040, N16039, N16038, N16037, N16036, N16035, N16034, N16033, N16032, N16031, N16030, N16029, N16028, N16027, N16026, N16025, N16024, N16023, N16022, N16021, N16020, N16019, N16018, N16017, N16016, N16015, N16014, N16013, N16012, N16011, N16010, N16009, N16008, N16007, N16006, N16005, N16004, N16003, N16002, N16001, N16000, N15999, N15998, N15997, N15996, N15995, N15994, N15993, N15992, N15991, N15990, N15989, N15988, N15987, N15986, N15985, N15984, N15983, N15982, N15981, N15980, N15979, N15978, N15977, N15976, N15975, N15974, N15973, N15972, N15971, N15970, N15969, N15968, N15967, N15966, N15965, N15964, N15963, N15962, N15961, N15960, N15959, N15958, N15957, N15956, N15955, N15954, N15953, N15952, N15951, N15950, N15949, N15948, N15947, N15946, N15945, N15944, N15943, N15942, N15941, N15940, N15939, N15938, N15937, N15936, N15935, N15934, N15933, N15932, N15931, N15930, N15929, N15928, N15927, N15926, N15925, N15924, N15923, N15922, N15921, N15920, N15919, N15918, N15917, N15916, N15915, N15914, N15913, N15912, N15911, N15910, N15909, N15908, N15907, N15906, N15905, N15904, N15903, N15902, N15901, N15900, N15899, N15898, N15897, N15896, N15895, N15894, N15893, N15892, N15891, N15890, N15889, N15888, N15887, N15886, N15885, N15884, N15883, N15882, N15881, N15880, N15879, N15878, N15877, N15876, N15875, N15874, N15873, N15872, N15871, N15870, N15869, N15868, N15867, N15866, N15865, N15864, N15863, N15862, N15861, N15860, N15859, N15858, N15857, N15856, N15855, N15854, N15853, N15852, N15851, N15850, N15849, N15848, N15847, N15846, N15845, N15844, N15843, N15842, N15841, N15840, N15839, N15838, N15837, N15836, N15835, N15834, N15833, N15832, N15831, N15830, N15829, N15828, N15827, N15826, N15825, N15824, N15823, N15822, N15821, N15820, N15819, N15818, N15817, N15816, N15815, N15814, N15813, N15812, N15811, N15810, N15809, N15808, N15807, N15806, N15805, N15804, N15803, N15802, N15801, N15800, N15799, N15798, N15797, N15796, N15795, N15794, N15793, N15792, N15791, N15790, N15789, N15788, N15787, N15786, N15785, N15784, N15783, N15782, N15781, N15780, N15779, N15778, N15777, N15776, N15775, N15774, N15773, N15772, N15771, N15770, N15769, N15768, N15767, N15766, N15765, N15764, N15763, N15762, N15761, N15760, N15759, N15758, N15757, N15756, N15755, N15754, N15753, N15752, N15751, N15750, N15749, N15748, N15747, N15746, N15745, N15744, N15743, N15742, N15741, N15740, N15739, N15738, N15737, N15736, N15735, N15734, N15733, N15732, N15731, N15730, N15729, N15728, N15727, N15726, N15725, N15724, N15723, N15722, N15721, N15720, N15719, N15718, N15717, N15716, N15715, N15714, N15713, N15712, N15711, N15710, N15709, N15708, N15707, N15706, N15705, N15704, N15703, N15702, N15701, N15700, N15699, N15698, N15697, N15696, N15695, N15694, N15693, N15692, N15691, N15690, N15689, N15688, N15687, N15686, N15685, N15684, N15683, N15682, N15681, N15680, N15679, N15678, N15677, N15676, N15675, N15674, N15673, N15672, N15671, N15670, N15669, N15668, N15667, N15666, N15665, N15664, N15663, N15662, N15661, N15660, N15659, N15658, N15657, N15656, N15655, N15654, N15653, N15652, N15651, N15650, N15649, N15648, N15647, N15646, N15645, N15644, N15643, N15642, N15641, N15640, N15639, N15638, N15637, N15636, N15635, N15634, N15633, N15632, N15631, N15630, N15629, N15628, N15627, N15626, N15625, N15624, N15623, N15622, N15621, N15620, N15619, N15618, N15617, N15616, N15615, N15614, N15613, N15612, N15611, N15610, N15609, N15608, N15607, N15606, N15605, N15604, N15603, N15602, N15601, N15600, N15599, N15598, N15597, N15596, N15595, N15594, N15593, N15592, N15591, N15590, N15589, N15588, N15587, N15586, N15585, N15584, N15583, N15582, N15581, N15580, N15579, N15578, N15577, N15576, N15575, N15574, N15573, N15572, N15571, N15570, N15569, N15568, N15567, N15566, N15565, N15564, N15563, N15562, N15561, N15560, N15559, N15558, N15557, N15556, N15555, N15554, N15553, N15552, N15551, N15550, N15549, N15548, N15547, N15546, N15545, N15544, N15543, N15542, N15541, N15540, N15539, N15538, N15537, N15536, N15535, N15534, N15533, N15532, N15531, N15530, N15529, N15528, N15527, N15526, N15525, N15524, N15523, N15522, N15521, N15520, N15519, N15518, N15517, N15516, N15515, N15514, N15513, N15512, N15511, N15510, N15509, N15508, N15507, N15506, N15505, N15504, N15503, N15502, N15501, N15500, N15499, N15498, N15497, N15496, N15495, N15494, N15493, N15492, N15491, N15490, N15489, N15488, N15487, N15486, N15485, N15484, N15483, N15482, N15481, N15480, N15479, N15478, N15477, N15476, N15475, N15474, N15473, N15472, N15471, N15470, N15469, N15468, N15467, N15466, N15465, N15464, N15463, N15462, N15461, N15460, N15459, N15458, N15457, N15456, N15455, N15454, N15453, N15452, N15451, N15450, N15449, N15448, N15447, N15446, N15445, N15444, N15443, N15442, N15441, N15440, N15439, N15438, N15437, N15436, N15435, N15434, N15433, N15432, N15431, N15430, N15429, N15428, N15427, N15426, N15425, N15424, N15423, N15422, N15421, N15420, N15419, N15418, N15417, N15416, N15415, N15414, N15413, N15412, N15411, N15410, N15409, N15408, N15407, N15406, N15405, N15404, N15403, N15402, N15401, N15400, N15399, N15398, N15397, N15396, N15395, N15394, N15393, N15392, N15391, N15390, N15389, N15388, N15387, N15386, N15385, N15384, N15383, N15382, N15381, N15380, N15379, N15378, N15377, N15376, N15375, N15374, N15373, N15372, N15371, N15370, N15369, N15368, N15367, N15366, N15365, N15364, N15363, N15362, N15361, N15360, N15359, N15358, N15357, N15356, N15355, N15354, N15353, N15352, N15351, N15350, N15349, N15348, N15347, N15346, N15345, N15344, N15343, N15342, N15341, N15340, N15339, N15338, N15337, N15336, N15335, N15334, N15333, N15332, N15331, N15330, N15329, N15328, N15327, N15326, N15325, N15324, N15323, N15322, N15321, N15320, N15319, N15318, N15317, N15316, N15315, N15314, N15313, N15312, N15311, N15310, N15309, N15308, N15307, N15306, N15305, N15304, N15303, N15302, N15301, N15300, N15299, N15298, N15297, N15296, N15295, N15294, N15293, N15292, N15291, N15290, N15289, N15288, N15287, N15286, N15285, N15284, N15283, N15282, N15281, N15280, N15279, N15278, N15277, N15276, N15275, N15274, N15273, N15272, N15271, N15270, N15269, N15268, N15267, N15266, N15265, N15264, N15263, N15262, N15261, N15260 } = (N179)? { N14223, N14222, N14221, N14220, N14219, N14218, N14217, N14216, N14215, N14214, N14213, N14212, N14211, N14210, N14209, N14208, N14207, N14206, N14205, N14204, N14203, N14202, N14201, N14200, N14199, N14198, N14197, N14196, N14195, N14194, N14193, N14192, N14191, N14190, N14189, N14188, N14187, N14186, N14185, N14184, N14183, N14182, N14181, N14180, N14179, N14178, N14177, N14176, N14175, N14174, N14173, N14172, N14171, N14170, N14169, N14168, N14167, N14166, N14165, N14164, N14163, N14162, N14161, N14160, N14159, N14158, N14157, N14156, N14155, N14154, N14153, N14152, N14151, N14150, N14149, N14148, N14147, N14146, N14145, N14144, N14143, N14142, N14141, N14140, N14139, N14138, N14137, N14136, N14135, N14134, N14133, N14132, N14131, N14130, N14129, N14128, N14127, N14126, N14125, N14124, N14123, N14122, N14121, N14120, N14119, N14118, N14117, N14116, N14115, N14114, N14113, N14112, N14111, N14110, N14109, N14108, N14107, N14106, N14105, N14104, N14103, N14102, N14101, N14100, N14099, N14098, N14097, N14096, N14095, N14094, N14093, N14092, N14091, N14090, N14089, N14088, N14087, N14086, N14085, N14084, N14083, N14082, N14081, N14080, N14079, N14078, N14077, N14076, N14075, N14074, N14073, N14072, N14071, N14070, N14069, N14068, N14067, N14066, N14065, N14064, N14063, N14062, N14061, N14060, N14059, N14058, N14057, N14056, N14055, N14054, N14053, N14052, N14051, N14050, N14049, N14048, N14047, N14046, N14045, N14044, N14043, N14042, N14041, N14040, N14039, N14038, N14037, N14036, N14035, N14034, N14033, N14032, N14031, N14030, N14029, N14028, N14027, N14026, N14025, N14024, N14023, N14022, N14021, N14020, N14019, N14018, N14017, N14016, N14015, N14014, N14013, N14012, N14011, N14010, N14009, N14008, N14007, N14006, N14005, N14004, N14003, N14002, N14001, N14000, N13999, N13998, N13997, N13996, N13995, N13994, N13993, N13992, N13991, N13990, N13989, N13988, N13987, N13986, N13985, N13984, N13983, N13982, N13981, N13980, N13979, N13978, N13977, N13976, N13975, N13974, N13973, N13972, N13971, N13970, N13969, N13968, N13967, N13966, N13965, N13964, N13963, N13962, N13961, N13960, N13959, N13958, N13957, N13956, N13955, N13954, N13953, N13952, N13951, N13950, N13949, N13948, N13947, N13946, N13945, N13944, N13943, N13942, N13941, N13940, N13939, N13938, N13937, N13936, N13935, N13934, N13933, N13932, N13931, N13930, N13929, N13928, N13927, N13926, N13925, N13924, N13923, N13922, N13921, N13920, N13919, N13918, N13917, N13916, N13915, N13914, N13913, N13912, N13911, N13910, N13909, N13908, N13907, N13906, N13905, N13904, N13903, N13902, N13901, N13900, N13899, N13898, N13897, N13896, N13895, N13894, N13893, N13892, N13891, N13890, N13889, N13888, N13887, N13886, N13885, N13884, N13883, N13882, N13881, N13880, N13879, N13878, N13877, N13876, N13875, N13874, N13873, N13872, N13871, N13870, N13869, N13868, N13867, N13866, N13865, N13864, N13863, N13862, N13861, N13860, N13859, N13858, N13857, N13856, N13855, N13854, N13853, N13852, N13851, N13850, N13849, N13848, N13847, N13846, N13845, N13844, N13843, N13842, N13841, N13840, N13839, N13838, N13837, N13836, N13835, N13834, N13833, N13832, N13831, N13830, N13829, N13828, N13827, N13826, N13825, N13824, N13823, N13822, N13821, N13820, N13819, N13818, N13817, N13816, N13815, N13814, N13813, N13812, N13811, N13810, N13809, N13808, N13807, N13806, N13805, N13804, N13803, N13802, N13801, N13800, N13799, N13798, N13797, N13796, N13795, N13794, N13793, N13792, N13791, N13790, N13789, N13788, N13787, N13786, N13785, N13784, N13783, N13782, N13781, N13780, N13779, N13778, N13777, N13776, N13775, N13774, N13773, N13772, N13771, N13770, N13769, N13768, N13767, N13766, N13765, N13764, N13763, N13762, N13761, N13760, N13759, N13758, N13757, N13756, N13755, N13754, N13753, N13752, N13751, N13750, N13749, N13748, N13747, N13746, N13745, N13744, N13743, N13742, N13741, N13740, N13739, N13738, N13737, N13736, N13735, N13734, N13733, N13732, N13731, N13730, N13729, N13728, N13727, N13726, N13725, N13724, N13723, N13722, N13721, N13720, N13719, N13718, N13717, N13716, N13715, N13714, N13713, N13712, N13711, N13710, N13709, N13708, N13707, N13706, N13705, N13704, N13703, N13702, N13701, N13700, N13699, N13698, N13697, N13696, N13695, N13694, N13693, N13692, N13691, N13690, N13689, N13688, N13687, N13686, N13685, N13684, N13683, N13682, N13681, N13680, N13679, N13678, N13677, N13676, N13675, N13674, N13673, N13672, N13671, N13670, N13669, N13668, N13667, N13666, N13665, N13664, N13663, N13662, N13661, N13660, N13659, N13658, N13657, N13656, N13655, N13654, N13653, N13652, N13651, N13650, N13649, N13648, N13647, N13646, N13645, N13644, N13643, N13642, N13641, N13640, N13639, N13638, N13637, N13636, N13635, N13634, N13633, N13632, N13631, N13630, N13629, N13628, N13627, N13626, N13625, N13624, N13623, N13622, N13621, N13620, N13619, N13618, N13617, N13616, N13615, N13614, N13613, N13612, N13611, N13610, N13609, N13608, N13607, N13606, N13605, N13604, N13603, N13602, N13601, N13600, N13599, N13598, N13597, N13596, N13595, N13594, N13593, N13592, N13591, N13590, N13589, N13588, N13587, N13586, N13585, N13584, N13583, N13582, N13581, N13580, N13579, N13578, N13577, N13576, N13575, N13574, N13573, N13572, N13571, N13570, N13569, N13568, N13567, N13566, N13565, N13564, N13563, N13562, N13561, N13560, N13559, N13558, N13557, N13556, N13555, N13554, N13553, N13552, N13551, N13550, N13549, N13548, N13547, N13546, N13545, N13544, N13543, N13542, N13541, N13540, N13539, N13538, N13537, N13536, N13535, N13534, N13533, N13532, N13531, N13530, N13529, N13528, N13527, N13526, N13525, N13524, N13523, N13522, N13521, N13520, N13519, N13518, N13517, N13516, N13515, N13514, N13513, N13512, N13511, N13510, N13509, N13508, N13507, N13506, N13505, N13504, N13503, N13502, N13501, N13500, N13499, N13498, N13497, N13496, N13495, N13494, N13493, N13492, N13491, N13490, N13489, N13488, N13487, N13486, N13485, N13484, N13483, N13482, N13481, N13480, N13479, N13478, N13477, N13476, N13475, N13474, N13473, N13472, N13471, N13470, N13469, N13468, N13467, N13466, N13465, N13464, N13463, N13462, N13461, N13460, N13459, N13458, N13457, N13456, N13455, N13454, N13453, N13452, N13451, N13450, N13449, N13448, N13447, N13446, N13445, N13444, N13443, N13442, N13441, N13440, N13439, N13438, N13437, N13436, N13435, N13434, N13433, N13432, N13431, N13430, N13429, N13428, N13427, N13426, N13425, N13424, N13423, N13422, N13421, N13420, N13419, N13418, N13417, N13416, N13415, N13414, N13413, N13412, N13411, N13410, N13409, N13408, N13407, N13406, N13405, N13404, N13403, N13402, N13401, N13400, N13399, N13398, N13397, N13396, N13395, N13394, N13393, N13392, N13391, N13390, N13389, N13388, N13387, N13386, N13385, N13384, N13383, N13382, N13381, N13380, N13379, N13378, N13377, N13376, N13375, N13374, N13373, N13372, N13371, N13370, N13369, N13368, N13367, N13366, N13365, N13364, N13363, N13362, N13361, N13360, N13359, N13358, N13357, N13356, N13355, N13354, N13353, N13352, N13351, N13350, N13349, N13348, N13347, N13346, N13345, N13344, N13343, N13342, N13341, N13340, N13339, N13338, N13337, N13336, N13335, N13334, N13333, N13332, N13331, N13330, N13329, N13328, N13327, N13326, N13325, N13324, N13323, N13322, N13321, N13320, N13319, N13318, N13317, N13316, N13315, N13314, N13313, N13312, N13311, N13310, N13309, N13308, N13307, N13306, N13305, N13304, N13303, N13302, N13301, N13300, N13299, N13298, N13297, N13296, N13295, N13294, N13293, N13292, N13291, N13290, N13289, N13288, N13287, N13286, N13285, N13284, N13283, N13282, N13281, N13280, N13279, N13278, N13277, N13276, N13275, N13274, N13273, N13272, N13271, N13270, N13269, N13268, N13267, N13266, N13265, N13264, N13263, N13262, N13261, N13260, N13259, N13258, N13257, N13256, N13255, N13254, N13253, N13252, N13251, N13250, N13249, N13248, N13247, N13246, N13245, N13244, N13243, N13242, N13241, N13240, N13239, N13238, N13237, N13236, N13235, N13234, N13233, N13232, N13231, N13230, N13229, N13228, N13227, N13226, N13225, N13224, N13223, N13222, N13221, N13220, N13219, N13218, N13217, N13216, N13215, N13214, N13213, N13212, N13211, N13210, N13209, N13208, N13207, N13206, N13205, N13204, N13203, N13202, N13201, N13200, N13199, N13198, N13197, N13196, N13195, N13194, N13193, N13192 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N13191)? { N15259, N15258, N15257, N15256, N15255, N15254, N15253, N15252, N15251, N15250, N15249, N15248, N15247, N15246, N15245, N15244, N15243, N15242, N15241, N15240, N15239, N15238, N15237, N15236, N15235, N15234, N15233, N15232, N15231, N15230, N15229, N15228, N15227, N15226, N15225, N15224, N15223, N15222, N15221, N15220, N15219, N15218, N15217, N15216, N15215, N15214, N15213, N15212, N15211, N15210, N15209, N15208, N15207, N15206, N15205, N15204, N15203, N15202, N15201, N15200, N15199, N15198, N15197, N15196, N11991, N11990, N11989, N11988, N11987, N11986, N11985, N11984, N11983, N11982, N11981, N11980, N11979, N11978, N11977, N11976, N11975, N11974, N11973, N11972, N11971, N11970, N11969, N11968, N11967, N11966, N11965, N11964, N11963, N11962, N11961, N11960, N11959, N11958, N11957, N11956, N11955, N11954, N11953, N11952, N11951, N11950, N11949, N11948, N11947, N11946, N11945, N11944, N11943, N11942, N11941, N11940, N11939, N11938, N11937, N11936, N11935, N11934, N11933, N11932, N11931, N11930, N11929, N11928, N11927, N15195, N15194, N15193, N15192, N15191, N15190, N15189, N15188, N15187, N15186, N15185, N15184, N15183, N15182, N15181, N15180, N15179, N15178, N15177, N15176, N15175, N15174, N15173, N15172, N15171, N15170, N15169, N15168, N15167, N15166, N15165, N15164, N15163, N15162, N15161, N15160, N15159, N15158, N15157, N15156, N15155, N15154, N15153, N15152, N15151, N15150, N15149, N15148, N15147, N15146, N15145, N15144, N15143, N15142, N15141, N15140, N15139, N15138, N15137, N15136, N15135, N15134, N15133, N15132, N11733, N11732, N11731, N11730, N11729, N11728, N11727, N11726, N11725, N11724, N11723, N11722, N11721, N11720, N11719, N11718, N11717, N11716, N11715, N11714, N11713, N11712, N11711, N11710, N11709, N11708, N11707, N11706, N11705, N11704, N11703, N11702, N11701, N11700, N11699, N11698, N11697, N11696, N11695, N11694, N11693, N11692, N11691, N11690, N11689, N11688, N11687, N11686, N11685, N11684, N11683, N11682, N11681, N11680, N11679, N11678, N11677, N11676, N11675, N11674, N11673, N11672, N11671, N11670, N11669, N15131, N15130, N15129, N15128, N15127, N15126, N15125, N15124, N15123, N15122, N15121, N15120, N15119, N15118, N15117, N15116, N15115, N15114, N15113, N15112, N15111, N15110, N15109, N15108, N15107, N15106, N15105, N15104, N15103, N15102, N15101, N15100, N15099, N15098, N15097, N15096, N15095, N15094, N15093, N15092, N15091, N15090, N15089, N15088, N15087, N15086, N15085, N15084, N15083, N15082, N15081, N15080, N15079, N15078, N15077, N15076, N15075, N15074, N15073, N15072, N15071, N15070, N15069, N15068, N11475, N11474, N11473, N11472, N11471, N11470, N11469, N11468, N11467, N11466, N11465, N11464, N11463, N11462, N11461, N11460, N11459, N11458, N11457, N11456, N11455, N11454, N11453, N11452, N11451, N11450, N11449, N11448, N11447, N11446, N11445, N11444, N11443, N11442, N11441, N11440, N11439, N11438, N11437, N11436, N11435, N11434, N11433, N11432, N11431, N11430, N11429, N11428, N11427, N11426, N11425, N11424, N11423, N11422, N11421, N11420, N11419, N11418, N11417, N11416, N11415, N11414, N11413, N11412, N11411, N15067, N15066, N15065, N15064, N15063, N15062, N15061, N15060, N15059, N15058, N15057, N15056, N15055, N15054, N15053, N15052, N15051, N15050, N15049, N15048, N15047, N15046, N15045, N15044, N15043, N15042, N15041, N15040, N15039, N15038, N15037, N15036, N15035, N15034, N15033, N15032, N15031, N15030, N15029, N15028, N15027, N15026, N15025, N15024, N15023, N15022, N15021, N15020, N15019, N15018, N15017, N15016, N15015, N15014, N15013, N15012, N15011, N15010, N15009, N15008, N15007, N15006, N15005, N15004, N11217, N11216, N11215, N11214, N11213, N11212, N11211, N11210, N11209, N11208, N11207, N11206, N11205, N11204, N11203, N11202, N11201, N11200, N11199, N11198, N11197, N11196, N11195, N11194, N11193, N11192, N11191, N11190, N11189, N11188, N11187, N11186, N11185, N11184, N11183, N11182, N11181, N11180, N11179, N11178, N11177, N11176, N11175, N11174, N11173, N11172, N11171, N11170, N11169, N11168, N11167, N11166, N11165, N11164, N11163, N11162, N11161, N11160, N11159, N11158, N11157, N11156, N11155, N11154, N11153, N15003, N15002, N15001, N15000, N14999, N14998, N14997, N14996, N14995, N14994, N14993, N14992, N14991, N14990, N14989, N14988, N14987, N14986, N14985, N14984, N14983, N14982, N14981, N14980, N14979, N14978, N14977, N14976, N14975, N14974, N14973, N14972, N14971, N14970, N14969, N14968, N14967, N14966, N14965, N14964, N14963, N14962, N14961, N14960, N14959, N14958, N14957, N14956, N14955, N14954, N14953, N14952, N14951, N14950, N14949, N14948, N14947, N14946, N14945, N14944, N14943, N14942, N14941, N14940, N10959, N10958, N10957, N10956, N10955, N10954, N10953, N10952, N10951, N10950, N10949, N10948, N10947, N10946, N10945, N10944, N10943, N10942, N10941, N10940, N10939, N10938, N10937, N10936, N10935, N10934, N10933, N10932, N10931, N10930, N10929, N10928, N10927, N10926, N10925, N10924, N10923, N10922, N10921, N10920, N10919, N10918, N10917, N10916, N10915, N10914, N10913, N10912, N10911, N10910, N10909, N10908, N10907, N10906, N10905, N10904, N10903, N10902, N10901, N10900, N10899, N10898, N10897, N10896, N10895, N14939, N14938, N14937, N14936, N14935, N14934, N14933, N14932, N14931, N14930, N14929, N14928, N14927, N14926, N14925, N14924, N14923, N14922, N14921, N14920, N14919, N14918, N14917, N14916, N14915, N14914, N14913, N14912, N14911, N14910, N14909, N14908, N14907, N14906, N14905, N14904, N14903, N14902, N14901, N14900, N14899, N14898, N14897, N14896, N14895, N14894, N14893, N14892, N14891, N14890, N14889, N14888, N14887, N14886, N14885, N14884, N14883, N14882, N14881, N14880, N14879, N14878, N14877, N14876, N10701, N10700, N10699, N10698, N10697, N10696, N10695, N10694, N10693, N10692, N10691, N10690, N10689, N10688, N10687, N10686, N10685, N10684, N10683, N10682, N10681, N10680, N10679, N10678, N10677, N10676, N10675, N10674, N10673, N10672, N10671, N10670, N10669, N10668, N10667, N10666, N10665, N10664, N10663, N10662, N10661, N10660, N10659, N10658, N10657, N10656, N10655, N10654, N10653, N10652, N10651, N10650, N10649, N10648, N10647, N10646, N10645, N10644, N10643, N10642, N10641, N10640, N10639, N10638, N10637, N14875, N14874, N14873, N14872, N14871, N14870, N14869, N14868, N14867, N14866, N14865, N14864, N14863, N14862, N14861, N14860, N14859, N14858, N14857, N14856, N14855, N14854, N14853, N14852, N14851, N14850, N14849, N14848, N14847, N14846, N14845, N14844, N14843, N14842, N14841, N14840, N14839, N14838, N14837, N14836, N14835, N14834, N14833, N14832, N14831, N14830, N14829, N14828, N14827, N14826, N14825, N14824, N14823, N14822, N14821, N14820, N14819, N14818, N14817, N14816, N14815, N14814, N14813, N14812, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422, N10421, N10420, N10419, N10418, N10417, N10416, N10415, N10414, N10413, N10412, N10411, N10410, N10409, N10408, N10407, N10406, N10405, N10404, N10403, N10402, N10401, N10400, N10399, N10398, N10397, N10396, N10395, N10394, N10393, N10392, N10391, N10390, N10389, N10388, N10387, N10386, N10385, N10384, N10383, N10382, N10381, N10380, N10379, N14811, N14810, N14809, N14808, N14807, N14806, N14805, N14804, N14803, N14802, N14801, N14800, N14799, N14798, N14797, N14796, N14795, N14794, N14793, N14792, N14791, N14790, N14789, N14788, N14787, N14786, N14785, N14784, N14783, N14782, N14781, N14780, N14779, N14778, N14777, N14776, N14775, N14774, N14773, N14772, N14771, N14770, N14769, N14768, N14767, N14766, N14765, N14764, N14763, N14762, N14761, N14760, N14759, N14758, N14757, N14756, N14755, N14754, N14753, N14752, N14751, N14750, N14749, N14748, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121 } : 1'b0;
  assign N179 = ex_i[129];
  assign { N18355, N18354, N18353, N18352, N18351, N18350, N18349, N18348, N18347, N18346, N18345, N18344, N18343, N18342, N18341, N18340, N18339, N18338, N18337, N18336, N18335, N18334, N18333, N18332, N18331, N18330, N18329, N18328, N18327, N18326, N18325, N18324, N18323, N18322, N18321, N18320, N18319, N18318, N18317, N18316, N18315, N18314, N18313, N18312, N18311, N18310, N18309, N18308, N18307, N18306, N18305, N18304, N18303, N18302, N18301, N18300, N18299, N18298, N18297, N18296, N18295, N18294, N18293, N18292, N18291, N18290, N18289, N18288, N18287, N18286, N18285, N18284, N18283, N18282, N18281, N18280, N18279, N18278, N18277, N18276, N18275, N18274, N18273, N18272, N18271, N18270, N18269, N18268, N18267, N18266, N18265, N18264, N18263, N18262, N18261, N18260, N18259, N18258, N18257, N18256, N18255, N18254, N18253, N18252, N18251, N18250, N18249, N18248, N18247, N18246, N18245, N18244, N18243, N18242, N18241, N18240, N18239, N18238, N18237, N18236, N18235, N18234, N18233, N18232, N18231, N18230, N18229, N18228, N18227, N18226, N18225, N18224, N18223, N18222, N18221, N18220, N18219, N18218, N18217, N18216, N18215, N18214, N18213, N18212, N18211, N18210, N18209, N18208, N18207, N18206, N18205, N18204, N18203, N18202, N18201, N18200, N18199, N18198, N18197, N18196, N18195, N18194, N18193, N18192, N18191, N18190, N18189, N18188, N18187, N18186, N18185, N18184, N18183, N18182, N18181, N18180, N18179, N18178, N18177, N18176, N18175, N18174, N18173, N18172, N18171, N18170, N18169, N18168, N18167, N18166, N18165, N18164, N18163, N18162, N18161, N18160, N18159, N18158, N18157, N18156, N18155, N18154, N18153, N18152, N18151, N18150, N18149, N18148, N18147, N18146, N18145, N18144, N18143, N18142, N18141, N18140, N18139, N18138, N18137, N18136, N18135, N18134, N18133, N18132, N18131, N18130, N18129, N18128, N18127, N18126, N18125, N18124, N18123, N18122, N18121, N18120, N18119, N18118, N18117, N18116, N18115, N18114, N18113, N18112, N18111, N18110, N18109, N18108, N18107, N18106, N18105, N18104, N18103, N18102, N18101, N18100, N18099, N18098, N18097, N18096, N18095, N18094, N18093, N18092, N18091, N18090, N18089, N18088, N18087, N18086, N18085, N18084, N18083, N18082, N18081, N18080, N18079, N18078, N18077, N18076, N18075, N18074, N18073, N18072, N18071, N18070, N18069, N18068, N18067, N18066, N18065, N18064, N18063, N18062, N18061, N18060, N18059, N18058, N18057, N18056, N18055, N18054, N18053, N18052, N18051, N18050, N18049, N18048, N18047, N18046, N18045, N18044, N18043, N18042, N18041, N18040, N18039, N18038, N18037, N18036, N18035, N18034, N18033, N18032, N18031, N18030, N18029, N18028, N18027, N18026, N18025, N18024, N18023, N18022, N18021, N18020, N18019, N18018, N18017, N18016, N18015, N18014, N18013, N18012, N18011, N18010, N18009, N18008, N18007, N18006, N18005, N18004, N18003, N18002, N18001, N18000, N17999, N17998, N17997, N17996, N17995, N17994, N17993, N17992, N17991, N17990, N17989, N17988, N17987, N17986, N17985, N17984, N17983, N17982, N17981, N17980, N17979, N17978, N17977, N17976, N17975, N17974, N17973, N17972, N17971, N17970, N17969, N17968, N17967, N17966, N17965, N17964, N17963, N17962, N17961, N17960, N17959, N17958, N17957, N17956, N17955, N17954, N17953, N17952, N17951, N17950, N17949, N17948, N17947, N17946, N17945, N17944, N17943, N17942, N17941, N17940, N17939, N17938, N17937, N17936, N17935, N17934, N17933, N17932, N17931, N17930, N17929, N17928, N17927, N17926, N17925, N17924, N17923, N17922, N17921, N17920, N17919, N17918, N17917, N17916, N17915, N17914, N17913, N17912, N17911, N17910, N17909, N17908, N17907, N17906, N17905, N17904, N17903, N17902, N17901, N17900, N17899, N17898, N17897, N17896, N17895, N17894, N17893, N17892, N17891, N17890, N17889, N17888, N17887, N17886, N17885, N17884, N17883, N17882, N17881, N17880, N17879, N17878, N17877, N17876, N17875, N17874, N17873, N17872, N17871, N17870, N17869, N17868, N17867, N17866, N17865, N17864, N17863, N17862, N17861, N17860, N17859, N17858, N17857, N17856, N17855, N17854, N17853, N17852, N17851, N17850, N17849, N17848, N17847, N17846, N17845, N17844, N17843, N17842, N17841, N17840, N17839, N17838, N17837, N17836, N17835, N17834, N17833, N17832, N17831, N17830, N17829, N17828, N17827, N17826, N17825, N17824, N17823, N17822, N17821, N17820, N17819, N17818, N17817, N17816, N17815, N17814, N17813, N17812, N17811, N17810, N17809, N17808, N17807, N17806, N17805, N17804, N17803, N17802, N17801, N17800, N17799, N17798, N17797, N17796, N17795, N17794, N17793, N17792, N17791, N17790, N17789, N17788, N17787, N17786, N17785, N17784, N17783, N17782, N17781, N17780, N17779, N17778, N17777, N17776, N17775, N17774, N17773, N17772, N17771, N17770, N17769, N17768, N17767, N17766, N17765, N17764, N17763, N17762, N17761, N17760, N17759, N17758, N17757, N17756, N17755, N17754, N17753, N17752, N17751, N17750, N17749, N17748, N17747, N17746, N17745, N17744, N17743, N17742, N17741, N17740, N17739, N17738, N17737, N17736, N17735, N17734, N17733, N17732, N17731, N17730, N17729, N17728, N17727, N17726, N17725, N17724, N17723, N17722, N17721, N17720, N17719, N17718, N17717, N17716, N17715, N17714, N17713, N17712, N17711, N17710, N17709, N17708, N17707, N17706, N17705, N17704, N17703, N17702, N17701, N17700, N17699, N17698, N17697, N17696, N17695, N17694, N17693, N17692, N17691, N17690, N17689, N17688, N17687, N17686, N17685, N17684, N17683, N17682, N17681, N17680, N17679, N17678, N17677, N17676, N17675, N17674, N17673, N17672, N17671, N17670, N17669, N17668, N17667, N17666, N17665, N17664, N17663, N17662, N17661, N17660, N17659, N17658, N17657, N17656, N17655, N17654, N17653, N17652, N17651, N17650, N17649, N17648, N17647, N17646, N17645, N17644, N17643, N17642, N17641, N17640, N17639, N17638, N17637, N17636, N17635, N17634, N17633, N17632, N17631, N17630, N17629, N17628, N17627, N17626, N17625, N17624, N17623, N17622, N17621, N17620, N17619, N17618, N17617, N17616, N17615, N17614, N17613, N17612, N17611, N17610, N17609, N17608, N17607, N17606, N17605, N17604, N17603, N17602, N17601, N17600, N17599, N17598, N17597, N17596, N17595, N17594, N17593, N17592, N17591, N17590, N17589, N17588, N17587, N17586, N17585, N17584, N17583, N17582, N17581, N17580, N17579, N17578, N17577, N17576, N17575, N17574, N17573, N17572, N17571, N17570, N17569, N17568, N17567, N17566, N17565, N17564, N17563, N17562, N17561, N17560, N17559, N17558, N17557, N17556, N17555, N17554, N17553, N17552, N17551, N17550, N17549, N17548, N17547, N17546, N17545, N17544, N17543, N17542, N17541, N17540, N17539, N17538, N17537, N17536, N17535, N17534, N17533, N17532, N17531, N17530, N17529, N17528, N17527, N17526, N17525, N17524, N17523, N17522, N17521, N17520, N17519, N17518, N17517, N17516, N17515, N17514, N17513, N17512, N17511, N17510, N17509, N17508, N17507, N17506, N17505, N17504, N17503, N17502, N17501, N17500, N17499, N17498, N17497, N17496, N17495, N17494, N17493, N17492, N17491, N17490, N17489, N17488, N17487, N17486, N17485, N17484, N17483, N17482, N17481, N17480, N17479, N17478, N17477, N17476, N17475, N17474, N17473, N17472, N17471, N17470, N17469, N17468, N17467, N17466, N17465, N17464, N17463, N17462, N17461, N17460, N17459, N17458, N17457, N17456, N17455, N17454, N17453, N17452, N17451, N17450, N17449, N17448, N17447, N17446, N17445, N17444, N17443, N17442, N17441, N17440, N17439, N17438, N17437, N17436, N17435, N17434, N17433, N17432, N17431, N17430, N17429, N17428, N17427, N17426, N17425, N17424, N17423, N17422, N17421, N17420, N17419, N17418, N17417, N17416, N17415, N17414, N17413, N17412, N17411, N17410, N17409, N17408, N17407, N17406, N17405, N17404, N17403, N17402, N17401, N17400, N17399, N17398, N17397, N17396, N17395, N17394, N17393, N17392, N17391, N17390, N17389, N17388, N17387, N17386, N17385, N17384, N17383, N17382, N17381, N17380, N17379, N17378, N17377, N17376, N17375, N17374, N17373, N17372, N17371, N17370, N17369, N17368, N17367, N17366, N17365, N17364, N17363, N17362, N17361, N17360, N17359, N17358, N17357, N17356, N17355, N17354, N17353, N17352, N17351, N17350, N17349, N17348, N17347, N17346, N17345, N17344, N17343, N17342, N17341, N17340, N17339, N17338, N17337, N17336, N17335, N17334, N17333, N17332, N17331, N17330, N17329, N17328, N17327, N17326, N17325, N17324, N17323, N17322, N17321, N17320, N17319, N17318, N17317, N17316, N17315, N17314, N17313, N17312, N17311, N17310, N17309, N17308, N17307, N17306, N17305, N17304, N17303, N17302, N17301, N17300, N17299, N17298, N17297, N17296, N17295, N17294, N17293, N17292, N17291, N17290, N17289, N17288, N17287, N17286, N17285, N17284, N17283, N17282, N17281, N17280, N17279, N17278, N17277, N17276, N17275, N17274, N17273, N17272, N17271, N17270, N17269, N17268, N17267, N17266, N17265, N17264, N17263, N17262, N17261, N17260, N17259, N17258, N17257, N17256, N17255, N17254, N17253, N17252, N17251, N17250, N17249, N17248, N17247, N17246, N17245, N17244, N17243, N17242, N17241, N17240, N17239, N17238, N17237, N17236, N17235, N17234, N17233, N17232, N17231, N17230, N17229, N17228, N17227, N17226, N17225, N17224, N17223, N17222, N17221, N17220, N17219, N17218, N17217, N17216, N17215, N17214, N17213, N17212, N17211, N17210, N17209, N17208, N17207, N17206, N17205, N17204, N17203, N17202, N17201, N17200, N17199, N17198, N17197, N17196, N17195, N17194, N17193, N17192, N17191, N17190, N17189, N17188, N17187, N17186, N17185, N17184, N17183, N17182, N17181, N17180, N17179, N17178, N17177, N17176, N17175, N17174, N17173, N17172, N17171, N17170, N17169, N17168, N17167, N17166, N17165, N17164, N17163, N17162, N17161, N17160, N17159, N17158, N17157, N17156, N17155, N17154, N17153, N17152, N17151, N17150, N17149, N17148, N17147, N17146, N17145, N17144, N17143, N17142, N17141, N17140, N17139, N17138, N17137, N17136, N17135, N17134, N17133, N17132, N17131, N17130, N17129, N17128, N17127, N17126, N17125, N17124, N17123, N17122, N17121, N17120, N17119, N17118, N17117, N17116, N17115, N17114, N17113, N17112, N17111, N17110, N17109, N17108, N17107, N17106, N17105, N17104, N17103, N17102, N17101, N17100, N17099, N17098, N17097, N17096, N17095, N17094, N17093, N17092, N17091, N17090, N17089, N17088, N17087, N17086, N17085, N17084, N17083, N17082, N17081, N17080, N17079, N17078, N17077, N17076, N17075, N17074, N17073, N17072, N17071, N17070, N17069, N17068, N17067, N17066, N17065, N17064, N17063, N17062, N17061, N17060, N17059, N17058, N17057, N17056, N17055, N17054, N17053, N17052, N17051, N17050, N17049, N17048, N17047, N17046, N17045, N17044, N17043, N17042, N17041, N17040, N17039, N17038, N17037, N17036, N17035, N17034, N17033, N17032, N17031, N17030, N17029, N17028, N17027, N17026, N17025, N17024, N17023, N17022, N17021, N17020, N17019, N17018, N17017, N17016, N17015, N17014, N17013, N17012, N17011, N17010, N17009, N17008, N17007, N17006, N17005, N17004, N17003, N17002, N17001, N17000, N16999, N16998, N16997, N16996, N16995, N16994, N16993, N16992, N16991, N16990, N16989, N16988, N16987, N16986, N16985, N16984, N16983, N16982, N16981, N16980, N16979, N16978, N16977, N16976, N16975, N16974, N16973, N16972, N16971, N16970, N16969, N16968, N16967, N16966, N16965, N16964, N16963, N16962, N16961, N16960, N16959, N16958, N16957, N16956, N16955, N16954, N16953, N16952, N16951, N16950, N16949, N16948, N16947, N16946, N16945, N16944, N16943, N16942, N16941, N16940, N16939, N16938, N16937, N16936, N16935, N16934, N16933, N16932, N16931, N16930, N16929, N16928, N16927, N16926, N16925, N16924, N16923, N16922, N16921, N16920, N16919, N16918, N16917, N16916, N16915, N16914, N16913, N16912, N16911, N16910, N16909, N16908, N16907, N16906, N16905, N16904, N16903, N16902, N16901, N16900, N16899, N16898, N16897, N16896, N16895, N16894, N16893, N16892, N16891, N16890, N16889, N16888, N16887, N16886, N16885, N16884, N16883, N16882, N16881, N16880, N16879, N16878, N16877, N16876, N16875, N16874, N16873, N16872, N16871, N16870, N16869, N16868, N16867, N16866, N16865, N16864, N16863, N16862, N16861, N16860, N16859, N16858, N16857, N16856, N16855, N16854, N16853, N16852, N16851, N16850, N16849, N16848, N16847, N16846, N16845, N16844, N16843, N16842, N16841, N16840, N16839, N16838, N16837, N16836, N16835, N16834, N16833, N16832, N16831, N16830, N16829, N16828, N16827, N16826, N16825, N16824, N16823, N16822, N16821, N16820, N16819, N16818, N16817, N16816, N16815, N16814, N16813, N16812, N16811, N16810, N16809, N16808, N16807, N16806, N16805, N16804, N16803, N16802, N16801, N16800, N16799, N16798, N16797, N16796, N16795, N16794, N16793, N16792, N16791, N16790, N16789, N16788, N16787, N16786, N16785, N16784, N16783, N16782, N16781, N16780, N16779, N16778, N16777, N16776, N16775, N16774, N16773, N16772, N16771, N16770, N16769, N16768, N16767, N16766, N16765, N16764, N16763, N16762, N16761, N16760, N16759, N16758, N16757, N16756, N16755, N16754, N16753, N16752, N16751, N16750, N16749, N16748, N16747, N16746, N16745, N16744, N16743, N16742, N16741, N16740, N16739, N16738, N16737, N16736, N16735, N16734, N16733, N16732, N16731, N16730, N16729, N16728, N16727, N16726, N16725, N16724, N16723, N16722, N16721, N16720, N16719, N16718, N16717, N16716, N16715, N16714, N16713, N16712, N16711, N16710, N16709, N16708, N16707, N16706, N16705, N16704, N16703, N16702, N16701, N16700, N16699, N16698, N16697, N16696, N16695, N16694, N16693, N16692, N16691, N16690, N16689, N16688, N16687, N16686, N16685, N16684, N16683, N16682, N16681, N16680, N16679, N16678, N16677, N16676, N16675, N16674, N16673, N16672, N16671, N16670, N16669, N16668, N16667, N16666, N16665, N16664, N16663, N16662, N16661, N16660, N16659, N16658, N16657, N16656, N16655, N16654, N16653, N16652, N16651, N16650, N16649, N16648, N16647, N16646, N16645, N16644, N16643, N16642, N16641, N16640, N16639, N16638, N16637, N16636, N16635, N16634, N16633, N16632, N16631, N16630, N16629, N16628, N16627, N16626, N16625, N16624, N16623, N16622, N16621, N16620, N16619, N16618, N16617, N16616, N16615, N16614, N16613, N16612, N16611, N16610, N16609, N16608, N16607, N16606, N16605, N16604, N16603, N16602, N16601, N16600, N16599, N16598, N16597, N16596, N16595, N16594, N16593, N16592, N16591, N16590, N16589, N16588, N16587, N16586, N16585, N16584, N16583, N16582, N16581, N16580, N16579, N16578, N16577, N16576, N16575, N16574, N16573, N16572, N16571, N16570, N16569, N16568, N16567, N16566, N16565, N16564, N16563, N16562, N16561, N16560, N16559, N16558, N16557, N16556, N16555, N16554, N16553, N16552, N16551, N16550, N16549, N16548, N16547, N16546, N16545, N16544, N16543, N16542, N16541, N16540, N16539, N16538, N16537, N16536, N16535, N16534, N16533, N16532, N16531, N16530, N16529, N16528, N16527, N16526, N16525, N16524, N16523, N16522, N16521, N16520, N16519, N16518, N16517, N16516, N16515, N16514, N16513, N16512, N16511, N16510, N16509, N16508, N16507, N16506, N16505, N16504, N16503, N16502, N16501, N16500, N16499, N16498, N16497, N16496, N16495, N16494, N16493, N16492, N16491, N16490, N16489, N16488, N16487, N16486, N16485, N16484, N16483, N16482, N16481, N16480, N16479, N16478, N16477, N16476, N16475, N16474, N16473, N16472, N16471, N16470, N16469, N16468, N16467, N16466, N16465, N16464, N16463, N16462, N16461, N16460, N16459, N16458, N16457, N16456, N16455, N16454, N16453, N16452, N16451, N16450, N16449, N16448, N16447, N16446, N16445, N16444, N16443, N16442, N16441, N16440, N16439, N16438, N16437, N16436, N16435, N16434, N16433, N16432, N16431, N16430, N16429, N16428, N16427, N16426, N16425, N16424, N16423, N16422, N16421, N16420, N16419, N16418, N16417, N16416, N16415, N16414, N16413, N16412, N16411, N16410, N16409, N16408, N16407, N16406, N16405, N16404, N16403, N16402, N16401, N16400, N16399, N16398, N16397, N16396, N16395, N16394, N16393, N16392, N16391, N16390, N16389, N16388, N16387, N16386, N16385, N16384, N16383, N16382, N16381, N16380, N16379, N16378, N16377, N16376, N16375, N16374, N16373, N16372, N16371, N16370, N16369, N16368, N16367, N16366, N16365, N16364, N16363, N16362, N16361, N16360, N16359, N16358, N16357, N16356, N16355, N16354, N16353, N16352, N16351, N16350, N16349, N16348, N16347, N16346, N16345, N16344, N16343, N16342, N16341, N16340, N16339, N16338, N16337, N16336, N16335, N16334, N16333, N16332, N16331, N16330, N16329, N16328, N16327, N16326, N16325, N16324, N16323, N16322, N16321, N16320, N16319, N16318, N16317, N16316, N16315, N16314, N16313, N16312, N16311, N16310, N16309, N16308, N16307, N16306, N16305, N16304, N16303, N16302, N16301, N16300, N16299, N16298, N16297, N16296, N16295, N16294, N16293, N16292 } = (N180)? { N12674, N12673, N12672, N12671, N12670, N12669, N12668, N12667, N12666, N12665, N12664, N12663, N12662, N12661, N12660, N12659, N12658, N12657, N12656, N12655, N12654, N12653, N12652, N12651, N12650, N12649, N12648, N12647, N12646, N12645, N12644, N12643, N12642, N12641, N12640, N12639, N12638, N12637, N12636, N12635, N12634, N12633, N12632, N12631, N12630, N12629, N12628, N12627, N12626, N12625, N12624, N12623, N12622, N12621, N12620, N12619, N12618, N12617, N12616, N12615, N12614, N12613, N12612, N12611, N12146, N16291, N16290, N16289, N16288, N16287, N16286, N16285, N16284, N16283, N16282, N16281, N16280, N16279, N16278, N16277, N16276, N16275, N16274, N16273, N16272, N16271, N16270, N16269, N16268, N16267, N16266, N16265, N16264, N16263, N16262, N16261, N16260, N16259, N16258, N16257, N16256, N16255, N16254, N16253, N16252, N16251, N16250, N16249, N16248, N16247, N16246, N16245, N16244, N16243, N16242, N16241, N16240, N16239, N16238, N16237, N16236, N16235, N16234, N16233, N16232, N16231, N16230, N16229, N16228, N16227, N16226, N16225, N16224, N16223, N16222, N16221, N16220, N16219, N16218, N16217, N16216, N16215, N16214, N16213, N16212, N16211, N16210, N16209, N16208, N16207, N16206, N16205, N16204, N16203, N16202, N16201, N16200, N16199, N16198, N16197, N16196, N16195, N16194, N16193, N16192, N16191, N16190, N16189, N16188, N16187, N16186, N16185, N16184, N16183, N16182, N16181, N16180, N16179, N16178, N16177, N16176, N16175, N16174, N16173, N16172, N16171, N16170, N16169, N16168, N16167, N16166, N16165, N16164, N16163, N13186, N13185, N13184, N13183, N13182, N13181, N13180, N13179, N13178, N13177, N13176, N13175, N13174, N13173, N13172, N13171, N13170, N13169, N13168, N13167, N13166, N13165, N13164, N13163, N13162, N13161, N13160, N13159, N13158, N13157, N13156, N13155, N13154, N13153, N13152, N13151, N13150, N13149, N13148, N13147, N13146, N13145, N13144, N13143, N13142, N13141, N13140, N13139, N13138, N13137, N13136, N13135, N13134, N13133, N13132, N13131, N13130, N13129, N13128, N13127, N13126, N13125, N13124, N13123, N12609, N12608, N12607, N12606, N12605, N12604, N12603, N12602, N12601, N12600, N12599, N12598, N12597, N12596, N12595, N12594, N12593, N12592, N12591, N12590, N12589, N12588, N12587, N12586, N12585, N12584, N12583, N12582, N12581, N12580, N12579, N12578, N12577, N12576, N12575, N12574, N12573, N12572, N12571, N12570, N12569, N12568, N12567, N12566, N12565, N12564, N12563, N12562, N12561, N12560, N12559, N12558, N12557, N12556, N12555, N12554, N12553, N12552, N12551, N12550, N12549, N12548, N12547, N12546, N12145, N16162, N16161, N16160, N16159, N16158, N16157, N16156, N16155, N16154, N16153, N16152, N16151, N16150, N16149, N16148, N16147, N16146, N16145, N16144, N16143, N16142, N16141, N16140, N16139, N16138, N16137, N16136, N16135, N16134, N16133, N16132, N16131, N16130, N16129, N16128, N16127, N16126, N16125, N16124, N16123, N16122, N16121, N16120, N16119, N16118, N16117, N16116, N16115, N16114, N16113, N16112, N16111, N16110, N16109, N16108, N16107, N16106, N16105, N16104, N16103, N16102, N16101, N16100, N16099, N16098, N16097, N16096, N16095, N16094, N16093, N16092, N16091, N16090, N16089, N16088, N16087, N16086, N16085, N16084, N16083, N16082, N16081, N16080, N16079, N16078, N16077, N16076, N16075, N16074, N16073, N16072, N16071, N16070, N16069, N16068, N16067, N16066, N16065, N16064, N16063, N16062, N16061, N16060, N16059, N16058, N16057, N16056, N16055, N16054, N16053, N16052, N16051, N16050, N16049, N16048, N16047, N16046, N16045, N16044, N16043, N16042, N16041, N16040, N16039, N16038, N16037, N16036, N16035, N16034, N13122, N13121, N13120, N13119, N13118, N13117, N13116, N13115, N13114, N13113, N13112, N13111, N13110, N13109, N13108, N13107, N13106, N13105, N13104, N13103, N13102, N13101, N13100, N13099, N13098, N13097, N13096, N13095, N13094, N13093, N13092, N13091, N13090, N13089, N13088, N13087, N13086, N13085, N13084, N13083, N13082, N13081, N13080, N13079, N13078, N13077, N13076, N13075, N13074, N13073, N13072, N13071, N13070, N13069, N13068, N13067, N13066, N13065, N13064, N13063, N13062, N13061, N13060, N13059, N12544, N12543, N12542, N12541, N12540, N12539, N12538, N12537, N12536, N12535, N12534, N12533, N12532, N12531, N12530, N12529, N12528, N12527, N12526, N12525, N12524, N12523, N12522, N12521, N12520, N12519, N12518, N12517, N12516, N12515, N12514, N12513, N12512, N12511, N12510, N12509, N12508, N12507, N12506, N12505, N12504, N12503, N12502, N12501, N12500, N12499, N12498, N12497, N12496, N12495, N12494, N12493, N12492, N12491, N12490, N12489, N12488, N12487, N12486, N12485, N12484, N12483, N12482, N12481, N12144, N16033, N16032, N16031, N16030, N16029, N16028, N16027, N16026, N16025, N16024, N16023, N16022, N16021, N16020, N16019, N16018, N16017, N16016, N16015, N16014, N16013, N16012, N16011, N16010, N16009, N16008, N16007, N16006, N16005, N16004, N16003, N16002, N16001, N16000, N15999, N15998, N15997, N15996, N15995, N15994, N15993, N15992, N15991, N15990, N15989, N15988, N15987, N15986, N15985, N15984, N15983, N15982, N15981, N15980, N15979, N15978, N15977, N15976, N15975, N15974, N15973, N15972, N15971, N15970, N15969, N15968, N15967, N15966, N15965, N15964, N15963, N15962, N15961, N15960, N15959, N15958, N15957, N15956, N15955, N15954, N15953, N15952, N15951, N15950, N15949, N15948, N15947, N15946, N15945, N15944, N15943, N15942, N15941, N15940, N15939, N15938, N15937, N15936, N15935, N15934, N15933, N15932, N15931, N15930, N15929, N15928, N15927, N15926, N15925, N15924, N15923, N15922, N15921, N15920, N15919, N15918, N15917, N15916, N15915, N15914, N15913, N15912, N15911, N15910, N15909, N15908, N15907, N15906, N15905, N13058, N13057, N13056, N13055, N13054, N13053, N13052, N13051, N13050, N13049, N13048, N13047, N13046, N13045, N13044, N13043, N13042, N13041, N13040, N13039, N13038, N13037, N13036, N13035, N13034, N13033, N13032, N13031, N13030, N13029, N13028, N13027, N13026, N13025, N13024, N13023, N13022, N13021, N13020, N13019, N13018, N13017, N13016, N13015, N13014, N13013, N13012, N13011, N13010, N13009, N13008, N13007, N13006, N13005, N13004, N13003, N13002, N13001, N13000, N12999, N12998, N12997, N12996, N12995, N12479, N12478, N12477, N12476, N12475, N12474, N12473, N12472, N12471, N12470, N12469, N12468, N12467, N12466, N12465, N12464, N12463, N12462, N12461, N12460, N12459, N12458, N12457, N12456, N12455, N12454, N12453, N12452, N12451, N12450, N12449, N12448, N12447, N12446, N12445, N12444, N12443, N12442, N12441, N12440, N12439, N12438, N12437, N12436, N12435, N12434, N12433, N12432, N12431, N12430, N12429, N12428, N12427, N12426, N12425, N12424, N12423, N12422, N12421, N12420, N12419, N12418, N12417, N12416, N12143, N15904, N15903, N15902, N15901, N15900, N15899, N15898, N15897, N15896, N15895, N15894, N15893, N15892, N15891, N15890, N15889, N15888, N15887, N15886, N15885, N15884, N15883, N15882, N15881, N15880, N15879, N15878, N15877, N15876, N15875, N15874, N15873, N15872, N15871, N15870, N15869, N15868, N15867, N15866, N15865, N15864, N15863, N15862, N15861, N15860, N15859, N15858, N15857, N15856, N15855, N15854, N15853, N15852, N15851, N15850, N15849, N15848, N15847, N15846, N15845, N15844, N15843, N15842, N15841, N15840, N15839, N15838, N15837, N15836, N15835, N15834, N15833, N15832, N15831, N15830, N15829, N15828, N15827, N15826, N15825, N15824, N15823, N15822, N15821, N15820, N15819, N15818, N15817, N15816, N15815, N15814, N15813, N15812, N15811, N15810, N15809, N15808, N15807, N15806, N15805, N15804, N15803, N15802, N15801, N15800, N15799, N15798, N15797, N15796, N15795, N15794, N15793, N15792, N15791, N15790, N15789, N15788, N15787, N15786, N15785, N15784, N15783, N15782, N15781, N15780, N15779, N15778, N15777, N15776, N12994, N12993, N12992, N12991, N12990, N12989, N12988, N12987, N12986, N12985, N12984, N12983, N12982, N12981, N12980, N12979, N12978, N12977, N12976, N12975, N12974, N12973, N12972, N12971, N12970, N12969, N12968, N12967, N12966, N12965, N12964, N12963, N12962, N12961, N12960, N12959, N12958, N12957, N12956, N12955, N12954, N12953, N12952, N12951, N12950, N12949, N12948, N12947, N12946, N12945, N12944, N12943, N12942, N12941, N12940, N12939, N12938, N12937, N12936, N12935, N12934, N12933, N12932, N12931, N12414, N12413, N12412, N12411, N12410, N12409, N12408, N12407, N12406, N12405, N12404, N12403, N12402, N12401, N12400, N12399, N12398, N12397, N12396, N12395, N12394, N12393, N12392, N12391, N12390, N12389, N12388, N12387, N12386, N12385, N12384, N12383, N12382, N12381, N12380, N12379, N12378, N12377, N12376, N12375, N12374, N12373, N12372, N12371, N12370, N12369, N12368, N12367, N12366, N12365, N12364, N12363, N12362, N12361, N12360, N12359, N12358, N12357, N12356, N12355, N12354, N12353, N12352, N12351, N12142, N15775, N15774, N15773, N15772, N15771, N15770, N15769, N15768, N15767, N15766, N15765, N15764, N15763, N15762, N15761, N15760, N15759, N15758, N15757, N15756, N15755, N15754, N15753, N15752, N15751, N15750, N15749, N15748, N15747, N15746, N15745, N15744, N15743, N15742, N15741, N15740, N15739, N15738, N15737, N15736, N15735, N15734, N15733, N15732, N15731, N15730, N15729, N15728, N15727, N15726, N15725, N15724, N15723, N15722, N15721, N15720, N15719, N15718, N15717, N15716, N15715, N15714, N15713, N15712, N15711, N15710, N15709, N15708, N15707, N15706, N15705, N15704, N15703, N15702, N15701, N15700, N15699, N15698, N15697, N15696, N15695, N15694, N15693, N15692, N15691, N15690, N15689, N15688, N15687, N15686, N15685, N15684, N15683, N15682, N15681, N15680, N15679, N15678, N15677, N15676, N15675, N15674, N15673, N15672, N15671, N15670, N15669, N15668, N15667, N15666, N15665, N15664, N15663, N15662, N15661, N15660, N15659, N15658, N15657, N15656, N15655, N15654, N15653, N15652, N15651, N15650, N15649, N15648, N15647, N12930, N12929, N12928, N12927, N12926, N12925, N12924, N12923, N12922, N12921, N12920, N12919, N12918, N12917, N12916, N12915, N12914, N12913, N12912, N12911, N12910, N12909, N12908, N12907, N12906, N12905, N12904, N12903, N12902, N12901, N12900, N12899, N12898, N12897, N12896, N12895, N12894, N12893, N12892, N12891, N12890, N12889, N12888, N12887, N12886, N12885, N12884, N12883, N12882, N12881, N12880, N12879, N12878, N12877, N12876, N12875, N12874, N12873, N12872, N12871, N12870, N12869, N12868, N12867, N12349, N12348, N12347, N12346, N12345, N12344, N12343, N12342, N12341, N12340, N12339, N12338, N12337, N12336, N12335, N12334, N12333, N12332, N12331, N12330, N12329, N12328, N12327, N12326, N12325, N12324, N12323, N12322, N12321, N12320, N12319, N12318, N12317, N12316, N12315, N12314, N12313, N12312, N12311, N12310, N12309, N12308, N12307, N12306, N12305, N12304, N12303, N12302, N12301, N12300, N12299, N12298, N12297, N12296, N12295, N12294, N12293, N12292, N12291, N12290, N12289, N12288, N12287, N12286, N12141, N15646, N15645, N15644, N15643, N15642, N15641, N15640, N15639, N15638, N15637, N15636, N15635, N15634, N15633, N15632, N15631, N15630, N15629, N15628, N15627, N15626, N15625, N15624, N15623, N15622, N15621, N15620, N15619, N15618, N15617, N15616, N15615, N15614, N15613, N15612, N15611, N15610, N15609, N15608, N15607, N15606, N15605, N15604, N15603, N15602, N15601, N15600, N15599, N15598, N15597, N15596, N15595, N15594, N15593, N15592, N15591, N15590, N15589, N15588, N15587, N15586, N15585, N15584, N15583, N15582, N15581, N15580, N15579, N15578, N15577, N15576, N15575, N15574, N15573, N15572, N15571, N15570, N15569, N15568, N15567, N15566, N15565, N15564, N15563, N15562, N15561, N15560, N15559, N15558, N15557, N15556, N15555, N15554, N15553, N15552, N15551, N15550, N15549, N15548, N15547, N15546, N15545, N15544, N15543, N15542, N15541, N15540, N15539, N15538, N15537, N15536, N15535, N15534, N15533, N15532, N15531, N15530, N15529, N15528, N15527, N15526, N15525, N15524, N15523, N15522, N15521, N15520, N15519, N15518, N12866, N12865, N12864, N12863, N12862, N12861, N12860, N12859, N12858, N12857, N12856, N12855, N12854, N12853, N12852, N12851, N12850, N12849, N12848, N12847, N12846, N12845, N12844, N12843, N12842, N12841, N12840, N12839, N12838, N12837, N12836, N12835, N12834, N12833, N12832, N12831, N12830, N12829, N12828, N12827, N12826, N12825, N12824, N12823, N12822, N12821, N12820, N12819, N12818, N12817, N12816, N12815, N12814, N12813, N12812, N12811, N12810, N12809, N12808, N12807, N12806, N12805, N12804, N12803, N12284, N12283, N12282, N12281, N12280, N12279, N12278, N12277, N12276, N12275, N12274, N12273, N12272, N12271, N12270, N12269, N12268, N12267, N12266, N12265, N12264, N12263, N12262, N12261, N12260, N12259, N12258, N12257, N12256, N12255, N12254, N12253, N12252, N12251, N12250, N12249, N12248, N12247, N12246, N12245, N12244, N12243, N12242, N12241, N12240, N12239, N12238, N12237, N12236, N12235, N12234, N12233, N12232, N12231, N12230, N12229, N12228, N12227, N12226, N12225, N12224, N12223, N12222, N12221, N12140, N15517, N15516, N15515, N15514, N15513, N15512, N15511, N15510, N15509, N15508, N15507, N15506, N15505, N15504, N15503, N15502, N15501, N15500, N15499, N15498, N15497, N15496, N15495, N15494, N15493, N15492, N15491, N15490, N15489, N15488, N15487, N15486, N15485, N15484, N15483, N15482, N15481, N15480, N15479, N15478, N15477, N15476, N15475, N15474, N15473, N15472, N15471, N15470, N15469, N15468, N15467, N15466, N15465, N15464, N15463, N15462, N15461, N15460, N15459, N15458, N15457, N15456, N15455, N15454, N15453, N15452, N15451, N15450, N15449, N15448, N15447, N15446, N15445, N15444, N15443, N15442, N15441, N15440, N15439, N15438, N15437, N15436, N15435, N15434, N15433, N15432, N15431, N15430, N15429, N15428, N15427, N15426, N15425, N15424, N15423, N15422, N15421, N15420, N15419, N15418, N15417, N15416, N15415, N15414, N15413, N15412, N15411, N15410, N15409, N15408, N15407, N15406, N15405, N15404, N15403, N15402, N15401, N15400, N15399, N15398, N15397, N15396, N15395, N15394, N15393, N15392, N15391, N15390, N15389, N12802, N12801, N12800, N12799, N12798, N12797, N12796, N12795, N12794, N12793, N12792, N12791, N12790, N12789, N12788, N12787, N12786, N12785, N12784, N12783, N12782, N12781, N12780, N12779, N12778, N12777, N12776, N12775, N12774, N12773, N12772, N12771, N12770, N12769, N12768, N12767, N12766, N12765, N12764, N12763, N12762, N12761, N12760, N12759, N12758, N12757, N12756, N12755, N12754, N12753, N12752, N12751, N12750, N12749, N12748, N12747, N12746, N12745, N12744, N12743, N12742, N12741, N12740, N12739, N12219, N12218, N12217, N12216, N12215, N12214, N12213, N12212, N12211, N12210, N12209, N12208, N12207, N12206, N12205, N12204, N12203, N12202, N12201, N12200, N12199, N12198, N12197, N12196, N12195, N12194, N12193, N12192, N12191, N12190, N12189, N12188, N12187, N12186, N12185, N12184, N12183, N12182, N12181, N12180, N12179, N12178, N12177, N12176, N12175, N12174, N12173, N12172, N12171, N12170, N12169, N12168, N12167, N12166, N12165, N12164, N12163, N12162, N12161, N12160, N12159, N12158, N12157, N12156, N12139, N15388, N15387, N15386, N15385, N15384, N15383, N15382, N15381, N15380, N15379, N15378, N15377, N15376, N15375, N15374, N15373, N15372, N15371, N15370, N15369, N15368, N15367, N15366, N15365, N15364, N15363, N15362, N15361, N15360, N15359, N15358, N15357, N15356, N15355, N15354, N15353, N15352, N15351, N15350, N15349, N15348, N15347, N15346, N15345, N15344, N15343, N15342, N15341, N15340, N15339, N15338, N15337, N15336, N15335, N15334, N15333, N15332, N15331, N15330, N15329, N15328, N15327, N15326, N15325, N15324, N15323, N15322, N15321, N15320, N15319, N15318, N15317, N15316, N15315, N15314, N15313, N15312, N15311, N15310, N15309, N15308, N15307, N15306, N15305, N15304, N15303, N15302, N15301, N15300, N15299, N15298, N15297, N15296, N15295, N15294, N15293, N15292, N15291, N15290, N15289, N15288, N15287, N15286, N15285, N15284, N15283, N15282, N15281, N15280, N15279, N15278, N15277, N15276, N15275, N15274, N15273, N15272, N15271, N15270, N15269, N15268, N15267, N15266, N15265, N15264, N15263, N15262, N15261, N15260, N12738, N12737, N12736, N12735, N12734, N12733, N12732, N12731, N12730, N12729, N12728, N12727, N12726, N12725, N12724, N12723, N12722, N12721, N12720, N12719, N12718, N12717, N12716, N12715, N12714, N12713, N12712, N12711, N12710, N12709, N12708, N12707, N12706, N12705, N12704, N12703, N12702, N12701, N12700, N12699, N12698, N12697, N12696, N12695, N12694, N12693, N12692, N12691, N12690, N12689, N12688, N12687, N12686, N12685, N12684, N12683, N12682, N12681, N12680, N12679, N12678, N12677, N12676, N12675 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12138)? { N12120, N12119, N12118, N12117, N12116, N12115, N12114, N12113, N12112, N12111, N12110, N12109, N12108, N12107, N12106, N12105, N12104, N12103, N12102, N12101, N12100, N12099, N12098, N12097, N12096, N12095, N12094, N12093, N12092, N12091, N12090, N12089, N12088, N12087, N12086, N12085, N12084, N12083, N12082, N12081, N12080, N12079, N12078, N12077, N12076, N12075, N12074, N12073, N12072, N12071, N12070, N12069, N12068, N12067, N12066, N12065, N12064, N12063, N12062, N12061, N12060, N12059, N12058, N12057, N12056, N12055, N12054, N12053, N12052, N12051, N12050, N12049, N12048, N12047, N12046, N12045, N12044, N12043, N12042, N12041, N12040, N12039, N12038, N12037, N12036, N12035, N12034, N12033, N12032, N12031, N12030, N12029, N12028, N12027, N12026, N12025, N12024, N12023, N12022, N12021, N12020, N12019, N12018, N12017, N12016, N12015, N12014, N12013, N12012, N12011, N12010, N12009, N12008, N12007, N12006, N12005, N12004, N12003, N12002, N12001, N12000, N11999, N11998, N11997, N11996, N11995, N11994, N11993, N11992, N11991, N11990, N11989, N11988, N11987, N11986, N11985, N11984, N11983, N11982, N11981, N11980, N11979, N11978, N11977, N11976, N11975, N11974, N11973, N11972, N11971, N11970, N11969, N11968, N11967, N11966, N11965, N11964, N11963, N11962, N11961, N11960, N11959, N11958, N11957, N11956, N11955, N11954, N11953, N11952, N11951, N11950, N11949, N11948, N11947, N11946, N11945, N11944, N11943, N11942, N11941, N11940, N11939, N11938, N11937, N11936, N11935, N11934, N11933, N11932, N11931, N11930, N11929, N11928, N11927, N11926, N11925, N11924, N11923, N11922, N11921, N11920, N11919, N11918, N11917, N11916, N11915, N11914, N11913, N11912, N11911, N11910, N11909, N11908, N11907, N11906, N11905, N11904, N11903, N11902, N11901, N11900, N11899, N11898, N11897, N11896, N11895, N11894, N11893, N11892, N11891, N11890, N11889, N11888, N11887, N11886, N11885, N11884, N11883, N11882, N11881, N11880, N11879, N11878, N11877, N11876, N11875, N11874, N11873, N11872, N11871, N11870, N11869, N11868, N11867, N11866, N11865, N11864, N11863, N11862, N11861, N11860, N11859, N11858, N11857, N11856, N11855, N11854, N11853, N11852, N11851, N11850, N11849, N11848, N11847, N11846, N11845, N11844, N11843, N11842, N11841, N11840, N11839, N11838, N11837, N11836, N11835, N11834, N11833, N11832, N11831, N11830, N11829, N11828, N11827, N11826, N11825, N11824, N11823, N11822, N11821, N11820, N11819, N11818, N11817, N11816, N11815, N11814, N11813, N11812, N11811, N11810, N11809, N11808, N11807, N11806, N11805, N11804, N11803, N11802, N11801, N11800, N11799, N11798, N11797, N11796, N11795, N11794, N11793, N11792, N11791, N11790, N11789, N11788, N11787, N11786, N11785, N11784, N11783, N11782, N11781, N11780, N11779, N11778, N11777, N11776, N11775, N11774, N11773, N11772, N11771, N11770, N11769, N11768, N11767, N11766, N11765, N11764, N11763, N11762, N11761, N11760, N11759, N11758, N11757, N11756, N11755, N11754, N11753, N11752, N11751, N11750, N11749, N11748, N11747, N11746, N11745, N11744, N11743, N11742, N11741, N11740, N11739, N11738, N11737, N11736, N11735, N11734, N11733, N11732, N11731, N11730, N11729, N11728, N11727, N11726, N11725, N11724, N11723, N11722, N11721, N11720, N11719, N11718, N11717, N11716, N11715, N11714, N11713, N11712, N11711, N11710, N11709, N11708, N11707, N11706, N11705, N11704, N11703, N11702, N11701, N11700, N11699, N11698, N11697, N11696, N11695, N11694, N11693, N11692, N11691, N11690, N11689, N11688, N11687, N11686, N11685, N11684, N11683, N11682, N11681, N11680, N11679, N11678, N11677, N11676, N11675, N11674, N11673, N11672, N11671, N11670, N11669, N11668, N11667, N11666, N11665, N11664, N11663, N11662, N11661, N11660, N11659, N11658, N11657, N11656, N11655, N11654, N11653, N11652, N11651, N11650, N11649, N11648, N11647, N11646, N11645, N11644, N11643, N11642, N11641, N11640, N11639, N11638, N11637, N11636, N11635, N11634, N11633, N11632, N11631, N11630, N11629, N11628, N11627, N11626, N11625, N11624, N11623, N11622, N11621, N11620, N11619, N11618, N11617, N11616, N11615, N11614, N11613, N11612, N11611, N11610, N11609, N11608, N11607, N11606, N11605, N11604, N11603, N11602, N11601, N11600, N11599, N11598, N11597, N11596, N11595, N11594, N11593, N11592, N11591, N11590, N11589, N11588, N11587, N11586, N11585, N11584, N11583, N11582, N11581, N11580, N11579, N11578, N11577, N11576, N11575, N11574, N11573, N11572, N11571, N11570, N11569, N11568, N11567, N11566, N11565, N11564, N11563, N11562, N11561, N11560, N11559, N11558, N11557, N11556, N11555, N11554, N11553, N11552, N11551, N11550, N11549, N11548, N11547, N11546, N11545, N11544, N11543, N11542, N11541, N11540, N11539, N11538, N11537, N11536, N11535, N11534, N11533, N11532, N11531, N11530, N11529, N11528, N11527, N11526, N11525, N11524, N11523, N11522, N11521, N11520, N11519, N11518, N11517, N11516, N11515, N11514, N11513, N11512, N11511, N11510, N11509, N11508, N11507, N11506, N11505, N11504, N11503, N11502, N11501, N11500, N11499, N11498, N11497, N11496, N11495, N11494, N11493, N11492, N11491, N11490, N11489, N11488, N11487, N11486, N11485, N11484, N11483, N11482, N11481, N11480, N11479, N11478, N11477, N11476, N11475, N11474, N11473, N11472, N11471, N11470, N11469, N11468, N11467, N11466, N11465, N11464, N11463, N11462, N11461, N11460, N11459, N11458, N11457, N11456, N11455, N11454, N11453, N11452, N11451, N11450, N11449, N11448, N11447, N11446, N11445, N11444, N11443, N11442, N11441, N11440, N11439, N11438, N11437, N11436, N11435, N11434, N11433, N11432, N11431, N11430, N11429, N11428, N11427, N11426, N11425, N11424, N11423, N11422, N11421, N11420, N11419, N11418, N11417, N11416, N11415, N11414, N11413, N11412, N11411, N11410, N11409, N11408, N11407, N11406, N11405, N11404, N11403, N11402, N11401, N11400, N11399, N11398, N11397, N11396, N11395, N11394, N11393, N11392, N11391, N11390, N11389, N11388, N11387, N11386, N11385, N11384, N11383, N11382, N11381, N11380, N11379, N11378, N11377, N11376, N11375, N11374, N11373, N11372, N11371, N11370, N11369, N11368, N11367, N11366, N11365, N11364, N11363, N11362, N11361, N11360, N11359, N11358, N11357, N11356, N11355, N11354, N11353, N11352, N11351, N11350, N11349, N11348, N11347, N11346, N11345, N11344, N11343, N11342, N11341, N11340, N11339, N11338, N11337, N11336, N11335, N11334, N11333, N11332, N11331, N11330, N11329, N11328, N11327, N11326, N11325, N11324, N11323, N11322, N11321, N11320, N11319, N11318, N11317, N11316, N11315, N11314, N11313, N11312, N11311, N11310, N11309, N11308, N11307, N11306, N11305, N11304, N11303, N11302, N11301, N11300, N11299, N11298, N11297, N11296, N11295, N11294, N11293, N11292, N11291, N11290, N11289, N11288, N11287, N11286, N11285, N11284, N11283, N11282, N11281, N11280, N11279, N11278, N11277, N11276, N11275, N11274, N11273, N11272, N11271, N11270, N11269, N11268, N11267, N11266, N11265, N11264, N11263, N11262, N11261, N11260, N11259, N11258, N11257, N11256, N11255, N11254, N11253, N11252, N11251, N11250, N11249, N11248, N11247, N11246, N11245, N11244, N11243, N11242, N11241, N11240, N11239, N11238, N11237, N11236, N11235, N11234, N11233, N11232, N11231, N11230, N11229, N11228, N11227, N11226, N11225, N11224, N11223, N11222, N11221, N11220, N11219, N11218, N11217, N11216, N11215, N11214, N11213, N11212, N11211, N11210, N11209, N11208, N11207, N11206, N11205, N11204, N11203, N11202, N11201, N11200, N11199, N11198, N11197, N11196, N11195, N11194, N11193, N11192, N11191, N11190, N11189, N11188, N11187, N11186, N11185, N11184, N11183, N11182, N11181, N11180, N11179, N11178, N11177, N11176, N11175, N11174, N11173, N11172, N11171, N11170, N11169, N11168, N11167, N11166, N11165, N11164, N11163, N11162, N11161, N11160, N11159, N11158, N11157, N11156, N11155, N11154, N11153, N11152, N11151, N11150, N11149, N11148, N11147, N11146, N11145, N11144, N11143, N11142, N11141, N11140, N11139, N11138, N11137, N11136, N11135, N11134, N11133, N11132, N11131, N11130, N11129, N11128, N11127, N11126, N11125, N11124, N11123, N11122, N11121, N11120, N11119, N11118, N11117, N11116, N11115, N11114, N11113, N11112, N11111, N11110, N11109, N11108, N11107, N11106, N11105, N11104, N11103, N11102, N11101, N11100, N11099, N11098, N11097, N11096, N11095, N11094, N11093, N11092, N11091, N11090, N11089, N11088, N11087, N11086, N11085, N11084, N11083, N11082, N11081, N11080, N11079, N11078, N11077, N11076, N11075, N11074, N11073, N11072, N11071, N11070, N11069, N11068, N11067, N11066, N11065, N11064, N11063, N11062, N11061, N11060, N11059, N11058, N11057, N11056, N11055, N11054, N11053, N11052, N11051, N11050, N11049, N11048, N11047, N11046, N11045, N11044, N11043, N11042, N11041, N11040, N11039, N11038, N11037, N11036, N11035, N11034, N11033, N11032, N11031, N11030, N11029, N11028, N11027, N11026, N11025, N11024, N11023, N11022, N11021, N11020, N11019, N11018, N11017, N11016, N11015, N11014, N11013, N11012, N11011, N11010, N11009, N11008, N11007, N11006, N11005, N11004, N11003, N11002, N11001, N11000, N10999, N10998, N10997, N10996, N10995, N10994, N10993, N10992, N10991, N10990, N10989, N10988, N10987, N10986, N10985, N10984, N10983, N10982, N10981, N10980, N10979, N10978, N10977, N10976, N10975, N10974, N10973, N10972, N10971, N10970, N10969, N10968, N10967, N10966, N10965, N10964, N10963, N10962, N10961, N10960, N10959, N10958, N10957, N10956, N10955, N10954, N10953, N10952, N10951, N10950, N10949, N10948, N10947, N10946, N10945, N10944, N10943, N10942, N10941, N10940, N10939, N10938, N10937, N10936, N10935, N10934, N10933, N10932, N10931, N10930, N10929, N10928, N10927, N10926, N10925, N10924, N10923, N10922, N10921, N10920, N10919, N10918, N10917, N10916, N10915, N10914, N10913, N10912, N10911, N10910, N10909, N10908, N10907, N10906, N10905, N10904, N10903, N10902, N10901, N10900, N10899, N10898, N10897, N10896, N10895, N10894, N10893, N10892, N10891, N10890, N10889, N10888, N10887, N10886, N10885, N10884, N10883, N10882, N10881, N10880, N10879, N10878, N10877, N10876, N10875, N10874, N10873, N10872, N10871, N10870, N10869, N10868, N10867, N10866, N10865, N10864, N10863, N10862, N10861, N10860, N10859, N10858, N10857, N10856, N10855, N10854, N10853, N10852, N10851, N10850, N10849, N10848, N10847, N10846, N10845, N10844, N10843, N10842, N10841, N10840, N10839, N10838, N10837, N10836, N10835, N10834, N10833, N10832, N10831, N10830, N10829, N10828, N10827, N10826, N10825, N10824, N10823, N10822, N10821, N10820, N10819, N10818, N10817, N10816, N10815, N10814, N10813, N10812, N10811, N10810, N10809, N10808, N10807, N10806, N10805, N10804, N10803, N10802, N10801, N10800, N10799, N10798, N10797, N10796, N10795, N10794, N10793, N10792, N10791, N10790, N10789, N10788, N10787, N10786, N10785, N10784, N10783, N10782, N10781, N10780, N10779, N10778, N10777, N10776, N10775, N10774, N10773, N10772, N10771, N10770, N10769, N10768, N10767, N10766, N10765, N10764, N10763, N10762, N10761, N10760, N10759, N10758, N10757, N10756, N10755, N10754, N10753, N10752, N10751, N10750, N10749, N10748, N10747, N10746, N10745, N10744, N10743, N10742, N10741, N10740, N10739, N10738, N10737, N10736, N10735, N10734, N10733, N10732, N10731, N10730, N10729, N10728, N10727, N10726, N10725, N10724, N10723, N10722, N10721, N10720, N10719, N10718, N10717, N10716, N10715, N10714, N10713, N10712, N10711, N10710, N10709, N10708, N10707, N10706, N10705, N10704, N10703, N10702, N10701, N10700, N10699, N10698, N10697, N10696, N10695, N10694, N10693, N10692, N10691, N10690, N10689, N10688, N10687, N10686, N10685, N10684, N10683, N10682, N10681, N10680, N10679, N10678, N10677, N10676, N10675, N10674, N10673, N10672, N10671, N10670, N10669, N10668, N10667, N10666, N10665, N10664, N10663, N10662, N10661, N10660, N10659, N10658, N10657, N10656, N10655, N10654, N10653, N10652, N10651, N10650, N10649, N10648, N10647, N10646, N10645, N10644, N10643, N10642, N10641, N10640, N10639, N10638, N10637, N10636, N10635, N10634, N10633, N10632, N10631, N10630, N10629, N10628, N10627, N10626, N10625, N10624, N10623, N10622, N10621, N10620, N10619, N10618, N10617, N10616, N10615, N10614, N10613, N10612, N10611, N10610, N10609, N10608, N10607, N10606, N10605, N10604, N10603, N10602, N10601, N10600, N10599, N10598, N10597, N10596, N10595, N10594, N10593, N10592, N10591, N10590, N10589, N10588, N10587, N10586, N10585, N10584, N10583, N10582, N10581, N10580, N10579, N10578, N10577, N10576, N10575, N10574, N10573, N10572, N10571, N10570, N10569, N10568, N10567, N10566, N10565, N10564, N10563, N10562, N10561, N10560, N10559, N10558, N10557, N10556, N10555, N10554, N10553, N10552, N10551, N10550, N10549, N10548, N10547, N10546, N10545, N10544, N10543, N10542, N10541, N10540, N10539, N10538, N10537, N10536, N10535, N10534, N10533, N10532, N10531, N10530, N10529, N10528, N10527, N10526, N10525, N10524, N10523, N10522, N10521, N10520, N10519, N10518, N10517, N10516, N10515, N10514, N10513, N10512, N10511, N10510, N10509, N10508, N10507, N10506, N10505, N10504, N10503, N10502, N10501, N10500, N10499, N10498, N10497, N10496, N10495, N10494, N10493, N10492, N10491, N10490, N10489, N10488, N10487, N10486, N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422, N10421, N10420, N10419, N10418, N10417, N10416, N10415, N10414, N10413, N10412, N10411, N10410, N10409, N10408, N10407, N10406, N10405, N10404, N10403, N10402, N10401, N10400, N10399, N10398, N10397, N10396, N10395, N10394, N10393, N10392, N10391, N10390, N10389, N10388, N10387, N10386, N10385, N10384, N10383, N10382, N10381, N10380, N10379, N10378, N10377, N10376, N10375, N10374, N10373, N10372, N10371, N10370, N10369, N10368, N10367, N10366, N10365, N10364, N10363, N10362, N10361, N10360, N10359, N10358, N10357, N10356, N10355, N10354, N10353, N10352, N10351, N10350, N10349, N10348, N10347, N10346, N10345, N10344, N10343, N10342, N10341, N10340, N10339, N10338, N10337, N10336, N10335, N10334, N10333, N10332, N10331, N10330, N10329, N10328, N10327, N10326, N10325, N10324, N10323, N10322, N10321, N10320, N10319, N10318, N10317, N10316, N10315, N10314, N10313, N10312, N10311, N10310, N10309, N10308, N10307, N10306, N10305, N10304, N10303, N10302, N10301, N10300, N10299, N10298, N10297, N10296, N10295, N10294, N10293, N10292, N10291, N10290, N10289, N10288, N10287, N10286, N10285, N10284, N10283, N10282, N10281, N10280, N10279, N10278, N10277, N10276, N10275, N10274, N10273, N10272, N10271, N10270, N10269, N10268, N10267, N10266, N10265, N10264, N10263, N10262, N10261, N10260, N10259, N10258, N10257, N10256, N10255, N10254, N10253, N10252, N10251, N10250, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057 } : 1'b0;
  assign N180 = N12137;
  assign N18374 = (N181)? 1'b1 : 
                  (N18390)? N16485 : 1'b0;
  assign N181 = N18382;
  assign N18375 = (N182)? 1'b1 : 
                  (N18455)? N16743 : 1'b0;
  assign N182 = N18383;
  assign N18376 = (N183)? 1'b1 : 
                  (N18520)? N17001 : 1'b0;
  assign N183 = N18384;
  assign N18377 = (N184)? 1'b1 : 
                  (N18585)? N17259 : 1'b0;
  assign N184 = N18385;
  assign N18378 = (N185)? 1'b1 : 
                  (N18650)? N17517 : 1'b0;
  assign N185 = N18386;
  assign N18379 = (N186)? 1'b1 : 
                  (N18715)? N17775 : 1'b0;
  assign N186 = N18387;
  assign N18380 = (N187)? 1'b1 : 
                  (N18780)? N18033 : 1'b0;
  assign N187 = N18388;
  assign N18381 = (N188)? 1'b1 : 
                  (N18845)? N18291 : 1'b0;
  assign N188 = N18389;
  assign { N18454, N18453, N18452, N18451, N18450, N18449, N18448, N18447, N18446, N18445, N18444, N18443, N18442, N18441, N18440, N18439, N18438, N18437, N18436, N18435, N18434, N18433, N18432, N18431, N18430, N18429, N18428, N18427, N18426, N18425, N18424, N18423, N18422, N18421, N18420, N18419, N18418, N18417, N18416, N18415, N18414, N18413, N18412, N18411, N18410, N18409, N18408, N18407, N18406, N18405, N18404, N18403, N18402, N18401, N18400, N18399, N18398, N18397, N18396, N18395, N18394, N18393, N18392, N18391 } = (N181)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18390)? { N16549, N16548, N16547, N16546, N16545, N16544, N16543, N16542, N16541, N16540, N16539, N16538, N16537, N16536, N16535, N16534, N16533, N16532, N16531, N16530, N16529, N16528, N16527, N16526, N16525, N16524, N16523, N16522, N16521, N16520, N16519, N16518, N16517, N16516, N16515, N16514, N16513, N16512, N16511, N16510, N16509, N16508, N16507, N16506, N16505, N16504, N16503, N16502, N16501, N16500, N16499, N16498, N16497, N16496, N16495, N16494, N16493, N16492, N16491, N16490, N16489, N16488, N16487, N16486 } : 1'b0;
  assign { N18519, N18518, N18517, N18516, N18515, N18514, N18513, N18512, N18511, N18510, N18509, N18508, N18507, N18506, N18505, N18504, N18503, N18502, N18501, N18500, N18499, N18498, N18497, N18496, N18495, N18494, N18493, N18492, N18491, N18490, N18489, N18488, N18487, N18486, N18485, N18484, N18483, N18482, N18481, N18480, N18479, N18478, N18477, N18476, N18475, N18474, N18473, N18472, N18471, N18470, N18469, N18468, N18467, N18466, N18465, N18464, N18463, N18462, N18461, N18460, N18459, N18458, N18457, N18456 } = (N182)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18455)? { N16807, N16806, N16805, N16804, N16803, N16802, N16801, N16800, N16799, N16798, N16797, N16796, N16795, N16794, N16793, N16792, N16791, N16790, N16789, N16788, N16787, N16786, N16785, N16784, N16783, N16782, N16781, N16780, N16779, N16778, N16777, N16776, N16775, N16774, N16773, N16772, N16771, N16770, N16769, N16768, N16767, N16766, N16765, N16764, N16763, N16762, N16761, N16760, N16759, N16758, N16757, N16756, N16755, N16754, N16753, N16752, N16751, N16750, N16749, N16748, N16747, N16746, N16745, N16744 } : 1'b0;
  assign { N18584, N18583, N18582, N18581, N18580, N18579, N18578, N18577, N18576, N18575, N18574, N18573, N18572, N18571, N18570, N18569, N18568, N18567, N18566, N18565, N18564, N18563, N18562, N18561, N18560, N18559, N18558, N18557, N18556, N18555, N18554, N18553, N18552, N18551, N18550, N18549, N18548, N18547, N18546, N18545, N18544, N18543, N18542, N18541, N18540, N18539, N18538, N18537, N18536, N18535, N18534, N18533, N18532, N18531, N18530, N18529, N18528, N18527, N18526, N18525, N18524, N18523, N18522, N18521 } = (N183)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18520)? { N17065, N17064, N17063, N17062, N17061, N17060, N17059, N17058, N17057, N17056, N17055, N17054, N17053, N17052, N17051, N17050, N17049, N17048, N17047, N17046, N17045, N17044, N17043, N17042, N17041, N17040, N17039, N17038, N17037, N17036, N17035, N17034, N17033, N17032, N17031, N17030, N17029, N17028, N17027, N17026, N17025, N17024, N17023, N17022, N17021, N17020, N17019, N17018, N17017, N17016, N17015, N17014, N17013, N17012, N17011, N17010, N17009, N17008, N17007, N17006, N17005, N17004, N17003, N17002 } : 1'b0;
  assign { N18649, N18648, N18647, N18646, N18645, N18644, N18643, N18642, N18641, N18640, N18639, N18638, N18637, N18636, N18635, N18634, N18633, N18632, N18631, N18630, N18629, N18628, N18627, N18626, N18625, N18624, N18623, N18622, N18621, N18620, N18619, N18618, N18617, N18616, N18615, N18614, N18613, N18612, N18611, N18610, N18609, N18608, N18607, N18606, N18605, N18604, N18603, N18602, N18601, N18600, N18599, N18598, N18597, N18596, N18595, N18594, N18593, N18592, N18591, N18590, N18589, N18588, N18587, N18586 } = (N184)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18585)? { N17323, N17322, N17321, N17320, N17319, N17318, N17317, N17316, N17315, N17314, N17313, N17312, N17311, N17310, N17309, N17308, N17307, N17306, N17305, N17304, N17303, N17302, N17301, N17300, N17299, N17298, N17297, N17296, N17295, N17294, N17293, N17292, N17291, N17290, N17289, N17288, N17287, N17286, N17285, N17284, N17283, N17282, N17281, N17280, N17279, N17278, N17277, N17276, N17275, N17274, N17273, N17272, N17271, N17270, N17269, N17268, N17267, N17266, N17265, N17264, N17263, N17262, N17261, N17260 } : 1'b0;
  assign { N18714, N18713, N18712, N18711, N18710, N18709, N18708, N18707, N18706, N18705, N18704, N18703, N18702, N18701, N18700, N18699, N18698, N18697, N18696, N18695, N18694, N18693, N18692, N18691, N18690, N18689, N18688, N18687, N18686, N18685, N18684, N18683, N18682, N18681, N18680, N18679, N18678, N18677, N18676, N18675, N18674, N18673, N18672, N18671, N18670, N18669, N18668, N18667, N18666, N18665, N18664, N18663, N18662, N18661, N18660, N18659, N18658, N18657, N18656, N18655, N18654, N18653, N18652, N18651 } = (N185)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18650)? { N17581, N17580, N17579, N17578, N17577, N17576, N17575, N17574, N17573, N17572, N17571, N17570, N17569, N17568, N17567, N17566, N17565, N17564, N17563, N17562, N17561, N17560, N17559, N17558, N17557, N17556, N17555, N17554, N17553, N17552, N17551, N17550, N17549, N17548, N17547, N17546, N17545, N17544, N17543, N17542, N17541, N17540, N17539, N17538, N17537, N17536, N17535, N17534, N17533, N17532, N17531, N17530, N17529, N17528, N17527, N17526, N17525, N17524, N17523, N17522, N17521, N17520, N17519, N17518 } : 1'b0;
  assign { N18779, N18778, N18777, N18776, N18775, N18774, N18773, N18772, N18771, N18770, N18769, N18768, N18767, N18766, N18765, N18764, N18763, N18762, N18761, N18760, N18759, N18758, N18757, N18756, N18755, N18754, N18753, N18752, N18751, N18750, N18749, N18748, N18747, N18746, N18745, N18744, N18743, N18742, N18741, N18740, N18739, N18738, N18737, N18736, N18735, N18734, N18733, N18732, N18731, N18730, N18729, N18728, N18727, N18726, N18725, N18724, N18723, N18722, N18721, N18720, N18719, N18718, N18717, N18716 } = (N186)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18715)? { N17839, N17838, N17837, N17836, N17835, N17834, N17833, N17832, N17831, N17830, N17829, N17828, N17827, N17826, N17825, N17824, N17823, N17822, N17821, N17820, N17819, N17818, N17817, N17816, N17815, N17814, N17813, N17812, N17811, N17810, N17809, N17808, N17807, N17806, N17805, N17804, N17803, N17802, N17801, N17800, N17799, N17798, N17797, N17796, N17795, N17794, N17793, N17792, N17791, N17790, N17789, N17788, N17787, N17786, N17785, N17784, N17783, N17782, N17781, N17780, N17779, N17778, N17777, N17776 } : 1'b0;
  assign { N18844, N18843, N18842, N18841, N18840, N18839, N18838, N18837, N18836, N18835, N18834, N18833, N18832, N18831, N18830, N18829, N18828, N18827, N18826, N18825, N18824, N18823, N18822, N18821, N18820, N18819, N18818, N18817, N18816, N18815, N18814, N18813, N18812, N18811, N18810, N18809, N18808, N18807, N18806, N18805, N18804, N18803, N18802, N18801, N18800, N18799, N18798, N18797, N18796, N18795, N18794, N18793, N18792, N18791, N18790, N18789, N18788, N18787, N18786, N18785, N18784, N18783, N18782, N18781 } = (N187)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18780)? { N18097, N18096, N18095, N18094, N18093, N18092, N18091, N18090, N18089, N18088, N18087, N18086, N18085, N18084, N18083, N18082, N18081, N18080, N18079, N18078, N18077, N18076, N18075, N18074, N18073, N18072, N18071, N18070, N18069, N18068, N18067, N18066, N18065, N18064, N18063, N18062, N18061, N18060, N18059, N18058, N18057, N18056, N18055, N18054, N18053, N18052, N18051, N18050, N18049, N18048, N18047, N18046, N18045, N18044, N18043, N18042, N18041, N18040, N18039, N18038, N18037, N18036, N18035, N18034 } : 1'b0;
  assign { N18909, N18908, N18907, N18906, N18905, N18904, N18903, N18902, N18901, N18900, N18899, N18898, N18897, N18896, N18895, N18894, N18893, N18892, N18891, N18890, N18889, N18888, N18887, N18886, N18885, N18884, N18883, N18882, N18881, N18880, N18879, N18878, N18877, N18876, N18875, N18874, N18873, N18872, N18871, N18870, N18869, N18868, N18867, N18866, N18865, N18864, N18863, N18862, N18861, N18860, N18859, N18858, N18857, N18856, N18855, N18854, N18853, N18852, N18851, N18850, N18849, N18848, N18847, N18846 } = (N188)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18845)? { N18355, N18354, N18353, N18352, N18351, N18350, N18349, N18348, N18347, N18346, N18345, N18344, N18343, N18342, N18341, N18340, N18339, N18338, N18337, N18336, N18335, N18334, N18333, N18332, N18331, N18330, N18329, N18328, N18327, N18326, N18325, N18324, N18323, N18322, N18321, N18320, N18319, N18318, N18317, N18316, N18315, N18314, N18313, N18312, N18311, N18310, N18309, N18308, N18307, N18306, N18305, N18304, N18303, N18302, N18301, N18300, N18299, N18298, N18297, N18296, N18295, N18294, N18293, N18292 } : 1'b0;
  assign { N18973, N18972, N18971, N18970, N18969, N18968, N18967, N18966, N18965, N18964, N18963, N18962, N18961, N18960, N18959, N18958, N18957, N18956, N18955, N18954, N18953, N18952, N18951, N18950, N18949, N18948, N18947, N18946, N18945, N18944, N18943, N18942, N18941, N18940, N18939, N18938, N18937, N18936, N18935, N18934, N18933, N18932, N18931, N18930, N18929, N18928, N18927, N18926, N18925, N18924, N18923, N18922, N18921, N18920, N18919, N18918, N18917, N18916, N18915, N18914, N18913, N18912, N18911, N18910 } = (N181)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18390)? { N16355, N16354, N16353, N16352, N16351, N16350, N16349, N16348, N16347, N16346, N16345, N16344, N16343, N16342, N16341, N16340, N16339, N16338, N16337, N16336, N16335, N16334, N16333, N16332, N16331, N16330, N16329, N16328, N16327, N16326, N16325, N16324, N16323, N16322, N16321, N16320, N16319, N16318, N16317, N16316, N16315, N16314, N16313, N16312, N16311, N16310, N16309, N16308, N16307, N16306, N16305, N16304, N16303, N16302, N16301, N16300, N16299, N16298, N16297, N16296, N16295, N16294, N16293, N16292 } : 1'b0;
  assign { N19037, N19036, N19035, N19034, N19033, N19032, N19031, N19030, N19029, N19028, N19027, N19026, N19025, N19024, N19023, N19022, N19021, N19020, N19019, N19018, N19017, N19016, N19015, N19014, N19013, N19012, N19011, N19010, N19009, N19008, N19007, N19006, N19005, N19004, N19003, N19002, N19001, N19000, N18999, N18998, N18997, N18996, N18995, N18994, N18993, N18992, N18991, N18990, N18989, N18988, N18987, N18986, N18985, N18984, N18983, N18982, N18981, N18980, N18979, N18978, N18977, N18976, N18975, N18974 } = (N182)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18455)? { N16613, N16612, N16611, N16610, N16609, N16608, N16607, N16606, N16605, N16604, N16603, N16602, N16601, N16600, N16599, N16598, N16597, N16596, N16595, N16594, N16593, N16592, N16591, N16590, N16589, N16588, N16587, N16586, N16585, N16584, N16583, N16582, N16581, N16580, N16579, N16578, N16577, N16576, N16575, N16574, N16573, N16572, N16571, N16570, N16569, N16568, N16567, N16566, N16565, N16564, N16563, N16562, N16561, N16560, N16559, N16558, N16557, N16556, N16555, N16554, N16553, N16552, N16551, N16550 } : 1'b0;
  assign { N19101, N19100, N19099, N19098, N19097, N19096, N19095, N19094, N19093, N19092, N19091, N19090, N19089, N19088, N19087, N19086, N19085, N19084, N19083, N19082, N19081, N19080, N19079, N19078, N19077, N19076, N19075, N19074, N19073, N19072, N19071, N19070, N19069, N19068, N19067, N19066, N19065, N19064, N19063, N19062, N19061, N19060, N19059, N19058, N19057, N19056, N19055, N19054, N19053, N19052, N19051, N19050, N19049, N19048, N19047, N19046, N19045, N19044, N19043, N19042, N19041, N19040, N19039, N19038 } = (N183)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18520)? { N16871, N16870, N16869, N16868, N16867, N16866, N16865, N16864, N16863, N16862, N16861, N16860, N16859, N16858, N16857, N16856, N16855, N16854, N16853, N16852, N16851, N16850, N16849, N16848, N16847, N16846, N16845, N16844, N16843, N16842, N16841, N16840, N16839, N16838, N16837, N16836, N16835, N16834, N16833, N16832, N16831, N16830, N16829, N16828, N16827, N16826, N16825, N16824, N16823, N16822, N16821, N16820, N16819, N16818, N16817, N16816, N16815, N16814, N16813, N16812, N16811, N16810, N16809, N16808 } : 1'b0;
  assign { N19165, N19164, N19163, N19162, N19161, N19160, N19159, N19158, N19157, N19156, N19155, N19154, N19153, N19152, N19151, N19150, N19149, N19148, N19147, N19146, N19145, N19144, N19143, N19142, N19141, N19140, N19139, N19138, N19137, N19136, N19135, N19134, N19133, N19132, N19131, N19130, N19129, N19128, N19127, N19126, N19125, N19124, N19123, N19122, N19121, N19120, N19119, N19118, N19117, N19116, N19115, N19114, N19113, N19112, N19111, N19110, N19109, N19108, N19107, N19106, N19105, N19104, N19103, N19102 } = (N184)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18585)? { N17129, N17128, N17127, N17126, N17125, N17124, N17123, N17122, N17121, N17120, N17119, N17118, N17117, N17116, N17115, N17114, N17113, N17112, N17111, N17110, N17109, N17108, N17107, N17106, N17105, N17104, N17103, N17102, N17101, N17100, N17099, N17098, N17097, N17096, N17095, N17094, N17093, N17092, N17091, N17090, N17089, N17088, N17087, N17086, N17085, N17084, N17083, N17082, N17081, N17080, N17079, N17078, N17077, N17076, N17075, N17074, N17073, N17072, N17071, N17070, N17069, N17068, N17067, N17066 } : 1'b0;
  assign { N19229, N19228, N19227, N19226, N19225, N19224, N19223, N19222, N19221, N19220, N19219, N19218, N19217, N19216, N19215, N19214, N19213, N19212, N19211, N19210, N19209, N19208, N19207, N19206, N19205, N19204, N19203, N19202, N19201, N19200, N19199, N19198, N19197, N19196, N19195, N19194, N19193, N19192, N19191, N19190, N19189, N19188, N19187, N19186, N19185, N19184, N19183, N19182, N19181, N19180, N19179, N19178, N19177, N19176, N19175, N19174, N19173, N19172, N19171, N19170, N19169, N19168, N19167, N19166 } = (N185)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18650)? { N17387, N17386, N17385, N17384, N17383, N17382, N17381, N17380, N17379, N17378, N17377, N17376, N17375, N17374, N17373, N17372, N17371, N17370, N17369, N17368, N17367, N17366, N17365, N17364, N17363, N17362, N17361, N17360, N17359, N17358, N17357, N17356, N17355, N17354, N17353, N17352, N17351, N17350, N17349, N17348, N17347, N17346, N17345, N17344, N17343, N17342, N17341, N17340, N17339, N17338, N17337, N17336, N17335, N17334, N17333, N17332, N17331, N17330, N17329, N17328, N17327, N17326, N17325, N17324 } : 1'b0;
  assign { N19293, N19292, N19291, N19290, N19289, N19288, N19287, N19286, N19285, N19284, N19283, N19282, N19281, N19280, N19279, N19278, N19277, N19276, N19275, N19274, N19273, N19272, N19271, N19270, N19269, N19268, N19267, N19266, N19265, N19264, N19263, N19262, N19261, N19260, N19259, N19258, N19257, N19256, N19255, N19254, N19253, N19252, N19251, N19250, N19249, N19248, N19247, N19246, N19245, N19244, N19243, N19242, N19241, N19240, N19239, N19238, N19237, N19236, N19235, N19234, N19233, N19232, N19231, N19230 } = (N186)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18715)? { N17645, N17644, N17643, N17642, N17641, N17640, N17639, N17638, N17637, N17636, N17635, N17634, N17633, N17632, N17631, N17630, N17629, N17628, N17627, N17626, N17625, N17624, N17623, N17622, N17621, N17620, N17619, N17618, N17617, N17616, N17615, N17614, N17613, N17612, N17611, N17610, N17609, N17608, N17607, N17606, N17605, N17604, N17603, N17602, N17601, N17600, N17599, N17598, N17597, N17596, N17595, N17594, N17593, N17592, N17591, N17590, N17589, N17588, N17587, N17586, N17585, N17584, N17583, N17582 } : 1'b0;
  assign { N19357, N19356, N19355, N19354, N19353, N19352, N19351, N19350, N19349, N19348, N19347, N19346, N19345, N19344, N19343, N19342, N19341, N19340, N19339, N19338, N19337, N19336, N19335, N19334, N19333, N19332, N19331, N19330, N19329, N19328, N19327, N19326, N19325, N19324, N19323, N19322, N19321, N19320, N19319, N19318, N19317, N19316, N19315, N19314, N19313, N19312, N19311, N19310, N19309, N19308, N19307, N19306, N19305, N19304, N19303, N19302, N19301, N19300, N19299, N19298, N19297, N19296, N19295, N19294 } = (N187)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18780)? { N17903, N17902, N17901, N17900, N17899, N17898, N17897, N17896, N17895, N17894, N17893, N17892, N17891, N17890, N17889, N17888, N17887, N17886, N17885, N17884, N17883, N17882, N17881, N17880, N17879, N17878, N17877, N17876, N17875, N17874, N17873, N17872, N17871, N17870, N17869, N17868, N17867, N17866, N17865, N17864, N17863, N17862, N17861, N17860, N17859, N17858, N17857, N17856, N17855, N17854, N17853, N17852, N17851, N17850, N17849, N17848, N17847, N17846, N17845, N17844, N17843, N17842, N17841, N17840 } : 1'b0;
  assign { N19421, N19420, N19419, N19418, N19417, N19416, N19415, N19414, N19413, N19412, N19411, N19410, N19409, N19408, N19407, N19406, N19405, N19404, N19403, N19402, N19401, N19400, N19399, N19398, N19397, N19396, N19395, N19394, N19393, N19392, N19391, N19390, N19389, N19388, N19387, N19386, N19385, N19384, N19383, N19382, N19381, N19380, N19379, N19378, N19377, N19376, N19375, N19374, N19373, N19372, N19371, N19370, N19369, N19368, N19367, N19366, N19365, N19364, N19363, N19362, N19361, N19360, N19359, N19358 } = (N188)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18845)? { N18161, N18160, N18159, N18158, N18157, N18156, N18155, N18154, N18153, N18152, N18151, N18150, N18149, N18148, N18147, N18146, N18145, N18144, N18143, N18142, N18141, N18140, N18139, N18138, N18137, N18136, N18135, N18134, N18133, N18132, N18131, N18130, N18129, N18128, N18127, N18126, N18125, N18124, N18123, N18122, N18121, N18120, N18119, N18118, N18117, N18116, N18115, N18114, N18113, N18112, N18111, N18110, N18109, N18108, N18107, N18106, N18105, N18104, N18103, N18102, N18101, N18100, N18099, N18098 } : 1'b0;
  assign { N19555, N19554, N19553, N19552, N19551, N19550, N19549, N19548, N19547, N19546, N19545, N19544, N19543, N19542, N19541, N19540, N19539, N19538, N19537, N19536, N19535, N19534, N19533, N19532, N19531, N19530, N19529, N19528, N19527, N19526, N19525, N19524, N19523, N19522, N19521, N19520, N19519, N19518, N19517, N19516, N19515, N19514, N19513, N19512, N19511, N19510, N19509, N19508, N19507, N19506, N19505, N19504, N19503, N19502, N19501, N19500, N19499, N19498, N19497, N19496, N19495, N19494, N19493, N19492, N19491, N19490, N19489, N19488, N19487, N19486, N19485, N19484, N19483, N19482, N19481, N19480, N19479, N19478, N19477, N19476, N19475, N19474, N19473, N19472, N19471, N19470, N19469, N19468, N19467, N19466, N19465, N19464, N19463, N19462, N19461, N19460, N19459, N19458, N19457, N19456, N19455, N19454, N19453, N19452, N19451, N19450, N19449, N19448, N19447, N19446, N19445, N19444, N19443, N19442, N19441, N19440, N19439, N19438, N19437, N19436, N19435, N19434, N19433, N19432, N19431, N19430, N19429, N19428, N19427 } = (N181)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18390)? { N16484, N16483, N16482, N16481, N16480, N16479, N16478, N16477, N16476, N16475, N16474, N16473, N16472, N16471, N16470, N16469, N16468, N16467, N16466, N16465, N16464, N16463, N16462, N16461, N16460, N16459, N16458, N16457, N16456, N16455, N16454, N16453, N16452, N16451, N16450, N16449, N16448, N16447, N16446, N16445, N16444, N16443, N16442, N16441, N16440, N16439, N16438, N16437, N16436, N16435, N16434, N16433, N16432, N16431, N16430, N16429, N16428, N16427, N16426, N16425, N16424, N16423, N16422, N16421, N16420, N16419, N16418, N16417, N16416, N16415, N16414, N16413, N16412, N16411, N16410, N16409, N16408, N16407, N16406, N16405, N16404, N16403, N16402, N16401, N16400, N16399, N16398, N16397, N16396, N16395, N16394, N16393, N16392, N16391, N16390, N16389, N16388, N16387, N16386, N16385, N16384, N16383, N16382, N16381, N16380, N16379, N16378, N16377, N16376, N16375, N16374, N16373, N16372, N16371, N16370, N16369, N16368, N16367, N16366, N16365, N16364, N16363, N16362, N16361, N16360, N16359, N16358, N16357, N16356 } : 1'b0;
  assign { N19684, N19683, N19682, N19681, N19680, N19679, N19678, N19677, N19676, N19675, N19674, N19673, N19672, N19671, N19670, N19669, N19668, N19667, N19666, N19665, N19664, N19663, N19662, N19661, N19660, N19659, N19658, N19657, N19656, N19655, N19654, N19653, N19652, N19651, N19650, N19649, N19648, N19647, N19646, N19645, N19644, N19643, N19642, N19641, N19640, N19639, N19638, N19637, N19636, N19635, N19634, N19633, N19632, N19631, N19630, N19629, N19628, N19627, N19626, N19625, N19624, N19623, N19622, N19621, N19620, N19619, N19618, N19617, N19616, N19615, N19614, N19613, N19612, N19611, N19610, N19609, N19608, N19607, N19606, N19605, N19604, N19603, N19602, N19601, N19600, N19599, N19598, N19597, N19596, N19595, N19594, N19593, N19592, N19591, N19590, N19589, N19588, N19587, N19586, N19585, N19584, N19583, N19582, N19581, N19580, N19579, N19578, N19577, N19576, N19575, N19574, N19573, N19572, N19571, N19570, N19569, N19568, N19567, N19566, N19565, N19564, N19563, N19562, N19561, N19560, N19559, N19558, N19557, N19556 } = (N182)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18455)? { N16742, N16741, N16740, N16739, N16738, N16737, N16736, N16735, N16734, N16733, N16732, N16731, N16730, N16729, N16728, N16727, N16726, N16725, N16724, N16723, N16722, N16721, N16720, N16719, N16718, N16717, N16716, N16715, N16714, N16713, N16712, N16711, N16710, N16709, N16708, N16707, N16706, N16705, N16704, N16703, N16702, N16701, N16700, N16699, N16698, N16697, N16696, N16695, N16694, N16693, N16692, N16691, N16690, N16689, N16688, N16687, N16686, N16685, N16684, N16683, N16682, N16681, N16680, N16679, N16678, N16677, N16676, N16675, N16674, N16673, N16672, N16671, N16670, N16669, N16668, N16667, N16666, N16665, N16664, N16663, N16662, N16661, N16660, N16659, N16658, N16657, N16656, N16655, N16654, N16653, N16652, N16651, N16650, N16649, N16648, N16647, N16646, N16645, N16644, N16643, N16642, N16641, N16640, N16639, N16638, N16637, N16636, N16635, N16634, N16633, N16632, N16631, N16630, N16629, N16628, N16627, N16626, N16625, N16624, N16623, N16622, N16621, N16620, N16619, N16618, N16617, N16616, N16615, N16614 } : 1'b0;
  assign { N19813, N19812, N19811, N19810, N19809, N19808, N19807, N19806, N19805, N19804, N19803, N19802, N19801, N19800, N19799, N19798, N19797, N19796, N19795, N19794, N19793, N19792, N19791, N19790, N19789, N19788, N19787, N19786, N19785, N19784, N19783, N19782, N19781, N19780, N19779, N19778, N19777, N19776, N19775, N19774, N19773, N19772, N19771, N19770, N19769, N19768, N19767, N19766, N19765, N19764, N19763, N19762, N19761, N19760, N19759, N19758, N19757, N19756, N19755, N19754, N19753, N19752, N19751, N19750, N19749, N19748, N19747, N19746, N19745, N19744, N19743, N19742, N19741, N19740, N19739, N19738, N19737, N19736, N19735, N19734, N19733, N19732, N19731, N19730, N19729, N19728, N19727, N19726, N19725, N19724, N19723, N19722, N19721, N19720, N19719, N19718, N19717, N19716, N19715, N19714, N19713, N19712, N19711, N19710, N19709, N19708, N19707, N19706, N19705, N19704, N19703, N19702, N19701, N19700, N19699, N19698, N19697, N19696, N19695, N19694, N19693, N19692, N19691, N19690, N19689, N19688, N19687, N19686, N19685 } = (N183)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18520)? { N17000, N16999, N16998, N16997, N16996, N16995, N16994, N16993, N16992, N16991, N16990, N16989, N16988, N16987, N16986, N16985, N16984, N16983, N16982, N16981, N16980, N16979, N16978, N16977, N16976, N16975, N16974, N16973, N16972, N16971, N16970, N16969, N16968, N16967, N16966, N16965, N16964, N16963, N16962, N16961, N16960, N16959, N16958, N16957, N16956, N16955, N16954, N16953, N16952, N16951, N16950, N16949, N16948, N16947, N16946, N16945, N16944, N16943, N16942, N16941, N16940, N16939, N16938, N16937, N16936, N16935, N16934, N16933, N16932, N16931, N16930, N16929, N16928, N16927, N16926, N16925, N16924, N16923, N16922, N16921, N16920, N16919, N16918, N16917, N16916, N16915, N16914, N16913, N16912, N16911, N16910, N16909, N16908, N16907, N16906, N16905, N16904, N16903, N16902, N16901, N16900, N16899, N16898, N16897, N16896, N16895, N16894, N16893, N16892, N16891, N16890, N16889, N16888, N16887, N16886, N16885, N16884, N16883, N16882, N16881, N16880, N16879, N16878, N16877, N16876, N16875, N16874, N16873, N16872 } : 1'b0;
  assign { N19942, N19941, N19940, N19939, N19938, N19937, N19936, N19935, N19934, N19933, N19932, N19931, N19930, N19929, N19928, N19927, N19926, N19925, N19924, N19923, N19922, N19921, N19920, N19919, N19918, N19917, N19916, N19915, N19914, N19913, N19912, N19911, N19910, N19909, N19908, N19907, N19906, N19905, N19904, N19903, N19902, N19901, N19900, N19899, N19898, N19897, N19896, N19895, N19894, N19893, N19892, N19891, N19890, N19889, N19888, N19887, N19886, N19885, N19884, N19883, N19882, N19881, N19880, N19879, N19878, N19877, N19876, N19875, N19874, N19873, N19872, N19871, N19870, N19869, N19868, N19867, N19866, N19865, N19864, N19863, N19862, N19861, N19860, N19859, N19858, N19857, N19856, N19855, N19854, N19853, N19852, N19851, N19850, N19849, N19848, N19847, N19846, N19845, N19844, N19843, N19842, N19841, N19840, N19839, N19838, N19837, N19836, N19835, N19834, N19833, N19832, N19831, N19830, N19829, N19828, N19827, N19826, N19825, N19824, N19823, N19822, N19821, N19820, N19819, N19818, N19817, N19816, N19815, N19814 } = (N184)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18585)? { N17258, N17257, N17256, N17255, N17254, N17253, N17252, N17251, N17250, N17249, N17248, N17247, N17246, N17245, N17244, N17243, N17242, N17241, N17240, N17239, N17238, N17237, N17236, N17235, N17234, N17233, N17232, N17231, N17230, N17229, N17228, N17227, N17226, N17225, N17224, N17223, N17222, N17221, N17220, N17219, N17218, N17217, N17216, N17215, N17214, N17213, N17212, N17211, N17210, N17209, N17208, N17207, N17206, N17205, N17204, N17203, N17202, N17201, N17200, N17199, N17198, N17197, N17196, N17195, N17194, N17193, N17192, N17191, N17190, N17189, N17188, N17187, N17186, N17185, N17184, N17183, N17182, N17181, N17180, N17179, N17178, N17177, N17176, N17175, N17174, N17173, N17172, N17171, N17170, N17169, N17168, N17167, N17166, N17165, N17164, N17163, N17162, N17161, N17160, N17159, N17158, N17157, N17156, N17155, N17154, N17153, N17152, N17151, N17150, N17149, N17148, N17147, N17146, N17145, N17144, N17143, N17142, N17141, N17140, N17139, N17138, N17137, N17136, N17135, N17134, N17133, N17132, N17131, N17130 } : 1'b0;
  assign { N20071, N20070, N20069, N20068, N20067, N20066, N20065, N20064, N20063, N20062, N20061, N20060, N20059, N20058, N20057, N20056, N20055, N20054, N20053, N20052, N20051, N20050, N20049, N20048, N20047, N20046, N20045, N20044, N20043, N20042, N20041, N20040, N20039, N20038, N20037, N20036, N20035, N20034, N20033, N20032, N20031, N20030, N20029, N20028, N20027, N20026, N20025, N20024, N20023, N20022, N20021, N20020, N20019, N20018, N20017, N20016, N20015, N20014, N20013, N20012, N20011, N20010, N20009, N20008, N20007, N20006, N20005, N20004, N20003, N20002, N20001, N20000, N19999, N19998, N19997, N19996, N19995, N19994, N19993, N19992, N19991, N19990, N19989, N19988, N19987, N19986, N19985, N19984, N19983, N19982, N19981, N19980, N19979, N19978, N19977, N19976, N19975, N19974, N19973, N19972, N19971, N19970, N19969, N19968, N19967, N19966, N19965, N19964, N19963, N19962, N19961, N19960, N19959, N19958, N19957, N19956, N19955, N19954, N19953, N19952, N19951, N19950, N19949, N19948, N19947, N19946, N19945, N19944, N19943 } = (N185)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18650)? { N17516, N17515, N17514, N17513, N17512, N17511, N17510, N17509, N17508, N17507, N17506, N17505, N17504, N17503, N17502, N17501, N17500, N17499, N17498, N17497, N17496, N17495, N17494, N17493, N17492, N17491, N17490, N17489, N17488, N17487, N17486, N17485, N17484, N17483, N17482, N17481, N17480, N17479, N17478, N17477, N17476, N17475, N17474, N17473, N17472, N17471, N17470, N17469, N17468, N17467, N17466, N17465, N17464, N17463, N17462, N17461, N17460, N17459, N17458, N17457, N17456, N17455, N17454, N17453, N17452, N17451, N17450, N17449, N17448, N17447, N17446, N17445, N17444, N17443, N17442, N17441, N17440, N17439, N17438, N17437, N17436, N17435, N17434, N17433, N17432, N17431, N17430, N17429, N17428, N17427, N17426, N17425, N17424, N17423, N17422, N17421, N17420, N17419, N17418, N17417, N17416, N17415, N17414, N17413, N17412, N17411, N17410, N17409, N17408, N17407, N17406, N17405, N17404, N17403, N17402, N17401, N17400, N17399, N17398, N17397, N17396, N17395, N17394, N17393, N17392, N17391, N17390, N17389, N17388 } : 1'b0;
  assign { N20200, N20199, N20198, N20197, N20196, N20195, N20194, N20193, N20192, N20191, N20190, N20189, N20188, N20187, N20186, N20185, N20184, N20183, N20182, N20181, N20180, N20179, N20178, N20177, N20176, N20175, N20174, N20173, N20172, N20171, N20170, N20169, N20168, N20167, N20166, N20165, N20164, N20163, N20162, N20161, N20160, N20159, N20158, N20157, N20156, N20155, N20154, N20153, N20152, N20151, N20150, N20149, N20148, N20147, N20146, N20145, N20144, N20143, N20142, N20141, N20140, N20139, N20138, N20137, N20136, N20135, N20134, N20133, N20132, N20131, N20130, N20129, N20128, N20127, N20126, N20125, N20124, N20123, N20122, N20121, N20120, N20119, N20118, N20117, N20116, N20115, N20114, N20113, N20112, N20111, N20110, N20109, N20108, N20107, N20106, N20105, N20104, N20103, N20102, N20101, N20100, N20099, N20098, N20097, N20096, N20095, N20094, N20093, N20092, N20091, N20090, N20089, N20088, N20087, N20086, N20085, N20084, N20083, N20082, N20081, N20080, N20079, N20078, N20077, N20076, N20075, N20074, N20073, N20072 } = (N186)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18715)? { N17774, N17773, N17772, N17771, N17770, N17769, N17768, N17767, N17766, N17765, N17764, N17763, N17762, N17761, N17760, N17759, N17758, N17757, N17756, N17755, N17754, N17753, N17752, N17751, N17750, N17749, N17748, N17747, N17746, N17745, N17744, N17743, N17742, N17741, N17740, N17739, N17738, N17737, N17736, N17735, N17734, N17733, N17732, N17731, N17730, N17729, N17728, N17727, N17726, N17725, N17724, N17723, N17722, N17721, N17720, N17719, N17718, N17717, N17716, N17715, N17714, N17713, N17712, N17711, N17710, N17709, N17708, N17707, N17706, N17705, N17704, N17703, N17702, N17701, N17700, N17699, N17698, N17697, N17696, N17695, N17694, N17693, N17692, N17691, N17690, N17689, N17688, N17687, N17686, N17685, N17684, N17683, N17682, N17681, N17680, N17679, N17678, N17677, N17676, N17675, N17674, N17673, N17672, N17671, N17670, N17669, N17668, N17667, N17666, N17665, N17664, N17663, N17662, N17661, N17660, N17659, N17658, N17657, N17656, N17655, N17654, N17653, N17652, N17651, N17650, N17649, N17648, N17647, N17646 } : 1'b0;
  assign { N20329, N20328, N20327, N20326, N20325, N20324, N20323, N20322, N20321, N20320, N20319, N20318, N20317, N20316, N20315, N20314, N20313, N20312, N20311, N20310, N20309, N20308, N20307, N20306, N20305, N20304, N20303, N20302, N20301, N20300, N20299, N20298, N20297, N20296, N20295, N20294, N20293, N20292, N20291, N20290, N20289, N20288, N20287, N20286, N20285, N20284, N20283, N20282, N20281, N20280, N20279, N20278, N20277, N20276, N20275, N20274, N20273, N20272, N20271, N20270, N20269, N20268, N20267, N20266, N20265, N20264, N20263, N20262, N20261, N20260, N20259, N20258, N20257, N20256, N20255, N20254, N20253, N20252, N20251, N20250, N20249, N20248, N20247, N20246, N20245, N20244, N20243, N20242, N20241, N20240, N20239, N20238, N20237, N20236, N20235, N20234, N20233, N20232, N20231, N20230, N20229, N20228, N20227, N20226, N20225, N20224, N20223, N20222, N20221, N20220, N20219, N20218, N20217, N20216, N20215, N20214, N20213, N20212, N20211, N20210, N20209, N20208, N20207, N20206, N20205, N20204, N20203, N20202, N20201 } = (N187)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18780)? { N18032, N18031, N18030, N18029, N18028, N18027, N18026, N18025, N18024, N18023, N18022, N18021, N18020, N18019, N18018, N18017, N18016, N18015, N18014, N18013, N18012, N18011, N18010, N18009, N18008, N18007, N18006, N18005, N18004, N18003, N18002, N18001, N18000, N17999, N17998, N17997, N17996, N17995, N17994, N17993, N17992, N17991, N17990, N17989, N17988, N17987, N17986, N17985, N17984, N17983, N17982, N17981, N17980, N17979, N17978, N17977, N17976, N17975, N17974, N17973, N17972, N17971, N17970, N17969, N17968, N17967, N17966, N17965, N17964, N17963, N17962, N17961, N17960, N17959, N17958, N17957, N17956, N17955, N17954, N17953, N17952, N17951, N17950, N17949, N17948, N17947, N17946, N17945, N17944, N17943, N17942, N17941, N17940, N17939, N17938, N17937, N17936, N17935, N17934, N17933, N17932, N17931, N17930, N17929, N17928, N17927, N17926, N17925, N17924, N17923, N17922, N17921, N17920, N17919, N17918, N17917, N17916, N17915, N17914, N17913, N17912, N17911, N17910, N17909, N17908, N17907, N17906, N17905, N17904 } : 1'b0;
  assign { N20458, N20457, N20456, N20455, N20454, N20453, N20452, N20451, N20450, N20449, N20448, N20447, N20446, N20445, N20444, N20443, N20442, N20441, N20440, N20439, N20438, N20437, N20436, N20435, N20434, N20433, N20432, N20431, N20430, N20429, N20428, N20427, N20426, N20425, N20424, N20423, N20422, N20421, N20420, N20419, N20418, N20417, N20416, N20415, N20414, N20413, N20412, N20411, N20410, N20409, N20408, N20407, N20406, N20405, N20404, N20403, N20402, N20401, N20400, N20399, N20398, N20397, N20396, N20395, N20394, N20393, N20392, N20391, N20390, N20389, N20388, N20387, N20386, N20385, N20384, N20383, N20382, N20381, N20380, N20379, N20378, N20377, N20376, N20375, N20374, N20373, N20372, N20371, N20370, N20369, N20368, N20367, N20366, N20365, N20364, N20363, N20362, N20361, N20360, N20359, N20358, N20357, N20356, N20355, N20354, N20353, N20352, N20351, N20350, N20349, N20348, N20347, N20346, N20345, N20344, N20343, N20342, N20341, N20340, N20339, N20338, N20337, N20336, N20335, N20334, N20333, N20332, N20331, N20330 } = (N188)? ex_i[386:258] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N18845)? { N18290, N18289, N18288, N18287, N18286, N18285, N18284, N18283, N18282, N18281, N18280, N18279, N18278, N18277, N18276, N18275, N18274, N18273, N18272, N18271, N18270, N18269, N18268, N18267, N18266, N18265, N18264, N18263, N18262, N18261, N18260, N18259, N18258, N18257, N18256, N18255, N18254, N18253, N18252, N18251, N18250, N18249, N18248, N18247, N18246, N18245, N18244, N18243, N18242, N18241, N18240, N18239, N18238, N18237, N18236, N18235, N18234, N18233, N18232, N18231, N18230, N18229, N18228, N18227, N18226, N18225, N18224, N18223, N18222, N18221, N18220, N18219, N18218, N18217, N18216, N18215, N18214, N18213, N18212, N18211, N18210, N18209, N18208, N18207, N18206, N18205, N18204, N18203, N18202, N18201, N18200, N18199, N18198, N18197, N18196, N18195, N18194, N18193, N18192, N18191, N18190, N18189, N18188, N18187, N18186, N18185, N18184, N18183, N18182, N18181, N18180, N18179, N18178, N18177, N18176, N18175, N18174, N18173, N18172, N18171, N18170, N18169, N18168, N18167, N18166, N18165, N18164, N18163, N18162 } : 1'b0;
  assign { N20534, N20533, N20532, N20531, N20530, N20529, N20528, N20527, N20526, N20525, N20524, N20523, N20522, N20521, N20520, N20519, N20518, N20517, N20516, N20515, N20514, N20513, N20512, N20511, N20510, N20509, N20508, N20507, N20506, N20505, N20504, N20503, N20502, N20501, N20500, N20499, N20498, N20497, N20496, N20495, N20494, N20493, N20492, N20491, N20490, N20489, N20488, N20487, N20486, N20485, N20484, N20483, N20482, N20481, N20480, N20479, N20478, N20477, N20476, N20475, N20474, N20473, N20472, N20471 } = (N181)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18390)? { N16484, N16483, N16482, N16481, N16480, N16479, N16478, N16477, N16476, N16475, N16474, N16473, N16472, N16471, N16470, N16469, N16468, N16467, N16466, N16465, N16464, N16463, N16462, N16461, N16460, N16459, N16458, N16457, N16456, N16455, N16454, N16453, N16452, N16451, N16450, N16449, N16448, N16447, N16446, N16445, N16444, N16443, N16442, N16441, N16440, N16439, N16438, N16437, N16436, N16435, N16434, N16433, N16432, N16431, N16430, N16429, N16428, N16427, N16426, N16425, N16424, N16423, N16422, N16421 } : 1'b0;
  assign { N20598, N20597, N20596, N20595, N20594, N20593, N20592, N20591, N20590, N20589, N20588, N20587, N20586, N20585, N20584, N20583, N20582, N20581, N20580, N20579, N20578, N20577, N20576, N20575, N20574, N20573, N20572, N20571, N20570, N20569, N20568, N20567, N20566, N20565, N20564, N20563, N20562, N20561, N20560, N20559, N20558, N20557, N20556, N20555, N20554, N20553, N20552, N20551, N20550, N20549, N20548, N20547, N20546, N20545, N20544, N20543, N20542, N20541, N20540, N20539, N20538, N20537, N20536, N20535 } = (N182)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18455)? { N16742, N16741, N16740, N16739, N16738, N16737, N16736, N16735, N16734, N16733, N16732, N16731, N16730, N16729, N16728, N16727, N16726, N16725, N16724, N16723, N16722, N16721, N16720, N16719, N16718, N16717, N16716, N16715, N16714, N16713, N16712, N16711, N16710, N16709, N16708, N16707, N16706, N16705, N16704, N16703, N16702, N16701, N16700, N16699, N16698, N16697, N16696, N16695, N16694, N16693, N16692, N16691, N16690, N16689, N16688, N16687, N16686, N16685, N16684, N16683, N16682, N16681, N16680, N16679 } : 1'b0;
  assign { N20662, N20661, N20660, N20659, N20658, N20657, N20656, N20655, N20654, N20653, N20652, N20651, N20650, N20649, N20648, N20647, N20646, N20645, N20644, N20643, N20642, N20641, N20640, N20639, N20638, N20637, N20636, N20635, N20634, N20633, N20632, N20631, N20630, N20629, N20628, N20627, N20626, N20625, N20624, N20623, N20622, N20621, N20620, N20619, N20618, N20617, N20616, N20615, N20614, N20613, N20612, N20611, N20610, N20609, N20608, N20607, N20606, N20605, N20604, N20603, N20602, N20601, N20600, N20599 } = (N183)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18520)? { N17000, N16999, N16998, N16997, N16996, N16995, N16994, N16993, N16992, N16991, N16990, N16989, N16988, N16987, N16986, N16985, N16984, N16983, N16982, N16981, N16980, N16979, N16978, N16977, N16976, N16975, N16974, N16973, N16972, N16971, N16970, N16969, N16968, N16967, N16966, N16965, N16964, N16963, N16962, N16961, N16960, N16959, N16958, N16957, N16956, N16955, N16954, N16953, N16952, N16951, N16950, N16949, N16948, N16947, N16946, N16945, N16944, N16943, N16942, N16941, N16940, N16939, N16938, N16937 } : 1'b0;
  assign { N20726, N20725, N20724, N20723, N20722, N20721, N20720, N20719, N20718, N20717, N20716, N20715, N20714, N20713, N20712, N20711, N20710, N20709, N20708, N20707, N20706, N20705, N20704, N20703, N20702, N20701, N20700, N20699, N20698, N20697, N20696, N20695, N20694, N20693, N20692, N20691, N20690, N20689, N20688, N20687, N20686, N20685, N20684, N20683, N20682, N20681, N20680, N20679, N20678, N20677, N20676, N20675, N20674, N20673, N20672, N20671, N20670, N20669, N20668, N20667, N20666, N20665, N20664, N20663 } = (N184)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18585)? { N17258, N17257, N17256, N17255, N17254, N17253, N17252, N17251, N17250, N17249, N17248, N17247, N17246, N17245, N17244, N17243, N17242, N17241, N17240, N17239, N17238, N17237, N17236, N17235, N17234, N17233, N17232, N17231, N17230, N17229, N17228, N17227, N17226, N17225, N17224, N17223, N17222, N17221, N17220, N17219, N17218, N17217, N17216, N17215, N17214, N17213, N17212, N17211, N17210, N17209, N17208, N17207, N17206, N17205, N17204, N17203, N17202, N17201, N17200, N17199, N17198, N17197, N17196, N17195 } : 1'b0;
  assign { N20790, N20789, N20788, N20787, N20786, N20785, N20784, N20783, N20782, N20781, N20780, N20779, N20778, N20777, N20776, N20775, N20774, N20773, N20772, N20771, N20770, N20769, N20768, N20767, N20766, N20765, N20764, N20763, N20762, N20761, N20760, N20759, N20758, N20757, N20756, N20755, N20754, N20753, N20752, N20751, N20750, N20749, N20748, N20747, N20746, N20745, N20744, N20743, N20742, N20741, N20740, N20739, N20738, N20737, N20736, N20735, N20734, N20733, N20732, N20731, N20730, N20729, N20728, N20727 } = (N185)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18650)? { N17516, N17515, N17514, N17513, N17512, N17511, N17510, N17509, N17508, N17507, N17506, N17505, N17504, N17503, N17502, N17501, N17500, N17499, N17498, N17497, N17496, N17495, N17494, N17493, N17492, N17491, N17490, N17489, N17488, N17487, N17486, N17485, N17484, N17483, N17482, N17481, N17480, N17479, N17478, N17477, N17476, N17475, N17474, N17473, N17472, N17471, N17470, N17469, N17468, N17467, N17466, N17465, N17464, N17463, N17462, N17461, N17460, N17459, N17458, N17457, N17456, N17455, N17454, N17453 } : 1'b0;
  assign { N20854, N20853, N20852, N20851, N20850, N20849, N20848, N20847, N20846, N20845, N20844, N20843, N20842, N20841, N20840, N20839, N20838, N20837, N20836, N20835, N20834, N20833, N20832, N20831, N20830, N20829, N20828, N20827, N20826, N20825, N20824, N20823, N20822, N20821, N20820, N20819, N20818, N20817, N20816, N20815, N20814, N20813, N20812, N20811, N20810, N20809, N20808, N20807, N20806, N20805, N20804, N20803, N20802, N20801, N20800, N20799, N20798, N20797, N20796, N20795, N20794, N20793, N20792, N20791 } = (N186)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18715)? { N17774, N17773, N17772, N17771, N17770, N17769, N17768, N17767, N17766, N17765, N17764, N17763, N17762, N17761, N17760, N17759, N17758, N17757, N17756, N17755, N17754, N17753, N17752, N17751, N17750, N17749, N17748, N17747, N17746, N17745, N17744, N17743, N17742, N17741, N17740, N17739, N17738, N17737, N17736, N17735, N17734, N17733, N17732, N17731, N17730, N17729, N17728, N17727, N17726, N17725, N17724, N17723, N17722, N17721, N17720, N17719, N17718, N17717, N17716, N17715, N17714, N17713, N17712, N17711 } : 1'b0;
  assign { N20918, N20917, N20916, N20915, N20914, N20913, N20912, N20911, N20910, N20909, N20908, N20907, N20906, N20905, N20904, N20903, N20902, N20901, N20900, N20899, N20898, N20897, N20896, N20895, N20894, N20893, N20892, N20891, N20890, N20889, N20888, N20887, N20886, N20885, N20884, N20883, N20882, N20881, N20880, N20879, N20878, N20877, N20876, N20875, N20874, N20873, N20872, N20871, N20870, N20869, N20868, N20867, N20866, N20865, N20864, N20863, N20862, N20861, N20860, N20859, N20858, N20857, N20856, N20855 } = (N187)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18780)? { N18032, N18031, N18030, N18029, N18028, N18027, N18026, N18025, N18024, N18023, N18022, N18021, N18020, N18019, N18018, N18017, N18016, N18015, N18014, N18013, N18012, N18011, N18010, N18009, N18008, N18007, N18006, N18005, N18004, N18003, N18002, N18001, N18000, N17999, N17998, N17997, N17996, N17995, N17994, N17993, N17992, N17991, N17990, N17989, N17988, N17987, N17986, N17985, N17984, N17983, N17982, N17981, N17980, N17979, N17978, N17977, N17976, N17975, N17974, N17973, N17972, N17971, N17970, N17969 } : 1'b0;
  assign { N20982, N20981, N20980, N20979, N20978, N20977, N20976, N20975, N20974, N20973, N20972, N20971, N20970, N20969, N20968, N20967, N20966, N20965, N20964, N20963, N20962, N20961, N20960, N20959, N20958, N20957, N20956, N20955, N20954, N20953, N20952, N20951, N20950, N20949, N20948, N20947, N20946, N20945, N20944, N20943, N20942, N20941, N20940, N20939, N20938, N20937, N20936, N20935, N20934, N20933, N20932, N20931, N20930, N20929, N20928, N20927, N20926, N20925, N20924, N20923, N20922, N20921, N20920, N20919 } = (N188)? ex_i[386:323] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18845)? { N18290, N18289, N18288, N18287, N18286, N18285, N18284, N18283, N18282, N18281, N18280, N18279, N18278, N18277, N18276, N18275, N18274, N18273, N18272, N18271, N18270, N18269, N18268, N18267, N18266, N18265, N18264, N18263, N18262, N18261, N18260, N18259, N18258, N18257, N18256, N18255, N18254, N18253, N18252, N18251, N18250, N18249, N18248, N18247, N18246, N18245, N18244, N18243, N18242, N18241, N18240, N18239, N18238, N18237, N18236, N18235, N18234, N18233, N18232, N18231, N18230, N18229, N18228, N18227 } : 1'b0;
  assign { N21494, N21493, N21492, N21491, N21490, N21489, N21488, N21487, N21486, N21485, N21484, N21483, N21482, N21481, N21480, N21479, N21478, N21477, N21476, N21475, N21474, N21473, N21472, N21471, N21470, N21469, N21468, N21467, N21466, N21465, N21464, N21463, N21462, N21461, N21460, N21459, N21458, N21457, N21456, N21455, N21454, N21453, N21452, N21451, N21450, N21449, N21448, N21447, N21446, N21445, N21444, N21443, N21442, N21441, N21440, N21439, N21438, N21437, N21436, N21435, N21434, N21433, N21432, N21431, N21430, N21429, N21428, N21427, N21426, N21425, N21424, N21423, N21422, N21421, N21420, N21419, N21418, N21417, N21416, N21415, N21414, N21413, N21412, N21411, N21410, N21409, N21408, N21407, N21406, N21405, N21404, N21403, N21402, N21401, N21400, N21399, N21398, N21397, N21396, N21395, N21394, N21393, N21392, N21391, N21390, N21389, N21388, N21387, N21386, N21385, N21384, N21383, N21382, N21381, N21380, N21379, N21378, N21377, N21376, N21375, N21374, N21373, N21372, N21371, N21370, N21369, N21368, N21367, N21366, N21365, N21364, N21363, N21362, N21361, N21360, N21359, N21358, N21357, N21356, N21355, N21354, N21353, N21352, N21351, N21350, N21349, N21348, N21347, N21346, N21345, N21344, N21343, N21342, N21341, N21340, N21339, N21338, N21337, N21336, N21335, N21334, N21333, N21332, N21331, N21330, N21329, N21328, N21327, N21326, N21325, N21324, N21323, N21322, N21321, N21320, N21319, N21318, N21317, N21316, N21315, N21314, N21313, N21312, N21311, N21310, N21309, N21308, N21307, N21306, N21305, N21304, N21303, N21302, N21301, N21300, N21299, N21298, N21297, N21296, N21295, N21294, N21293, N21292, N21291, N21290, N21289, N21288, N21287, N21286, N21285, N21284, N21283, N21282, N21281, N21280, N21279, N21278, N21277, N21276, N21275, N21274, N21273, N21272, N21271, N21270, N21269, N21268, N21267, N21266, N21265, N21264, N21263, N21262, N21261, N21260, N21259, N21258, N21257, N21256, N21255, N21254, N21253, N21252, N21251, N21250, N21249, N21248, N21247, N21246, N21245, N21244, N21243, N21242, N21241, N21240, N21239, N21238, N21237, N21236, N21235, N21234, N21233, N21232, N21231, N21230, N21229, N21228, N21227, N21226, N21225, N21224, N21223, N21222, N21221, N21220, N21219, N21218, N21217, N21216, N21215, N21214, N21213, N21212, N21211, N21210, N21209, N21208, N21207, N21206, N21205, N21204, N21203, N21202, N21201, N21200, N21199, N21198, N21197, N21196, N21195, N21194, N21193, N21192, N21191, N21190, N21189, N21188, N21187, N21186, N21185, N21184, N21183, N21182, N21181, N21180, N21179, N21178, N21177, N21176, N21175, N21174, N21173, N21172, N21171, N21170, N21169, N21168, N21167, N21166, N21165, N21164, N21163, N21162, N21161, N21160, N21159, N21158, N21157, N21156, N21155, N21154, N21153, N21152, N21151, N21150, N21149, N21148, N21147, N21146, N21145, N21144, N21143, N21142, N21141, N21140, N21139, N21138, N21137, N21136, N21135, N21134, N21133, N21132, N21131, N21130, N21129, N21128, N21127, N21126, N21125, N21124, N21123, N21122, N21121, N21120, N21119, N21118, N21117, N21116, N21115, N21114, N21113, N21112, N21111, N21110, N21109, N21108, N21107, N21106, N21105, N21104, N21103, N21102, N21101, N21100, N21099, N21098, N21097, N21096, N21095, N21094, N21093, N21092, N21091, N21090, N21089, N21088, N21087, N21086, N21085, N21084, N21083, N21082, N21081, N21080, N21079, N21078, N21077, N21076, N21075, N21074, N21073, N21072, N21071, N21070, N21069, N21068, N21067, N21066, N21065, N21064, N21063, N21062, N21061, N21060, N21059, N21058, N21057, N21056, N21055, N21054, N21053, N21052, N21051, N21050, N21049, N21048, N21047, N21046, N21045, N21044, N21043, N21042, N21041, N21040, N21039, N21038, N21037, N21036, N21035, N21034, N21033, N21032, N21031, N21030, N21029, N21028, N21027, N21026, N21025, N21024, N21023, N21022, N21021, N21020, N21019, N21018, N21017, N21016, N21015, N21014, N21013, N21012, N21011, N21010, N21009, N21008, N21007, N21006, N21005, N21004, N21003, N21002, N21001, N21000, N20999, N20998, N20997, N20996, N20995, N20994, N20993, N20992, N20991, N20990, N20989, N20988, N20987, N20986, N20985, N20984, N20983 } = (N189)? { N20982, N20981, N20980, N20979, N20978, N20977, N20976, N20975, N20974, N20973, N20972, N20971, N20970, N20969, N20968, N20967, N20966, N20965, N20964, N20963, N20962, N20961, N20960, N20959, N20958, N20957, N20956, N20955, N20954, N20953, N20952, N20951, N20950, N20949, N20948, N20947, N20946, N20945, N20944, N20943, N20942, N20941, N20940, N20939, N20938, N20937, N20936, N20935, N20934, N20933, N20932, N20931, N20930, N20929, N20928, N20927, N20926, N20925, N20924, N20923, N20922, N20921, N20920, N20919, N20918, N20917, N20916, N20915, N20914, N20913, N20912, N20911, N20910, N20909, N20908, N20907, N20906, N20905, N20904, N20903, N20902, N20901, N20900, N20899, N20898, N20897, N20896, N20895, N20894, N20893, N20892, N20891, N20890, N20889, N20888, N20887, N20886, N20885, N20884, N20883, N20882, N20881, N20880, N20879, N20878, N20877, N20876, N20875, N20874, N20873, N20872, N20871, N20870, N20869, N20868, N20867, N20866, N20865, N20864, N20863, N20862, N20861, N20860, N20859, N20858, N20857, N20856, N20855, N20854, N20853, N20852, N20851, N20850, N20849, N20848, N20847, N20846, N20845, N20844, N20843, N20842, N20841, N20840, N20839, N20838, N20837, N20836, N20835, N20834, N20833, N20832, N20831, N20830, N20829, N20828, N20827, N20826, N20825, N20824, N20823, N20822, N20821, N20820, N20819, N20818, N20817, N20816, N20815, N20814, N20813, N20812, N20811, N20810, N20809, N20808, N20807, N20806, N20805, N20804, N20803, N20802, N20801, N20800, N20799, N20798, N20797, N20796, N20795, N20794, N20793, N20792, N20791, N20790, N20789, N20788, N20787, N20786, N20785, N20784, N20783, N20782, N20781, N20780, N20779, N20778, N20777, N20776, N20775, N20774, N20773, N20772, N20771, N20770, N20769, N20768, N20767, N20766, N20765, N20764, N20763, N20762, N20761, N20760, N20759, N20758, N20757, N20756, N20755, N20754, N20753, N20752, N20751, N20750, N20749, N20748, N20747, N20746, N20745, N20744, N20743, N20742, N20741, N20740, N20739, N20738, N20737, N20736, N20735, N20734, N20733, N20732, N20731, N20730, N20729, N20728, N20727, N20726, N20725, N20724, N20723, N20722, N20721, N20720, N20719, N20718, N20717, N20716, N20715, N20714, N20713, N20712, N20711, N20710, N20709, N20708, N20707, N20706, N20705, N20704, N20703, N20702, N20701, N20700, N20699, N20698, N20697, N20696, N20695, N20694, N20693, N20692, N20691, N20690, N20689, N20688, N20687, N20686, N20685, N20684, N20683, N20682, N20681, N20680, N20679, N20678, N20677, N20676, N20675, N20674, N20673, N20672, N20671, N20670, N20669, N20668, N20667, N20666, N20665, N20664, N20663, N20662, N20661, N20660, N20659, N20658, N20657, N20656, N20655, N20654, N20653, N20652, N20651, N20650, N20649, N20648, N20647, N20646, N20645, N20644, N20643, N20642, N20641, N20640, N20639, N20638, N20637, N20636, N20635, N20634, N20633, N20632, N20631, N20630, N20629, N20628, N20627, N20626, N20625, N20624, N20623, N20622, N20621, N20620, N20619, N20618, N20617, N20616, N20615, N20614, N20613, N20612, N20611, N20610, N20609, N20608, N20607, N20606, N20605, N20604, N20603, N20602, N20601, N20600, N20599, N20598, N20597, N20596, N20595, N20594, N20593, N20592, N20591, N20590, N20589, N20588, N20587, N20586, N20585, N20584, N20583, N20582, N20581, N20580, N20579, N20578, N20577, N20576, N20575, N20574, N20573, N20572, N20571, N20570, N20569, N20568, N20567, N20566, N20565, N20564, N20563, N20562, N20561, N20560, N20559, N20558, N20557, N20556, N20555, N20554, N20553, N20552, N20551, N20550, N20549, N20548, N20547, N20546, N20545, N20544, N20543, N20542, N20541, N20540, N20539, N20538, N20537, N20536, N20535, N20534, N20533, N20532, N20531, N20530, N20529, N20528, N20527, N20526, N20525, N20524, N20523, N20522, N20521, N20520, N20519, N20518, N20517, N20516, N20515, N20514, N20513, N20512, N20511, N20510, N20509, N20508, N20507, N20506, N20505, N20504, N20503, N20502, N20501, N20500, N20499, N20498, N20497, N20496, N20495, N20494, N20493, N20492, N20491, N20490, N20489, N20488, N20487, N20486, N20485, N20484, N20483, N20482, N20481, N20480, N20479, N20478, N20477, N20476, N20475, N20474, N20473, N20472, N20471 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N190)? { N18290, N18289, N18288, N18287, N18286, N18285, N18284, N18283, N18282, N18281, N18280, N18279, N18278, N18277, N18276, N18275, N18274, N18273, N18272, N18271, N18270, N18269, N18268, N18267, N18266, N18265, N18264, N18263, N18262, N18261, N18260, N18259, N18258, N18257, N18256, N18255, N18254, N18253, N18252, N18251, N18250, N18249, N18248, N18247, N18246, N18245, N18244, N18243, N18242, N18241, N18240, N18239, N18238, N18237, N18236, N18235, N18234, N18233, N18232, N18231, N18230, N18229, N18228, N18227, N18032, N18031, N18030, N18029, N18028, N18027, N18026, N18025, N18024, N18023, N18022, N18021, N18020, N18019, N18018, N18017, N18016, N18015, N18014, N18013, N18012, N18011, N18010, N18009, N18008, N18007, N18006, N18005, N18004, N18003, N18002, N18001, N18000, N17999, N17998, N17997, N17996, N17995, N17994, N17993, N17992, N17991, N17990, N17989, N17988, N17987, N17986, N17985, N17984, N17983, N17982, N17981, N17980, N17979, N17978, N17977, N17976, N17975, N17974, N17973, N17972, N17971, N17970, N17969, N17774, N17773, N17772, N17771, N17770, N17769, N17768, N17767, N17766, N17765, N17764, N17763, N17762, N17761, N17760, N17759, N17758, N17757, N17756, N17755, N17754, N17753, N17752, N17751, N17750, N17749, N17748, N17747, N17746, N17745, N17744, N17743, N17742, N17741, N17740, N17739, N17738, N17737, N17736, N17735, N17734, N17733, N17732, N17731, N17730, N17729, N17728, N17727, N17726, N17725, N17724, N17723, N17722, N17721, N17720, N17719, N17718, N17717, N17716, N17715, N17714, N17713, N17712, N17711, N17516, N17515, N17514, N17513, N17512, N17511, N17510, N17509, N17508, N17507, N17506, N17505, N17504, N17503, N17502, N17501, N17500, N17499, N17498, N17497, N17496, N17495, N17494, N17493, N17492, N17491, N17490, N17489, N17488, N17487, N17486, N17485, N17484, N17483, N17482, N17481, N17480, N17479, N17478, N17477, N17476, N17475, N17474, N17473, N17472, N17471, N17470, N17469, N17468, N17467, N17466, N17465, N17464, N17463, N17462, N17461, N17460, N17459, N17458, N17457, N17456, N17455, N17454, N17453, N17258, N17257, N17256, N17255, N17254, N17253, N17252, N17251, N17250, N17249, N17248, N17247, N17246, N17245, N17244, N17243, N17242, N17241, N17240, N17239, N17238, N17237, N17236, N17235, N17234, N17233, N17232, N17231, N17230, N17229, N17228, N17227, N17226, N17225, N17224, N17223, N17222, N17221, N17220, N17219, N17218, N17217, N17216, N17215, N17214, N17213, N17212, N17211, N17210, N17209, N17208, N17207, N17206, N17205, N17204, N17203, N17202, N17201, N17200, N17199, N17198, N17197, N17196, N17195, N17000, N16999, N16998, N16997, N16996, N16995, N16994, N16993, N16992, N16991, N16990, N16989, N16988, N16987, N16986, N16985, N16984, N16983, N16982, N16981, N16980, N16979, N16978, N16977, N16976, N16975, N16974, N16973, N16972, N16971, N16970, N16969, N16968, N16967, N16966, N16965, N16964, N16963, N16962, N16961, N16960, N16959, N16958, N16957, N16956, N16955, N16954, N16953, N16952, N16951, N16950, N16949, N16948, N16947, N16946, N16945, N16944, N16943, N16942, N16941, N16940, N16939, N16938, N16937, N16742, N16741, N16740, N16739, N16738, N16737, N16736, N16735, N16734, N16733, N16732, N16731, N16730, N16729, N16728, N16727, N16726, N16725, N16724, N16723, N16722, N16721, N16720, N16719, N16718, N16717, N16716, N16715, N16714, N16713, N16712, N16711, N16710, N16709, N16708, N16707, N16706, N16705, N16704, N16703, N16702, N16701, N16700, N16699, N16698, N16697, N16696, N16695, N16694, N16693, N16692, N16691, N16690, N16689, N16688, N16687, N16686, N16685, N16684, N16683, N16682, N16681, N16680, N16679, N16484, N16483, N16482, N16481, N16480, N16479, N16478, N16477, N16476, N16475, N16474, N16473, N16472, N16471, N16470, N16469, N16468, N16467, N16466, N16465, N16464, N16463, N16462, N16461, N16460, N16459, N16458, N16457, N16456, N16455, N16454, N16453, N16452, N16451, N16450, N16449, N16448, N16447, N16446, N16445, N16444, N16443, N16442, N16441, N16440, N16439, N16438, N16437, N16436, N16435, N16434, N16433, N16432, N16431, N16430, N16429, N16428, N16427, N16426, N16425, N16424, N16423, N16422, N16421 } : 1'b0;
  assign N189 = N20469;
  assign N190 = N20470;
  assign { N22526, N22525, N22524, N22523, N22522, N22521, N22520, N22519, N22518, N22517, N22516, N22515, N22514, N22513, N22512, N22511, N22510, N22509, N22508, N22507, N22506, N22505, N22504, N22503, N22502, N22501, N22500, N22499, N22498, N22497, N22496, N22495, N22494, N22493, N22492, N22491, N22490, N22489, N22488, N22487, N22486, N22485, N22484, N22483, N22482, N22481, N22480, N22479, N22478, N22477, N22476, N22475, N22474, N22473, N22472, N22471, N22470, N22469, N22468, N22467, N22466, N22465, N22464, N22463, N22462, N22461, N22460, N22459, N22458, N22457, N22456, N22455, N22454, N22453, N22452, N22451, N22450, N22449, N22448, N22447, N22446, N22445, N22444, N22443, N22442, N22441, N22440, N22439, N22438, N22437, N22436, N22435, N22434, N22433, N22432, N22431, N22430, N22429, N22428, N22427, N22426, N22425, N22424, N22423, N22422, N22421, N22420, N22419, N22418, N22417, N22416, N22415, N22414, N22413, N22412, N22411, N22410, N22409, N22408, N22407, N22406, N22405, N22404, N22403, N22402, N22401, N22400, N22399, N22398, N22397, N22396, N22395, N22394, N22393, N22392, N22391, N22390, N22389, N22388, N22387, N22386, N22385, N22384, N22383, N22382, N22381, N22380, N22379, N22378, N22377, N22376, N22375, N22374, N22373, N22372, N22371, N22370, N22369, N22368, N22367, N22366, N22365, N22364, N22363, N22362, N22361, N22360, N22359, N22358, N22357, N22356, N22355, N22354, N22353, N22352, N22351, N22350, N22349, N22348, N22347, N22346, N22345, N22344, N22343, N22342, N22341, N22340, N22339, N22338, N22337, N22336, N22335, N22334, N22333, N22332, N22331, N22330, N22329, N22328, N22327, N22326, N22325, N22324, N22323, N22322, N22321, N22320, N22319, N22318, N22317, N22316, N22315, N22314, N22313, N22312, N22311, N22310, N22309, N22308, N22307, N22306, N22305, N22304, N22303, N22302, N22301, N22300, N22299, N22298, N22297, N22296, N22295, N22294, N22293, N22292, N22291, N22290, N22289, N22288, N22287, N22286, N22285, N22284, N22283, N22282, N22281, N22280, N22279, N22278, N22277, N22276, N22275, N22274, N22273, N22272, N22271, N22270, N22269, N22268, N22267, N22266, N22265, N22264, N22263, N22262, N22261, N22260, N22259, N22258, N22257, N22256, N22255, N22254, N22253, N22252, N22251, N22250, N22249, N22248, N22247, N22246, N22245, N22244, N22243, N22242, N22241, N22240, N22239, N22238, N22237, N22236, N22235, N22234, N22233, N22232, N22231, N22230, N22229, N22228, N22227, N22226, N22225, N22224, N22223, N22222, N22221, N22220, N22219, N22218, N22217, N22216, N22215, N22214, N22213, N22212, N22211, N22210, N22209, N22208, N22207, N22206, N22205, N22204, N22203, N22202, N22201, N22200, N22199, N22198, N22197, N22196, N22195, N22194, N22193, N22192, N22191, N22190, N22189, N22188, N22187, N22186, N22185, N22184, N22183, N22182, N22181, N22180, N22179, N22178, N22177, N22176, N22175, N22174, N22173, N22172, N22171, N22170, N22169, N22168, N22167, N22166, N22165, N22164, N22163, N22162, N22161, N22160, N22159, N22158, N22157, N22156, N22155, N22154, N22153, N22152, N22151, N22150, N22149, N22148, N22147, N22146, N22145, N22144, N22143, N22142, N22141, N22140, N22139, N22138, N22137, N22136, N22135, N22134, N22133, N22132, N22131, N22130, N22129, N22128, N22127, N22126, N22125, N22124, N22123, N22122, N22121, N22120, N22119, N22118, N22117, N22116, N22115, N22114, N22113, N22112, N22111, N22110, N22109, N22108, N22107, N22106, N22105, N22104, N22103, N22102, N22101, N22100, N22099, N22098, N22097, N22096, N22095, N22094, N22093, N22092, N22091, N22090, N22089, N22088, N22087, N22086, N22085, N22084, N22083, N22082, N22081, N22080, N22079, N22078, N22077, N22076, N22075, N22074, N22073, N22072, N22071, N22070, N22069, N22068, N22067, N22066, N22065, N22064, N22063, N22062, N22061, N22060, N22059, N22058, N22057, N22056, N22055, N22054, N22053, N22052, N22051, N22050, N22049, N22048, N22047, N22046, N22045, N22044, N22043, N22042, N22041, N22040, N22039, N22038, N22037, N22036, N22035, N22034, N22033, N22032, N22031, N22030, N22029, N22028, N22027, N22026, N22025, N22024, N22023, N22022, N22021, N22020, N22019, N22018, N22017, N22016, N22015, N22014, N22013, N22012, N22011, N22010, N22009, N22008, N22007, N22006, N22005, N22004, N22003, N22002, N22001, N22000, N21999, N21998, N21997, N21996, N21995, N21994, N21993, N21992, N21991, N21990, N21989, N21988, N21987, N21986, N21985, N21984, N21983, N21982, N21981, N21980, N21979, N21978, N21977, N21976, N21975, N21974, N21973, N21972, N21971, N21970, N21969, N21968, N21967, N21966, N21965, N21964, N21963, N21962, N21961, N21960, N21959, N21958, N21957, N21956, N21955, N21954, N21953, N21952, N21951, N21950, N21949, N21948, N21947, N21946, N21945, N21944, N21943, N21942, N21941, N21940, N21939, N21938, N21937, N21936, N21935, N21934, N21933, N21932, N21931, N21930, N21929, N21928, N21927, N21926, N21925, N21924, N21923, N21922, N21921, N21920, N21919, N21918, N21917, N21916, N21915, N21914, N21913, N21912, N21911, N21910, N21909, N21908, N21907, N21906, N21905, N21904, N21903, N21902, N21901, N21900, N21899, N21898, N21897, N21896, N21895, N21894, N21893, N21892, N21891, N21890, N21889, N21888, N21887, N21886, N21885, N21884, N21883, N21882, N21881, N21880, N21879, N21878, N21877, N21876, N21875, N21874, N21873, N21872, N21871, N21870, N21869, N21868, N21867, N21866, N21865, N21864, N21863, N21862, N21861, N21860, N21859, N21858, N21857, N21856, N21855, N21854, N21853, N21852, N21851, N21850, N21849, N21848, N21847, N21846, N21845, N21844, N21843, N21842, N21841, N21840, N21839, N21838, N21837, N21836, N21835, N21834, N21833, N21832, N21831, N21830, N21829, N21828, N21827, N21826, N21825, N21824, N21823, N21822, N21821, N21820, N21819, N21818, N21817, N21816, N21815, N21814, N21813, N21812, N21811, N21810, N21809, N21808, N21807, N21806, N21805, N21804, N21803, N21802, N21801, N21800, N21799, N21798, N21797, N21796, N21795, N21794, N21793, N21792, N21791, N21790, N21789, N21788, N21787, N21786, N21785, N21784, N21783, N21782, N21781, N21780, N21779, N21778, N21777, N21776, N21775, N21774, N21773, N21772, N21771, N21770, N21769, N21768, N21767, N21766, N21765, N21764, N21763, N21762, N21761, N21760, N21759, N21758, N21757, N21756, N21755, N21754, N21753, N21752, N21751, N21750, N21749, N21748, N21747, N21746, N21745, N21744, N21743, N21742, N21741, N21740, N21739, N21738, N21737, N21736, N21735, N21734, N21733, N21732, N21731, N21730, N21729, N21728, N21727, N21726, N21725, N21724, N21723, N21722, N21721, N21720, N21719, N21718, N21717, N21716, N21715, N21714, N21713, N21712, N21711, N21710, N21709, N21708, N21707, N21706, N21705, N21704, N21703, N21702, N21701, N21700, N21699, N21698, N21697, N21696, N21695, N21694, N21693, N21692, N21691, N21690, N21689, N21688, N21687, N21686, N21685, N21684, N21683, N21682, N21681, N21680, N21679, N21678, N21677, N21676, N21675, N21674, N21673, N21672, N21671, N21670, N21669, N21668, N21667, N21666, N21665, N21664, N21663, N21662, N21661, N21660, N21659, N21658, N21657, N21656, N21655, N21654, N21653, N21652, N21651, N21650, N21649, N21648, N21647, N21646, N21645, N21644, N21643, N21642, N21641, N21640, N21639, N21638, N21637, N21636, N21635, N21634, N21633, N21632, N21631, N21630, N21629, N21628, N21627, N21626, N21625, N21624, N21623, N21622, N21621, N21620, N21619, N21618, N21617, N21616, N21615, N21614, N21613, N21612, N21611, N21610, N21609, N21608, N21607, N21606, N21605, N21604, N21603, N21602, N21601, N21600, N21599, N21598, N21597, N21596, N21595, N21594, N21593, N21592, N21591, N21590, N21589, N21588, N21587, N21586, N21585, N21584, N21583, N21582, N21581, N21580, N21579, N21578, N21577, N21576, N21575, N21574, N21573, N21572, N21571, N21570, N21569, N21568, N21567, N21566, N21565, N21564, N21563, N21562, N21561, N21560, N21559, N21558, N21557, N21556, N21555, N21554, N21553, N21552, N21551, N21550, N21549, N21548, N21547, N21546, N21545, N21544, N21543, N21542, N21541, N21540, N21539, N21538, N21537, N21536, N21535, N21534, N21533, N21532, N21531, N21530, N21529, N21528, N21527, N21526, N21525, N21524, N21523, N21522, N21521, N21520, N21519, N21518, N21517, N21516, N21515, N21514, N21513, N21512, N21511, N21510, N21509, N21508, N21507, N21506, N21505, N21504, N21503, N21502, N21501, N21500, N21499, N21498, N21497, N21496, N21495 } = (N191)? { N20458, N20457, N20456, N20455, N20454, N20453, N20452, N20451, N20450, N20449, N20448, N20447, N20446, N20445, N20444, N20443, N20442, N20441, N20440, N20439, N20438, N20437, N20436, N20435, N20434, N20433, N20432, N20431, N20430, N20429, N20428, N20427, N20426, N20425, N20424, N20423, N20422, N20421, N20420, N20419, N20418, N20417, N20416, N20415, N20414, N20413, N20412, N20411, N20410, N20409, N20408, N20407, N20406, N20405, N20404, N20403, N20402, N20401, N20400, N20399, N20398, N20397, N20396, N20395, N20394, N20393, N20392, N20391, N20390, N20389, N20388, N20387, N20386, N20385, N20384, N20383, N20382, N20381, N20380, N20379, N20378, N20377, N20376, N20375, N20374, N20373, N20372, N20371, N20370, N20369, N20368, N20367, N20366, N20365, N20364, N20363, N20362, N20361, N20360, N20359, N20358, N20357, N20356, N20355, N20354, N20353, N20352, N20351, N20350, N20349, N20348, N20347, N20346, N20345, N20344, N20343, N20342, N20341, N20340, N20339, N20338, N20337, N20336, N20335, N20334, N20333, N20332, N20331, N20330, N20329, N20328, N20327, N20326, N20325, N20324, N20323, N20322, N20321, N20320, N20319, N20318, N20317, N20316, N20315, N20314, N20313, N20312, N20311, N20310, N20309, N20308, N20307, N20306, N20305, N20304, N20303, N20302, N20301, N20300, N20299, N20298, N20297, N20296, N20295, N20294, N20293, N20292, N20291, N20290, N20289, N20288, N20287, N20286, N20285, N20284, N20283, N20282, N20281, N20280, N20279, N20278, N20277, N20276, N20275, N20274, N20273, N20272, N20271, N20270, N20269, N20268, N20267, N20266, N20265, N20264, N20263, N20262, N20261, N20260, N20259, N20258, N20257, N20256, N20255, N20254, N20253, N20252, N20251, N20250, N20249, N20248, N20247, N20246, N20245, N20244, N20243, N20242, N20241, N20240, N20239, N20238, N20237, N20236, N20235, N20234, N20233, N20232, N20231, N20230, N20229, N20228, N20227, N20226, N20225, N20224, N20223, N20222, N20221, N20220, N20219, N20218, N20217, N20216, N20215, N20214, N20213, N20212, N20211, N20210, N20209, N20208, N20207, N20206, N20205, N20204, N20203, N20202, N20201, N20200, N20199, N20198, N20197, N20196, N20195, N20194, N20193, N20192, N20191, N20190, N20189, N20188, N20187, N20186, N20185, N20184, N20183, N20182, N20181, N20180, N20179, N20178, N20177, N20176, N20175, N20174, N20173, N20172, N20171, N20170, N20169, N20168, N20167, N20166, N20165, N20164, N20163, N20162, N20161, N20160, N20159, N20158, N20157, N20156, N20155, N20154, N20153, N20152, N20151, N20150, N20149, N20148, N20147, N20146, N20145, N20144, N20143, N20142, N20141, N20140, N20139, N20138, N20137, N20136, N20135, N20134, N20133, N20132, N20131, N20130, N20129, N20128, N20127, N20126, N20125, N20124, N20123, N20122, N20121, N20120, N20119, N20118, N20117, N20116, N20115, N20114, N20113, N20112, N20111, N20110, N20109, N20108, N20107, N20106, N20105, N20104, N20103, N20102, N20101, N20100, N20099, N20098, N20097, N20096, N20095, N20094, N20093, N20092, N20091, N20090, N20089, N20088, N20087, N20086, N20085, N20084, N20083, N20082, N20081, N20080, N20079, N20078, N20077, N20076, N20075, N20074, N20073, N20072, N20071, N20070, N20069, N20068, N20067, N20066, N20065, N20064, N20063, N20062, N20061, N20060, N20059, N20058, N20057, N20056, N20055, N20054, N20053, N20052, N20051, N20050, N20049, N20048, N20047, N20046, N20045, N20044, N20043, N20042, N20041, N20040, N20039, N20038, N20037, N20036, N20035, N20034, N20033, N20032, N20031, N20030, N20029, N20028, N20027, N20026, N20025, N20024, N20023, N20022, N20021, N20020, N20019, N20018, N20017, N20016, N20015, N20014, N20013, N20012, N20011, N20010, N20009, N20008, N20007, N20006, N20005, N20004, N20003, N20002, N20001, N20000, N19999, N19998, N19997, N19996, N19995, N19994, N19993, N19992, N19991, N19990, N19989, N19988, N19987, N19986, N19985, N19984, N19983, N19982, N19981, N19980, N19979, N19978, N19977, N19976, N19975, N19974, N19973, N19972, N19971, N19970, N19969, N19968, N19967, N19966, N19965, N19964, N19963, N19962, N19961, N19960, N19959, N19958, N19957, N19956, N19955, N19954, N19953, N19952, N19951, N19950, N19949, N19948, N19947, N19946, N19945, N19944, N19943, N19942, N19941, N19940, N19939, N19938, N19937, N19936, N19935, N19934, N19933, N19932, N19931, N19930, N19929, N19928, N19927, N19926, N19925, N19924, N19923, N19922, N19921, N19920, N19919, N19918, N19917, N19916, N19915, N19914, N19913, N19912, N19911, N19910, N19909, N19908, N19907, N19906, N19905, N19904, N19903, N19902, N19901, N19900, N19899, N19898, N19897, N19896, N19895, N19894, N19893, N19892, N19891, N19890, N19889, N19888, N19887, N19886, N19885, N19884, N19883, N19882, N19881, N19880, N19879, N19878, N19877, N19876, N19875, N19874, N19873, N19872, N19871, N19870, N19869, N19868, N19867, N19866, N19865, N19864, N19863, N19862, N19861, N19860, N19859, N19858, N19857, N19856, N19855, N19854, N19853, N19852, N19851, N19850, N19849, N19848, N19847, N19846, N19845, N19844, N19843, N19842, N19841, N19840, N19839, N19838, N19837, N19836, N19835, N19834, N19833, N19832, N19831, N19830, N19829, N19828, N19827, N19826, N19825, N19824, N19823, N19822, N19821, N19820, N19819, N19818, N19817, N19816, N19815, N19814, N19813, N19812, N19811, N19810, N19809, N19808, N19807, N19806, N19805, N19804, N19803, N19802, N19801, N19800, N19799, N19798, N19797, N19796, N19795, N19794, N19793, N19792, N19791, N19790, N19789, N19788, N19787, N19786, N19785, N19784, N19783, N19782, N19781, N19780, N19779, N19778, N19777, N19776, N19775, N19774, N19773, N19772, N19771, N19770, N19769, N19768, N19767, N19766, N19765, N19764, N19763, N19762, N19761, N19760, N19759, N19758, N19757, N19756, N19755, N19754, N19753, N19752, N19751, N19750, N19749, N19748, N19747, N19746, N19745, N19744, N19743, N19742, N19741, N19740, N19739, N19738, N19737, N19736, N19735, N19734, N19733, N19732, N19731, N19730, N19729, N19728, N19727, N19726, N19725, N19724, N19723, N19722, N19721, N19720, N19719, N19718, N19717, N19716, N19715, N19714, N19713, N19712, N19711, N19710, N19709, N19708, N19707, N19706, N19705, N19704, N19703, N19702, N19701, N19700, N19699, N19698, N19697, N19696, N19695, N19694, N19693, N19692, N19691, N19690, N19689, N19688, N19687, N19686, N19685, N19684, N19683, N19682, N19681, N19680, N19679, N19678, N19677, N19676, N19675, N19674, N19673, N19672, N19671, N19670, N19669, N19668, N19667, N19666, N19665, N19664, N19663, N19662, N19661, N19660, N19659, N19658, N19657, N19656, N19655, N19654, N19653, N19652, N19651, N19650, N19649, N19648, N19647, N19646, N19645, N19644, N19643, N19642, N19641, N19640, N19639, N19638, N19637, N19636, N19635, N19634, N19633, N19632, N19631, N19630, N19629, N19628, N19627, N19626, N19625, N19624, N19623, N19622, N19621, N19620, N19619, N19618, N19617, N19616, N19615, N19614, N19613, N19612, N19611, N19610, N19609, N19608, N19607, N19606, N19605, N19604, N19603, N19602, N19601, N19600, N19599, N19598, N19597, N19596, N19595, N19594, N19593, N19592, N19591, N19590, N19589, N19588, N19587, N19586, N19585, N19584, N19583, N19582, N19581, N19580, N19579, N19578, N19577, N19576, N19575, N19574, N19573, N19572, N19571, N19570, N19569, N19568, N19567, N19566, N19565, N19564, N19563, N19562, N19561, N19560, N19559, N19558, N19557, N19556, N19555, N19554, N19553, N19552, N19551, N19550, N19549, N19548, N19547, N19546, N19545, N19544, N19543, N19542, N19541, N19540, N19539, N19538, N19537, N19536, N19535, N19534, N19533, N19532, N19531, N19530, N19529, N19528, N19527, N19526, N19525, N19524, N19523, N19522, N19521, N19520, N19519, N19518, N19517, N19516, N19515, N19514, N19513, N19512, N19511, N19510, N19509, N19508, N19507, N19506, N19505, N19504, N19503, N19502, N19501, N19500, N19499, N19498, N19497, N19496, N19495, N19494, N19493, N19492, N19491, N19490, N19489, N19488, N19487, N19486, N19485, N19484, N19483, N19482, N19481, N19480, N19479, N19478, N19477, N19476, N19475, N19474, N19473, N19472, N19471, N19470, N19469, N19468, N19467, N19466, N19465, N19464, N19463, N19462, N19461, N19460, N19459, N19458, N19457, N19456, N19455, N19454, N19453, N19452, N19451, N19450, N19449, N19448, N19447, N19446, N19445, N19444, N19443, N19442, N19441, N19440, N19439, N19438, N19437, N19436, N19435, N19434, N19433, N19432, N19431, N19430, N19429, N19428, N19427 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N19426)? { N21494, N21493, N21492, N21491, N21490, N21489, N21488, N21487, N21486, N21485, N21484, N21483, N21482, N21481, N21480, N21479, N21478, N21477, N21476, N21475, N21474, N21473, N21472, N21471, N21470, N21469, N21468, N21467, N21466, N21465, N21464, N21463, N21462, N21461, N21460, N21459, N21458, N21457, N21456, N21455, N21454, N21453, N21452, N21451, N21450, N21449, N21448, N21447, N21446, N21445, N21444, N21443, N21442, N21441, N21440, N21439, N21438, N21437, N21436, N21435, N21434, N21433, N21432, N21431, N18226, N18225, N18224, N18223, N18222, N18221, N18220, N18219, N18218, N18217, N18216, N18215, N18214, N18213, N18212, N18211, N18210, N18209, N18208, N18207, N18206, N18205, N18204, N18203, N18202, N18201, N18200, N18199, N18198, N18197, N18196, N18195, N18194, N18193, N18192, N18191, N18190, N18189, N18188, N18187, N18186, N18185, N18184, N18183, N18182, N18181, N18180, N18179, N18178, N18177, N18176, N18175, N18174, N18173, N18172, N18171, N18170, N18169, N18168, N18167, N18166, N18165, N18164, N18163, N18162, N21430, N21429, N21428, N21427, N21426, N21425, N21424, N21423, N21422, N21421, N21420, N21419, N21418, N21417, N21416, N21415, N21414, N21413, N21412, N21411, N21410, N21409, N21408, N21407, N21406, N21405, N21404, N21403, N21402, N21401, N21400, N21399, N21398, N21397, N21396, N21395, N21394, N21393, N21392, N21391, N21390, N21389, N21388, N21387, N21386, N21385, N21384, N21383, N21382, N21381, N21380, N21379, N21378, N21377, N21376, N21375, N21374, N21373, N21372, N21371, N21370, N21369, N21368, N21367, N17968, N17967, N17966, N17965, N17964, N17963, N17962, N17961, N17960, N17959, N17958, N17957, N17956, N17955, N17954, N17953, N17952, N17951, N17950, N17949, N17948, N17947, N17946, N17945, N17944, N17943, N17942, N17941, N17940, N17939, N17938, N17937, N17936, N17935, N17934, N17933, N17932, N17931, N17930, N17929, N17928, N17927, N17926, N17925, N17924, N17923, N17922, N17921, N17920, N17919, N17918, N17917, N17916, N17915, N17914, N17913, N17912, N17911, N17910, N17909, N17908, N17907, N17906, N17905, N17904, N21366, N21365, N21364, N21363, N21362, N21361, N21360, N21359, N21358, N21357, N21356, N21355, N21354, N21353, N21352, N21351, N21350, N21349, N21348, N21347, N21346, N21345, N21344, N21343, N21342, N21341, N21340, N21339, N21338, N21337, N21336, N21335, N21334, N21333, N21332, N21331, N21330, N21329, N21328, N21327, N21326, N21325, N21324, N21323, N21322, N21321, N21320, N21319, N21318, N21317, N21316, N21315, N21314, N21313, N21312, N21311, N21310, N21309, N21308, N21307, N21306, N21305, N21304, N21303, N17710, N17709, N17708, N17707, N17706, N17705, N17704, N17703, N17702, N17701, N17700, N17699, N17698, N17697, N17696, N17695, N17694, N17693, N17692, N17691, N17690, N17689, N17688, N17687, N17686, N17685, N17684, N17683, N17682, N17681, N17680, N17679, N17678, N17677, N17676, N17675, N17674, N17673, N17672, N17671, N17670, N17669, N17668, N17667, N17666, N17665, N17664, N17663, N17662, N17661, N17660, N17659, N17658, N17657, N17656, N17655, N17654, N17653, N17652, N17651, N17650, N17649, N17648, N17647, N17646, N21302, N21301, N21300, N21299, N21298, N21297, N21296, N21295, N21294, N21293, N21292, N21291, N21290, N21289, N21288, N21287, N21286, N21285, N21284, N21283, N21282, N21281, N21280, N21279, N21278, N21277, N21276, N21275, N21274, N21273, N21272, N21271, N21270, N21269, N21268, N21267, N21266, N21265, N21264, N21263, N21262, N21261, N21260, N21259, N21258, N21257, N21256, N21255, N21254, N21253, N21252, N21251, N21250, N21249, N21248, N21247, N21246, N21245, N21244, N21243, N21242, N21241, N21240, N21239, N17452, N17451, N17450, N17449, N17448, N17447, N17446, N17445, N17444, N17443, N17442, N17441, N17440, N17439, N17438, N17437, N17436, N17435, N17434, N17433, N17432, N17431, N17430, N17429, N17428, N17427, N17426, N17425, N17424, N17423, N17422, N17421, N17420, N17419, N17418, N17417, N17416, N17415, N17414, N17413, N17412, N17411, N17410, N17409, N17408, N17407, N17406, N17405, N17404, N17403, N17402, N17401, N17400, N17399, N17398, N17397, N17396, N17395, N17394, N17393, N17392, N17391, N17390, N17389, N17388, N21238, N21237, N21236, N21235, N21234, N21233, N21232, N21231, N21230, N21229, N21228, N21227, N21226, N21225, N21224, N21223, N21222, N21221, N21220, N21219, N21218, N21217, N21216, N21215, N21214, N21213, N21212, N21211, N21210, N21209, N21208, N21207, N21206, N21205, N21204, N21203, N21202, N21201, N21200, N21199, N21198, N21197, N21196, N21195, N21194, N21193, N21192, N21191, N21190, N21189, N21188, N21187, N21186, N21185, N21184, N21183, N21182, N21181, N21180, N21179, N21178, N21177, N21176, N21175, N17194, N17193, N17192, N17191, N17190, N17189, N17188, N17187, N17186, N17185, N17184, N17183, N17182, N17181, N17180, N17179, N17178, N17177, N17176, N17175, N17174, N17173, N17172, N17171, N17170, N17169, N17168, N17167, N17166, N17165, N17164, N17163, N17162, N17161, N17160, N17159, N17158, N17157, N17156, N17155, N17154, N17153, N17152, N17151, N17150, N17149, N17148, N17147, N17146, N17145, N17144, N17143, N17142, N17141, N17140, N17139, N17138, N17137, N17136, N17135, N17134, N17133, N17132, N17131, N17130, N21174, N21173, N21172, N21171, N21170, N21169, N21168, N21167, N21166, N21165, N21164, N21163, N21162, N21161, N21160, N21159, N21158, N21157, N21156, N21155, N21154, N21153, N21152, N21151, N21150, N21149, N21148, N21147, N21146, N21145, N21144, N21143, N21142, N21141, N21140, N21139, N21138, N21137, N21136, N21135, N21134, N21133, N21132, N21131, N21130, N21129, N21128, N21127, N21126, N21125, N21124, N21123, N21122, N21121, N21120, N21119, N21118, N21117, N21116, N21115, N21114, N21113, N21112, N21111, N16936, N16935, N16934, N16933, N16932, N16931, N16930, N16929, N16928, N16927, N16926, N16925, N16924, N16923, N16922, N16921, N16920, N16919, N16918, N16917, N16916, N16915, N16914, N16913, N16912, N16911, N16910, N16909, N16908, N16907, N16906, N16905, N16904, N16903, N16902, N16901, N16900, N16899, N16898, N16897, N16896, N16895, N16894, N16893, N16892, N16891, N16890, N16889, N16888, N16887, N16886, N16885, N16884, N16883, N16882, N16881, N16880, N16879, N16878, N16877, N16876, N16875, N16874, N16873, N16872, N21110, N21109, N21108, N21107, N21106, N21105, N21104, N21103, N21102, N21101, N21100, N21099, N21098, N21097, N21096, N21095, N21094, N21093, N21092, N21091, N21090, N21089, N21088, N21087, N21086, N21085, N21084, N21083, N21082, N21081, N21080, N21079, N21078, N21077, N21076, N21075, N21074, N21073, N21072, N21071, N21070, N21069, N21068, N21067, N21066, N21065, N21064, N21063, N21062, N21061, N21060, N21059, N21058, N21057, N21056, N21055, N21054, N21053, N21052, N21051, N21050, N21049, N21048, N21047, N16678, N16677, N16676, N16675, N16674, N16673, N16672, N16671, N16670, N16669, N16668, N16667, N16666, N16665, N16664, N16663, N16662, N16661, N16660, N16659, N16658, N16657, N16656, N16655, N16654, N16653, N16652, N16651, N16650, N16649, N16648, N16647, N16646, N16645, N16644, N16643, N16642, N16641, N16640, N16639, N16638, N16637, N16636, N16635, N16634, N16633, N16632, N16631, N16630, N16629, N16628, N16627, N16626, N16625, N16624, N16623, N16622, N16621, N16620, N16619, N16618, N16617, N16616, N16615, N16614, N21046, N21045, N21044, N21043, N21042, N21041, N21040, N21039, N21038, N21037, N21036, N21035, N21034, N21033, N21032, N21031, N21030, N21029, N21028, N21027, N21026, N21025, N21024, N21023, N21022, N21021, N21020, N21019, N21018, N21017, N21016, N21015, N21014, N21013, N21012, N21011, N21010, N21009, N21008, N21007, N21006, N21005, N21004, N21003, N21002, N21001, N21000, N20999, N20998, N20997, N20996, N20995, N20994, N20993, N20992, N20991, N20990, N20989, N20988, N20987, N20986, N20985, N20984, N20983, N16420, N16419, N16418, N16417, N16416, N16415, N16414, N16413, N16412, N16411, N16410, N16409, N16408, N16407, N16406, N16405, N16404, N16403, N16402, N16401, N16400, N16399, N16398, N16397, N16396, N16395, N16394, N16393, N16392, N16391, N16390, N16389, N16388, N16387, N16386, N16385, N16384, N16383, N16382, N16381, N16380, N16379, N16378, N16377, N16376, N16375, N16374, N16373, N16372, N16371, N16370, N16369, N16368, N16367, N16366, N16365, N16364, N16363, N16362, N16361, N16360, N16359, N16358, N16357, N16356 } : 1'b0;
  assign N191 = ex_i[258];
  assign { N24590, N24589, N24588, N24587, N24586, N24585, N24584, N24583, N24582, N24581, N24580, N24579, N24578, N24577, N24576, N24575, N24574, N24573, N24572, N24571, N24570, N24569, N24568, N24567, N24566, N24565, N24564, N24563, N24562, N24561, N24560, N24559, N24558, N24557, N24556, N24555, N24554, N24553, N24552, N24551, N24550, N24549, N24548, N24547, N24546, N24545, N24544, N24543, N24542, N24541, N24540, N24539, N24538, N24537, N24536, N24535, N24534, N24533, N24532, N24531, N24530, N24529, N24528, N24527, N24526, N24525, N24524, N24523, N24522, N24521, N24520, N24519, N24518, N24517, N24516, N24515, N24514, N24513, N24512, N24511, N24510, N24509, N24508, N24507, N24506, N24505, N24504, N24503, N24502, N24501, N24500, N24499, N24498, N24497, N24496, N24495, N24494, N24493, N24492, N24491, N24490, N24489, N24488, N24487, N24486, N24485, N24484, N24483, N24482, N24481, N24480, N24479, N24478, N24477, N24476, N24475, N24474, N24473, N24472, N24471, N24470, N24469, N24468, N24467, N24466, N24465, N24464, N24463, N24462, N24461, N24460, N24459, N24458, N24457, N24456, N24455, N24454, N24453, N24452, N24451, N24450, N24449, N24448, N24447, N24446, N24445, N24444, N24443, N24442, N24441, N24440, N24439, N24438, N24437, N24436, N24435, N24434, N24433, N24432, N24431, N24430, N24429, N24428, N24427, N24426, N24425, N24424, N24423, N24422, N24421, N24420, N24419, N24418, N24417, N24416, N24415, N24414, N24413, N24412, N24411, N24410, N24409, N24408, N24407, N24406, N24405, N24404, N24403, N24402, N24401, N24400, N24399, N24398, N24397, N24396, N24395, N24394, N24393, N24392, N24391, N24390, N24389, N24388, N24387, N24386, N24385, N24384, N24383, N24382, N24381, N24380, N24379, N24378, N24377, N24376, N24375, N24374, N24373, N24372, N24371, N24370, N24369, N24368, N24367, N24366, N24365, N24364, N24363, N24362, N24361, N24360, N24359, N24358, N24357, N24356, N24355, N24354, N24353, N24352, N24351, N24350, N24349, N24348, N24347, N24346, N24345, N24344, N24343, N24342, N24341, N24340, N24339, N24338, N24337, N24336, N24335, N24334, N24333, N24332, N24331, N24330, N24329, N24328, N24327, N24326, N24325, N24324, N24323, N24322, N24321, N24320, N24319, N24318, N24317, N24316, N24315, N24314, N24313, N24312, N24311, N24310, N24309, N24308, N24307, N24306, N24305, N24304, N24303, N24302, N24301, N24300, N24299, N24298, N24297, N24296, N24295, N24294, N24293, N24292, N24291, N24290, N24289, N24288, N24287, N24286, N24285, N24284, N24283, N24282, N24281, N24280, N24279, N24278, N24277, N24276, N24275, N24274, N24273, N24272, N24271, N24270, N24269, N24268, N24267, N24266, N24265, N24264, N24263, N24262, N24261, N24260, N24259, N24258, N24257, N24256, N24255, N24254, N24253, N24252, N24251, N24250, N24249, N24248, N24247, N24246, N24245, N24244, N24243, N24242, N24241, N24240, N24239, N24238, N24237, N24236, N24235, N24234, N24233, N24232, N24231, N24230, N24229, N24228, N24227, N24226, N24225, N24224, N24223, N24222, N24221, N24220, N24219, N24218, N24217, N24216, N24215, N24214, N24213, N24212, N24211, N24210, N24209, N24208, N24207, N24206, N24205, N24204, N24203, N24202, N24201, N24200, N24199, N24198, N24197, N24196, N24195, N24194, N24193, N24192, N24191, N24190, N24189, N24188, N24187, N24186, N24185, N24184, N24183, N24182, N24181, N24180, N24179, N24178, N24177, N24176, N24175, N24174, N24173, N24172, N24171, N24170, N24169, N24168, N24167, N24166, N24165, N24164, N24163, N24162, N24161, N24160, N24159, N24158, N24157, N24156, N24155, N24154, N24153, N24152, N24151, N24150, N24149, N24148, N24147, N24146, N24145, N24144, N24143, N24142, N24141, N24140, N24139, N24138, N24137, N24136, N24135, N24134, N24133, N24132, N24131, N24130, N24129, N24128, N24127, N24126, N24125, N24124, N24123, N24122, N24121, N24120, N24119, N24118, N24117, N24116, N24115, N24114, N24113, N24112, N24111, N24110, N24109, N24108, N24107, N24106, N24105, N24104, N24103, N24102, N24101, N24100, N24099, N24098, N24097, N24096, N24095, N24094, N24093, N24092, N24091, N24090, N24089, N24088, N24087, N24086, N24085, N24084, N24083, N24082, N24081, N24080, N24079, N24078, N24077, N24076, N24075, N24074, N24073, N24072, N24071, N24070, N24069, N24068, N24067, N24066, N24065, N24064, N24063, N24062, N24061, N24060, N24059, N24058, N24057, N24056, N24055, N24054, N24053, N24052, N24051, N24050, N24049, N24048, N24047, N24046, N24045, N24044, N24043, N24042, N24041, N24040, N24039, N24038, N24037, N24036, N24035, N24034, N24033, N24032, N24031, N24030, N24029, N24028, N24027, N24026, N24025, N24024, N24023, N24022, N24021, N24020, N24019, N24018, N24017, N24016, N24015, N24014, N24013, N24012, N24011, N24010, N24009, N24008, N24007, N24006, N24005, N24004, N24003, N24002, N24001, N24000, N23999, N23998, N23997, N23996, N23995, N23994, N23993, N23992, N23991, N23990, N23989, N23988, N23987, N23986, N23985, N23984, N23983, N23982, N23981, N23980, N23979, N23978, N23977, N23976, N23975, N23974, N23973, N23972, N23971, N23970, N23969, N23968, N23967, N23966, N23965, N23964, N23963, N23962, N23961, N23960, N23959, N23958, N23957, N23956, N23955, N23954, N23953, N23952, N23951, N23950, N23949, N23948, N23947, N23946, N23945, N23944, N23943, N23942, N23941, N23940, N23939, N23938, N23937, N23936, N23935, N23934, N23933, N23932, N23931, N23930, N23929, N23928, N23927, N23926, N23925, N23924, N23923, N23922, N23921, N23920, N23919, N23918, N23917, N23916, N23915, N23914, N23913, N23912, N23911, N23910, N23909, N23908, N23907, N23906, N23905, N23904, N23903, N23902, N23901, N23900, N23899, N23898, N23897, N23896, N23895, N23894, N23893, N23892, N23891, N23890, N23889, N23888, N23887, N23886, N23885, N23884, N23883, N23882, N23881, N23880, N23879, N23878, N23877, N23876, N23875, N23874, N23873, N23872, N23871, N23870, N23869, N23868, N23867, N23866, N23865, N23864, N23863, N23862, N23861, N23860, N23859, N23858, N23857, N23856, N23855, N23854, N23853, N23852, N23851, N23850, N23849, N23848, N23847, N23846, N23845, N23844, N23843, N23842, N23841, N23840, N23839, N23838, N23837, N23836, N23835, N23834, N23833, N23832, N23831, N23830, N23829, N23828, N23827, N23826, N23825, N23824, N23823, N23822, N23821, N23820, N23819, N23818, N23817, N23816, N23815, N23814, N23813, N23812, N23811, N23810, N23809, N23808, N23807, N23806, N23805, N23804, N23803, N23802, N23801, N23800, N23799, N23798, N23797, N23796, N23795, N23794, N23793, N23792, N23791, N23790, N23789, N23788, N23787, N23786, N23785, N23784, N23783, N23782, N23781, N23780, N23779, N23778, N23777, N23776, N23775, N23774, N23773, N23772, N23771, N23770, N23769, N23768, N23767, N23766, N23765, N23764, N23763, N23762, N23761, N23760, N23759, N23758, N23757, N23756, N23755, N23754, N23753, N23752, N23751, N23750, N23749, N23748, N23747, N23746, N23745, N23744, N23743, N23742, N23741, N23740, N23739, N23738, N23737, N23736, N23735, N23734, N23733, N23732, N23731, N23730, N23729, N23728, N23727, N23726, N23725, N23724, N23723, N23722, N23721, N23720, N23719, N23718, N23717, N23716, N23715, N23714, N23713, N23712, N23711, N23710, N23709, N23708, N23707, N23706, N23705, N23704, N23703, N23702, N23701, N23700, N23699, N23698, N23697, N23696, N23695, N23694, N23693, N23692, N23691, N23690, N23689, N23688, N23687, N23686, N23685, N23684, N23683, N23682, N23681, N23680, N23679, N23678, N23677, N23676, N23675, N23674, N23673, N23672, N23671, N23670, N23669, N23668, N23667, N23666, N23665, N23664, N23663, N23662, N23661, N23660, N23659, N23658, N23657, N23656, N23655, N23654, N23653, N23652, N23651, N23650, N23649, N23648, N23647, N23646, N23645, N23644, N23643, N23642, N23641, N23640, N23639, N23638, N23637, N23636, N23635, N23634, N23633, N23632, N23631, N23630, N23629, N23628, N23627, N23626, N23625, N23624, N23623, N23622, N23621, N23620, N23619, N23618, N23617, N23616, N23615, N23614, N23613, N23612, N23611, N23610, N23609, N23608, N23607, N23606, N23605, N23604, N23603, N23602, N23601, N23600, N23599, N23598, N23597, N23596, N23595, N23594, N23593, N23592, N23591, N23590, N23589, N23588, N23587, N23586, N23585, N23584, N23583, N23582, N23581, N23580, N23579, N23578, N23577, N23576, N23575, N23574, N23573, N23572, N23571, N23570, N23569, N23568, N23567, N23566, N23565, N23564, N23563, N23562, N23561, N23560, N23559, N23558, N23557, N23556, N23555, N23554, N23553, N23552, N23551, N23550, N23549, N23548, N23547, N23546, N23545, N23544, N23543, N23542, N23541, N23540, N23539, N23538, N23537, N23536, N23535, N23534, N23533, N23532, N23531, N23530, N23529, N23528, N23527, N23526, N23525, N23524, N23523, N23522, N23521, N23520, N23519, N23518, N23517, N23516, N23515, N23514, N23513, N23512, N23511, N23510, N23509, N23508, N23507, N23506, N23505, N23504, N23503, N23502, N23501, N23500, N23499, N23498, N23497, N23496, N23495, N23494, N23493, N23492, N23491, N23490, N23489, N23488, N23487, N23486, N23485, N23484, N23483, N23482, N23481, N23480, N23479, N23478, N23477, N23476, N23475, N23474, N23473, N23472, N23471, N23470, N23469, N23468, N23467, N23466, N23465, N23464, N23463, N23462, N23461, N23460, N23459, N23458, N23457, N23456, N23455, N23454, N23453, N23452, N23451, N23450, N23449, N23448, N23447, N23446, N23445, N23444, N23443, N23442, N23441, N23440, N23439, N23438, N23437, N23436, N23435, N23434, N23433, N23432, N23431, N23430, N23429, N23428, N23427, N23426, N23425, N23424, N23423, N23422, N23421, N23420, N23419, N23418, N23417, N23416, N23415, N23414, N23413, N23412, N23411, N23410, N23409, N23408, N23407, N23406, N23405, N23404, N23403, N23402, N23401, N23400, N23399, N23398, N23397, N23396, N23395, N23394, N23393, N23392, N23391, N23390, N23389, N23388, N23387, N23386, N23385, N23384, N23383, N23382, N23381, N23380, N23379, N23378, N23377, N23376, N23375, N23374, N23373, N23372, N23371, N23370, N23369, N23368, N23367, N23366, N23365, N23364, N23363, N23362, N23361, N23360, N23359, N23358, N23357, N23356, N23355, N23354, N23353, N23352, N23351, N23350, N23349, N23348, N23347, N23346, N23345, N23344, N23343, N23342, N23341, N23340, N23339, N23338, N23337, N23336, N23335, N23334, N23333, N23332, N23331, N23330, N23329, N23328, N23327, N23326, N23325, N23324, N23323, N23322, N23321, N23320, N23319, N23318, N23317, N23316, N23315, N23314, N23313, N23312, N23311, N23310, N23309, N23308, N23307, N23306, N23305, N23304, N23303, N23302, N23301, N23300, N23299, N23298, N23297, N23296, N23295, N23294, N23293, N23292, N23291, N23290, N23289, N23288, N23287, N23286, N23285, N23284, N23283, N23282, N23281, N23280, N23279, N23278, N23277, N23276, N23275, N23274, N23273, N23272, N23271, N23270, N23269, N23268, N23267, N23266, N23265, N23264, N23263, N23262, N23261, N23260, N23259, N23258, N23257, N23256, N23255, N23254, N23253, N23252, N23251, N23250, N23249, N23248, N23247, N23246, N23245, N23244, N23243, N23242, N23241, N23240, N23239, N23238, N23237, N23236, N23235, N23234, N23233, N23232, N23231, N23230, N23229, N23228, N23227, N23226, N23225, N23224, N23223, N23222, N23221, N23220, N23219, N23218, N23217, N23216, N23215, N23214, N23213, N23212, N23211, N23210, N23209, N23208, N23207, N23206, N23205, N23204, N23203, N23202, N23201, N23200, N23199, N23198, N23197, N23196, N23195, N23194, N23193, N23192, N23191, N23190, N23189, N23188, N23187, N23186, N23185, N23184, N23183, N23182, N23181, N23180, N23179, N23178, N23177, N23176, N23175, N23174, N23173, N23172, N23171, N23170, N23169, N23168, N23167, N23166, N23165, N23164, N23163, N23162, N23161, N23160, N23159, N23158, N23157, N23156, N23155, N23154, N23153, N23152, N23151, N23150, N23149, N23148, N23147, N23146, N23145, N23144, N23143, N23142, N23141, N23140, N23139, N23138, N23137, N23136, N23135, N23134, N23133, N23132, N23131, N23130, N23129, N23128, N23127, N23126, N23125, N23124, N23123, N23122, N23121, N23120, N23119, N23118, N23117, N23116, N23115, N23114, N23113, N23112, N23111, N23110, N23109, N23108, N23107, N23106, N23105, N23104, N23103, N23102, N23101, N23100, N23099, N23098, N23097, N23096, N23095, N23094, N23093, N23092, N23091, N23090, N23089, N23088, N23087, N23086, N23085, N23084, N23083, N23082, N23081, N23080, N23079, N23078, N23077, N23076, N23075, N23074, N23073, N23072, N23071, N23070, N23069, N23068, N23067, N23066, N23065, N23064, N23063, N23062, N23061, N23060, N23059, N23058, N23057, N23056, N23055, N23054, N23053, N23052, N23051, N23050, N23049, N23048, N23047, N23046, N23045, N23044, N23043, N23042, N23041, N23040, N23039, N23038, N23037, N23036, N23035, N23034, N23033, N23032, N23031, N23030, N23029, N23028, N23027, N23026, N23025, N23024, N23023, N23022, N23021, N23020, N23019, N23018, N23017, N23016, N23015, N23014, N23013, N23012, N23011, N23010, N23009, N23008, N23007, N23006, N23005, N23004, N23003, N23002, N23001, N23000, N22999, N22998, N22997, N22996, N22995, N22994, N22993, N22992, N22991, N22990, N22989, N22988, N22987, N22986, N22985, N22984, N22983, N22982, N22981, N22980, N22979, N22978, N22977, N22976, N22975, N22974, N22973, N22972, N22971, N22970, N22969, N22968, N22967, N22966, N22965, N22964, N22963, N22962, N22961, N22960, N22959, N22958, N22957, N22956, N22955, N22954, N22953, N22952, N22951, N22950, N22949, N22948, N22947, N22946, N22945, N22944, N22943, N22942, N22941, N22940, N22939, N22938, N22937, N22936, N22935, N22934, N22933, N22932, N22931, N22930, N22929, N22928, N22927, N22926, N22925, N22924, N22923, N22922, N22921, N22920, N22919, N22918, N22917, N22916, N22915, N22914, N22913, N22912, N22911, N22910, N22909, N22908, N22907, N22906, N22905, N22904, N22903, N22902, N22901, N22900, N22899, N22898, N22897, N22896, N22895, N22894, N22893, N22892, N22891, N22890, N22889, N22888, N22887, N22886, N22885, N22884, N22883, N22882, N22881, N22880, N22879, N22878, N22877, N22876, N22875, N22874, N22873, N22872, N22871, N22870, N22869, N22868, N22867, N22866, N22865, N22864, N22863, N22862, N22861, N22860, N22859, N22858, N22857, N22856, N22855, N22854, N22853, N22852, N22851, N22850, N22849, N22848, N22847, N22846, N22845, N22844, N22843, N22842, N22841, N22840, N22839, N22838, N22837, N22836, N22835, N22834, N22833, N22832, N22831, N22830, N22829, N22828, N22827, N22826, N22825, N22824, N22823, N22822, N22821, N22820, N22819, N22818, N22817, N22816, N22815, N22814, N22813, N22812, N22811, N22810, N22809, N22808, N22807, N22806, N22805, N22804, N22803, N22802, N22801, N22800, N22799, N22798, N22797, N22796, N22795, N22794, N22793, N22792, N22791, N22790, N22789, N22788, N22787, N22786, N22785, N22784, N22783, N22782, N22781, N22780, N22779, N22778, N22777, N22776, N22775, N22774, N22773, N22772, N22771, N22770, N22769, N22768, N22767, N22766, N22765, N22764, N22763, N22762, N22761, N22760, N22759, N22758, N22757, N22756, N22755, N22754, N22753, N22752, N22751, N22750, N22749, N22748, N22747, N22746, N22745, N22744, N22743, N22742, N22741, N22740, N22739, N22738, N22737, N22736, N22735, N22734, N22733, N22732, N22731, N22730, N22729, N22728, N22727, N22726, N22725, N22724, N22723, N22722, N22721, N22720, N22719, N22718, N22717, N22716, N22715, N22714, N22713, N22712, N22711, N22710, N22709, N22708, N22707, N22706, N22705, N22704, N22703, N22702, N22701, N22700, N22699, N22698, N22697, N22696, N22695, N22694, N22693, N22692, N22691, N22690, N22689, N22688, N22687, N22686, N22685, N22684, N22683, N22682, N22681, N22680, N22679, N22678, N22677, N22676, N22675, N22674, N22673, N22672, N22671, N22670, N22669, N22668, N22667, N22666, N22665, N22664, N22663, N22662, N22661, N22660, N22659, N22658, N22657, N22656, N22655, N22654, N22653, N22652, N22651, N22650, N22649, N22648, N22647, N22646, N22645, N22644, N22643, N22642, N22641, N22640, N22639, N22638, N22637, N22636, N22635, N22634, N22633, N22632, N22631, N22630, N22629, N22628, N22627, N22626, N22625, N22624, N22623, N22622, N22621, N22620, N22619, N22618, N22617, N22616, N22615, N22614, N22613, N22612, N22611, N22610, N22609, N22608, N22607, N22606, N22605, N22604, N22603, N22602, N22601, N22600, N22599, N22598, N22597, N22596, N22595, N22594, N22593, N22592, N22591, N22590, N22589, N22588, N22587, N22586, N22585, N22584, N22583, N22582, N22581, N22580, N22579, N22578, N22577, N22576, N22575, N22574, N22573, N22572, N22571, N22570, N22569, N22568, N22567, N22566, N22565, N22564, N22563, N22562, N22561, N22560, N22559, N22558, N22557, N22556, N22555, N22554, N22553, N22552, N22551, N22550, N22549, N22548, N22547, N22546, N22545, N22544, N22543, N22542, N22541, N22540, N22539, N22538, N22537, N22536, N22535, N22534, N22533, N22532, N22531, N22530, N22529, N22528, N22527 } = (N192)? { N18909, N18908, N18907, N18906, N18905, N18904, N18903, N18902, N18901, N18900, N18899, N18898, N18897, N18896, N18895, N18894, N18893, N18892, N18891, N18890, N18889, N18888, N18887, N18886, N18885, N18884, N18883, N18882, N18881, N18880, N18879, N18878, N18877, N18876, N18875, N18874, N18873, N18872, N18871, N18870, N18869, N18868, N18867, N18866, N18865, N18864, N18863, N18862, N18861, N18860, N18859, N18858, N18857, N18856, N18855, N18854, N18853, N18852, N18851, N18850, N18849, N18848, N18847, N18846, N18381, N22526, N22525, N22524, N22523, N22522, N22521, N22520, N22519, N22518, N22517, N22516, N22515, N22514, N22513, N22512, N22511, N22510, N22509, N22508, N22507, N22506, N22505, N22504, N22503, N22502, N22501, N22500, N22499, N22498, N22497, N22496, N22495, N22494, N22493, N22492, N22491, N22490, N22489, N22488, N22487, N22486, N22485, N22484, N22483, N22482, N22481, N22480, N22479, N22478, N22477, N22476, N22475, N22474, N22473, N22472, N22471, N22470, N22469, N22468, N22467, N22466, N22465, N22464, N22463, N22462, N22461, N22460, N22459, N22458, N22457, N22456, N22455, N22454, N22453, N22452, N22451, N22450, N22449, N22448, N22447, N22446, N22445, N22444, N22443, N22442, N22441, N22440, N22439, N22438, N22437, N22436, N22435, N22434, N22433, N22432, N22431, N22430, N22429, N22428, N22427, N22426, N22425, N22424, N22423, N22422, N22421, N22420, N22419, N22418, N22417, N22416, N22415, N22414, N22413, N22412, N22411, N22410, N22409, N22408, N22407, N22406, N22405, N22404, N22403, N22402, N22401, N22400, N22399, N22398, N19421, N19420, N19419, N19418, N19417, N19416, N19415, N19414, N19413, N19412, N19411, N19410, N19409, N19408, N19407, N19406, N19405, N19404, N19403, N19402, N19401, N19400, N19399, N19398, N19397, N19396, N19395, N19394, N19393, N19392, N19391, N19390, N19389, N19388, N19387, N19386, N19385, N19384, N19383, N19382, N19381, N19380, N19379, N19378, N19377, N19376, N19375, N19374, N19373, N19372, N19371, N19370, N19369, N19368, N19367, N19366, N19365, N19364, N19363, N19362, N19361, N19360, N19359, N19358, N18844, N18843, N18842, N18841, N18840, N18839, N18838, N18837, N18836, N18835, N18834, N18833, N18832, N18831, N18830, N18829, N18828, N18827, N18826, N18825, N18824, N18823, N18822, N18821, N18820, N18819, N18818, N18817, N18816, N18815, N18814, N18813, N18812, N18811, N18810, N18809, N18808, N18807, N18806, N18805, N18804, N18803, N18802, N18801, N18800, N18799, N18798, N18797, N18796, N18795, N18794, N18793, N18792, N18791, N18790, N18789, N18788, N18787, N18786, N18785, N18784, N18783, N18782, N18781, N18380, N22397, N22396, N22395, N22394, N22393, N22392, N22391, N22390, N22389, N22388, N22387, N22386, N22385, N22384, N22383, N22382, N22381, N22380, N22379, N22378, N22377, N22376, N22375, N22374, N22373, N22372, N22371, N22370, N22369, N22368, N22367, N22366, N22365, N22364, N22363, N22362, N22361, N22360, N22359, N22358, N22357, N22356, N22355, N22354, N22353, N22352, N22351, N22350, N22349, N22348, N22347, N22346, N22345, N22344, N22343, N22342, N22341, N22340, N22339, N22338, N22337, N22336, N22335, N22334, N22333, N22332, N22331, N22330, N22329, N22328, N22327, N22326, N22325, N22324, N22323, N22322, N22321, N22320, N22319, N22318, N22317, N22316, N22315, N22314, N22313, N22312, N22311, N22310, N22309, N22308, N22307, N22306, N22305, N22304, N22303, N22302, N22301, N22300, N22299, N22298, N22297, N22296, N22295, N22294, N22293, N22292, N22291, N22290, N22289, N22288, N22287, N22286, N22285, N22284, N22283, N22282, N22281, N22280, N22279, N22278, N22277, N22276, N22275, N22274, N22273, N22272, N22271, N22270, N22269, N19357, N19356, N19355, N19354, N19353, N19352, N19351, N19350, N19349, N19348, N19347, N19346, N19345, N19344, N19343, N19342, N19341, N19340, N19339, N19338, N19337, N19336, N19335, N19334, N19333, N19332, N19331, N19330, N19329, N19328, N19327, N19326, N19325, N19324, N19323, N19322, N19321, N19320, N19319, N19318, N19317, N19316, N19315, N19314, N19313, N19312, N19311, N19310, N19309, N19308, N19307, N19306, N19305, N19304, N19303, N19302, N19301, N19300, N19299, N19298, N19297, N19296, N19295, N19294, N18779, N18778, N18777, N18776, N18775, N18774, N18773, N18772, N18771, N18770, N18769, N18768, N18767, N18766, N18765, N18764, N18763, N18762, N18761, N18760, N18759, N18758, N18757, N18756, N18755, N18754, N18753, N18752, N18751, N18750, N18749, N18748, N18747, N18746, N18745, N18744, N18743, N18742, N18741, N18740, N18739, N18738, N18737, N18736, N18735, N18734, N18733, N18732, N18731, N18730, N18729, N18728, N18727, N18726, N18725, N18724, N18723, N18722, N18721, N18720, N18719, N18718, N18717, N18716, N18379, N22268, N22267, N22266, N22265, N22264, N22263, N22262, N22261, N22260, N22259, N22258, N22257, N22256, N22255, N22254, N22253, N22252, N22251, N22250, N22249, N22248, N22247, N22246, N22245, N22244, N22243, N22242, N22241, N22240, N22239, N22238, N22237, N22236, N22235, N22234, N22233, N22232, N22231, N22230, N22229, N22228, N22227, N22226, N22225, N22224, N22223, N22222, N22221, N22220, N22219, N22218, N22217, N22216, N22215, N22214, N22213, N22212, N22211, N22210, N22209, N22208, N22207, N22206, N22205, N22204, N22203, N22202, N22201, N22200, N22199, N22198, N22197, N22196, N22195, N22194, N22193, N22192, N22191, N22190, N22189, N22188, N22187, N22186, N22185, N22184, N22183, N22182, N22181, N22180, N22179, N22178, N22177, N22176, N22175, N22174, N22173, N22172, N22171, N22170, N22169, N22168, N22167, N22166, N22165, N22164, N22163, N22162, N22161, N22160, N22159, N22158, N22157, N22156, N22155, N22154, N22153, N22152, N22151, N22150, N22149, N22148, N22147, N22146, N22145, N22144, N22143, N22142, N22141, N22140, N19293, N19292, N19291, N19290, N19289, N19288, N19287, N19286, N19285, N19284, N19283, N19282, N19281, N19280, N19279, N19278, N19277, N19276, N19275, N19274, N19273, N19272, N19271, N19270, N19269, N19268, N19267, N19266, N19265, N19264, N19263, N19262, N19261, N19260, N19259, N19258, N19257, N19256, N19255, N19254, N19253, N19252, N19251, N19250, N19249, N19248, N19247, N19246, N19245, N19244, N19243, N19242, N19241, N19240, N19239, N19238, N19237, N19236, N19235, N19234, N19233, N19232, N19231, N19230, N18714, N18713, N18712, N18711, N18710, N18709, N18708, N18707, N18706, N18705, N18704, N18703, N18702, N18701, N18700, N18699, N18698, N18697, N18696, N18695, N18694, N18693, N18692, N18691, N18690, N18689, N18688, N18687, N18686, N18685, N18684, N18683, N18682, N18681, N18680, N18679, N18678, N18677, N18676, N18675, N18674, N18673, N18672, N18671, N18670, N18669, N18668, N18667, N18666, N18665, N18664, N18663, N18662, N18661, N18660, N18659, N18658, N18657, N18656, N18655, N18654, N18653, N18652, N18651, N18378, N22139, N22138, N22137, N22136, N22135, N22134, N22133, N22132, N22131, N22130, N22129, N22128, N22127, N22126, N22125, N22124, N22123, N22122, N22121, N22120, N22119, N22118, N22117, N22116, N22115, N22114, N22113, N22112, N22111, N22110, N22109, N22108, N22107, N22106, N22105, N22104, N22103, N22102, N22101, N22100, N22099, N22098, N22097, N22096, N22095, N22094, N22093, N22092, N22091, N22090, N22089, N22088, N22087, N22086, N22085, N22084, N22083, N22082, N22081, N22080, N22079, N22078, N22077, N22076, N22075, N22074, N22073, N22072, N22071, N22070, N22069, N22068, N22067, N22066, N22065, N22064, N22063, N22062, N22061, N22060, N22059, N22058, N22057, N22056, N22055, N22054, N22053, N22052, N22051, N22050, N22049, N22048, N22047, N22046, N22045, N22044, N22043, N22042, N22041, N22040, N22039, N22038, N22037, N22036, N22035, N22034, N22033, N22032, N22031, N22030, N22029, N22028, N22027, N22026, N22025, N22024, N22023, N22022, N22021, N22020, N22019, N22018, N22017, N22016, N22015, N22014, N22013, N22012, N22011, N19229, N19228, N19227, N19226, N19225, N19224, N19223, N19222, N19221, N19220, N19219, N19218, N19217, N19216, N19215, N19214, N19213, N19212, N19211, N19210, N19209, N19208, N19207, N19206, N19205, N19204, N19203, N19202, N19201, N19200, N19199, N19198, N19197, N19196, N19195, N19194, N19193, N19192, N19191, N19190, N19189, N19188, N19187, N19186, N19185, N19184, N19183, N19182, N19181, N19180, N19179, N19178, N19177, N19176, N19175, N19174, N19173, N19172, N19171, N19170, N19169, N19168, N19167, N19166, N18649, N18648, N18647, N18646, N18645, N18644, N18643, N18642, N18641, N18640, N18639, N18638, N18637, N18636, N18635, N18634, N18633, N18632, N18631, N18630, N18629, N18628, N18627, N18626, N18625, N18624, N18623, N18622, N18621, N18620, N18619, N18618, N18617, N18616, N18615, N18614, N18613, N18612, N18611, N18610, N18609, N18608, N18607, N18606, N18605, N18604, N18603, N18602, N18601, N18600, N18599, N18598, N18597, N18596, N18595, N18594, N18593, N18592, N18591, N18590, N18589, N18588, N18587, N18586, N18377, N22010, N22009, N22008, N22007, N22006, N22005, N22004, N22003, N22002, N22001, N22000, N21999, N21998, N21997, N21996, N21995, N21994, N21993, N21992, N21991, N21990, N21989, N21988, N21987, N21986, N21985, N21984, N21983, N21982, N21981, N21980, N21979, N21978, N21977, N21976, N21975, N21974, N21973, N21972, N21971, N21970, N21969, N21968, N21967, N21966, N21965, N21964, N21963, N21962, N21961, N21960, N21959, N21958, N21957, N21956, N21955, N21954, N21953, N21952, N21951, N21950, N21949, N21948, N21947, N21946, N21945, N21944, N21943, N21942, N21941, N21940, N21939, N21938, N21937, N21936, N21935, N21934, N21933, N21932, N21931, N21930, N21929, N21928, N21927, N21926, N21925, N21924, N21923, N21922, N21921, N21920, N21919, N21918, N21917, N21916, N21915, N21914, N21913, N21912, N21911, N21910, N21909, N21908, N21907, N21906, N21905, N21904, N21903, N21902, N21901, N21900, N21899, N21898, N21897, N21896, N21895, N21894, N21893, N21892, N21891, N21890, N21889, N21888, N21887, N21886, N21885, N21884, N21883, N21882, N19165, N19164, N19163, N19162, N19161, N19160, N19159, N19158, N19157, N19156, N19155, N19154, N19153, N19152, N19151, N19150, N19149, N19148, N19147, N19146, N19145, N19144, N19143, N19142, N19141, N19140, N19139, N19138, N19137, N19136, N19135, N19134, N19133, N19132, N19131, N19130, N19129, N19128, N19127, N19126, N19125, N19124, N19123, N19122, N19121, N19120, N19119, N19118, N19117, N19116, N19115, N19114, N19113, N19112, N19111, N19110, N19109, N19108, N19107, N19106, N19105, N19104, N19103, N19102, N18584, N18583, N18582, N18581, N18580, N18579, N18578, N18577, N18576, N18575, N18574, N18573, N18572, N18571, N18570, N18569, N18568, N18567, N18566, N18565, N18564, N18563, N18562, N18561, N18560, N18559, N18558, N18557, N18556, N18555, N18554, N18553, N18552, N18551, N18550, N18549, N18548, N18547, N18546, N18545, N18544, N18543, N18542, N18541, N18540, N18539, N18538, N18537, N18536, N18535, N18534, N18533, N18532, N18531, N18530, N18529, N18528, N18527, N18526, N18525, N18524, N18523, N18522, N18521, N18376, N21881, N21880, N21879, N21878, N21877, N21876, N21875, N21874, N21873, N21872, N21871, N21870, N21869, N21868, N21867, N21866, N21865, N21864, N21863, N21862, N21861, N21860, N21859, N21858, N21857, N21856, N21855, N21854, N21853, N21852, N21851, N21850, N21849, N21848, N21847, N21846, N21845, N21844, N21843, N21842, N21841, N21840, N21839, N21838, N21837, N21836, N21835, N21834, N21833, N21832, N21831, N21830, N21829, N21828, N21827, N21826, N21825, N21824, N21823, N21822, N21821, N21820, N21819, N21818, N21817, N21816, N21815, N21814, N21813, N21812, N21811, N21810, N21809, N21808, N21807, N21806, N21805, N21804, N21803, N21802, N21801, N21800, N21799, N21798, N21797, N21796, N21795, N21794, N21793, N21792, N21791, N21790, N21789, N21788, N21787, N21786, N21785, N21784, N21783, N21782, N21781, N21780, N21779, N21778, N21777, N21776, N21775, N21774, N21773, N21772, N21771, N21770, N21769, N21768, N21767, N21766, N21765, N21764, N21763, N21762, N21761, N21760, N21759, N21758, N21757, N21756, N21755, N21754, N21753, N19101, N19100, N19099, N19098, N19097, N19096, N19095, N19094, N19093, N19092, N19091, N19090, N19089, N19088, N19087, N19086, N19085, N19084, N19083, N19082, N19081, N19080, N19079, N19078, N19077, N19076, N19075, N19074, N19073, N19072, N19071, N19070, N19069, N19068, N19067, N19066, N19065, N19064, N19063, N19062, N19061, N19060, N19059, N19058, N19057, N19056, N19055, N19054, N19053, N19052, N19051, N19050, N19049, N19048, N19047, N19046, N19045, N19044, N19043, N19042, N19041, N19040, N19039, N19038, N18519, N18518, N18517, N18516, N18515, N18514, N18513, N18512, N18511, N18510, N18509, N18508, N18507, N18506, N18505, N18504, N18503, N18502, N18501, N18500, N18499, N18498, N18497, N18496, N18495, N18494, N18493, N18492, N18491, N18490, N18489, N18488, N18487, N18486, N18485, N18484, N18483, N18482, N18481, N18480, N18479, N18478, N18477, N18476, N18475, N18474, N18473, N18472, N18471, N18470, N18469, N18468, N18467, N18466, N18465, N18464, N18463, N18462, N18461, N18460, N18459, N18458, N18457, N18456, N18375, N21752, N21751, N21750, N21749, N21748, N21747, N21746, N21745, N21744, N21743, N21742, N21741, N21740, N21739, N21738, N21737, N21736, N21735, N21734, N21733, N21732, N21731, N21730, N21729, N21728, N21727, N21726, N21725, N21724, N21723, N21722, N21721, N21720, N21719, N21718, N21717, N21716, N21715, N21714, N21713, N21712, N21711, N21710, N21709, N21708, N21707, N21706, N21705, N21704, N21703, N21702, N21701, N21700, N21699, N21698, N21697, N21696, N21695, N21694, N21693, N21692, N21691, N21690, N21689, N21688, N21687, N21686, N21685, N21684, N21683, N21682, N21681, N21680, N21679, N21678, N21677, N21676, N21675, N21674, N21673, N21672, N21671, N21670, N21669, N21668, N21667, N21666, N21665, N21664, N21663, N21662, N21661, N21660, N21659, N21658, N21657, N21656, N21655, N21654, N21653, N21652, N21651, N21650, N21649, N21648, N21647, N21646, N21645, N21644, N21643, N21642, N21641, N21640, N21639, N21638, N21637, N21636, N21635, N21634, N21633, N21632, N21631, N21630, N21629, N21628, N21627, N21626, N21625, N21624, N19037, N19036, N19035, N19034, N19033, N19032, N19031, N19030, N19029, N19028, N19027, N19026, N19025, N19024, N19023, N19022, N19021, N19020, N19019, N19018, N19017, N19016, N19015, N19014, N19013, N19012, N19011, N19010, N19009, N19008, N19007, N19006, N19005, N19004, N19003, N19002, N19001, N19000, N18999, N18998, N18997, N18996, N18995, N18994, N18993, N18992, N18991, N18990, N18989, N18988, N18987, N18986, N18985, N18984, N18983, N18982, N18981, N18980, N18979, N18978, N18977, N18976, N18975, N18974, N18454, N18453, N18452, N18451, N18450, N18449, N18448, N18447, N18446, N18445, N18444, N18443, N18442, N18441, N18440, N18439, N18438, N18437, N18436, N18435, N18434, N18433, N18432, N18431, N18430, N18429, N18428, N18427, N18426, N18425, N18424, N18423, N18422, N18421, N18420, N18419, N18418, N18417, N18416, N18415, N18414, N18413, N18412, N18411, N18410, N18409, N18408, N18407, N18406, N18405, N18404, N18403, N18402, N18401, N18400, N18399, N18398, N18397, N18396, N18395, N18394, N18393, N18392, N18391, N18374, N21623, N21622, N21621, N21620, N21619, N21618, N21617, N21616, N21615, N21614, N21613, N21612, N21611, N21610, N21609, N21608, N21607, N21606, N21605, N21604, N21603, N21602, N21601, N21600, N21599, N21598, N21597, N21596, N21595, N21594, N21593, N21592, N21591, N21590, N21589, N21588, N21587, N21586, N21585, N21584, N21583, N21582, N21581, N21580, N21579, N21578, N21577, N21576, N21575, N21574, N21573, N21572, N21571, N21570, N21569, N21568, N21567, N21566, N21565, N21564, N21563, N21562, N21561, N21560, N21559, N21558, N21557, N21556, N21555, N21554, N21553, N21552, N21551, N21550, N21549, N21548, N21547, N21546, N21545, N21544, N21543, N21542, N21541, N21540, N21539, N21538, N21537, N21536, N21535, N21534, N21533, N21532, N21531, N21530, N21529, N21528, N21527, N21526, N21525, N21524, N21523, N21522, N21521, N21520, N21519, N21518, N21517, N21516, N21515, N21514, N21513, N21512, N21511, N21510, N21509, N21508, N21507, N21506, N21505, N21504, N21503, N21502, N21501, N21500, N21499, N21498, N21497, N21496, N21495, N18973, N18972, N18971, N18970, N18969, N18968, N18967, N18966, N18965, N18964, N18963, N18962, N18961, N18960, N18959, N18958, N18957, N18956, N18955, N18954, N18953, N18952, N18951, N18950, N18949, N18948, N18947, N18946, N18945, N18944, N18943, N18942, N18941, N18940, N18939, N18938, N18937, N18936, N18935, N18934, N18933, N18932, N18931, N18930, N18929, N18928, N18927, N18926, N18925, N18924, N18923, N18922, N18921, N18920, N18919, N18918, N18917, N18916, N18915, N18914, N18913, N18912, N18911, N18910 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18373)? { N18355, N18354, N18353, N18352, N18351, N18350, N18349, N18348, N18347, N18346, N18345, N18344, N18343, N18342, N18341, N18340, N18339, N18338, N18337, N18336, N18335, N18334, N18333, N18332, N18331, N18330, N18329, N18328, N18327, N18326, N18325, N18324, N18323, N18322, N18321, N18320, N18319, N18318, N18317, N18316, N18315, N18314, N18313, N18312, N18311, N18310, N18309, N18308, N18307, N18306, N18305, N18304, N18303, N18302, N18301, N18300, N18299, N18298, N18297, N18296, N18295, N18294, N18293, N18292, N18291, N18290, N18289, N18288, N18287, N18286, N18285, N18284, N18283, N18282, N18281, N18280, N18279, N18278, N18277, N18276, N18275, N18274, N18273, N18272, N18271, N18270, N18269, N18268, N18267, N18266, N18265, N18264, N18263, N18262, N18261, N18260, N18259, N18258, N18257, N18256, N18255, N18254, N18253, N18252, N18251, N18250, N18249, N18248, N18247, N18246, N18245, N18244, N18243, N18242, N18241, N18240, N18239, N18238, N18237, N18236, N18235, N18234, N18233, N18232, N18231, N18230, N18229, N18228, N18227, N18226, N18225, N18224, N18223, N18222, N18221, N18220, N18219, N18218, N18217, N18216, N18215, N18214, N18213, N18212, N18211, N18210, N18209, N18208, N18207, N18206, N18205, N18204, N18203, N18202, N18201, N18200, N18199, N18198, N18197, N18196, N18195, N18194, N18193, N18192, N18191, N18190, N18189, N18188, N18187, N18186, N18185, N18184, N18183, N18182, N18181, N18180, N18179, N18178, N18177, N18176, N18175, N18174, N18173, N18172, N18171, N18170, N18169, N18168, N18167, N18166, N18165, N18164, N18163, N18162, N18161, N18160, N18159, N18158, N18157, N18156, N18155, N18154, N18153, N18152, N18151, N18150, N18149, N18148, N18147, N18146, N18145, N18144, N18143, N18142, N18141, N18140, N18139, N18138, N18137, N18136, N18135, N18134, N18133, N18132, N18131, N18130, N18129, N18128, N18127, N18126, N18125, N18124, N18123, N18122, N18121, N18120, N18119, N18118, N18117, N18116, N18115, N18114, N18113, N18112, N18111, N18110, N18109, N18108, N18107, N18106, N18105, N18104, N18103, N18102, N18101, N18100, N18099, N18098, N18097, N18096, N18095, N18094, N18093, N18092, N18091, N18090, N18089, N18088, N18087, N18086, N18085, N18084, N18083, N18082, N18081, N18080, N18079, N18078, N18077, N18076, N18075, N18074, N18073, N18072, N18071, N18070, N18069, N18068, N18067, N18066, N18065, N18064, N18063, N18062, N18061, N18060, N18059, N18058, N18057, N18056, N18055, N18054, N18053, N18052, N18051, N18050, N18049, N18048, N18047, N18046, N18045, N18044, N18043, N18042, N18041, N18040, N18039, N18038, N18037, N18036, N18035, N18034, N18033, N18032, N18031, N18030, N18029, N18028, N18027, N18026, N18025, N18024, N18023, N18022, N18021, N18020, N18019, N18018, N18017, N18016, N18015, N18014, N18013, N18012, N18011, N18010, N18009, N18008, N18007, N18006, N18005, N18004, N18003, N18002, N18001, N18000, N17999, N17998, N17997, N17996, N17995, N17994, N17993, N17992, N17991, N17990, N17989, N17988, N17987, N17986, N17985, N17984, N17983, N17982, N17981, N17980, N17979, N17978, N17977, N17976, N17975, N17974, N17973, N17972, N17971, N17970, N17969, N17968, N17967, N17966, N17965, N17964, N17963, N17962, N17961, N17960, N17959, N17958, N17957, N17956, N17955, N17954, N17953, N17952, N17951, N17950, N17949, N17948, N17947, N17946, N17945, N17944, N17943, N17942, N17941, N17940, N17939, N17938, N17937, N17936, N17935, N17934, N17933, N17932, N17931, N17930, N17929, N17928, N17927, N17926, N17925, N17924, N17923, N17922, N17921, N17920, N17919, N17918, N17917, N17916, N17915, N17914, N17913, N17912, N17911, N17910, N17909, N17908, N17907, N17906, N17905, N17904, N17903, N17902, N17901, N17900, N17899, N17898, N17897, N17896, N17895, N17894, N17893, N17892, N17891, N17890, N17889, N17888, N17887, N17886, N17885, N17884, N17883, N17882, N17881, N17880, N17879, N17878, N17877, N17876, N17875, N17874, N17873, N17872, N17871, N17870, N17869, N17868, N17867, N17866, N17865, N17864, N17863, N17862, N17861, N17860, N17859, N17858, N17857, N17856, N17855, N17854, N17853, N17852, N17851, N17850, N17849, N17848, N17847, N17846, N17845, N17844, N17843, N17842, N17841, N17840, N17839, N17838, N17837, N17836, N17835, N17834, N17833, N17832, N17831, N17830, N17829, N17828, N17827, N17826, N17825, N17824, N17823, N17822, N17821, N17820, N17819, N17818, N17817, N17816, N17815, N17814, N17813, N17812, N17811, N17810, N17809, N17808, N17807, N17806, N17805, N17804, N17803, N17802, N17801, N17800, N17799, N17798, N17797, N17796, N17795, N17794, N17793, N17792, N17791, N17790, N17789, N17788, N17787, N17786, N17785, N17784, N17783, N17782, N17781, N17780, N17779, N17778, N17777, N17776, N17775, N17774, N17773, N17772, N17771, N17770, N17769, N17768, N17767, N17766, N17765, N17764, N17763, N17762, N17761, N17760, N17759, N17758, N17757, N17756, N17755, N17754, N17753, N17752, N17751, N17750, N17749, N17748, N17747, N17746, N17745, N17744, N17743, N17742, N17741, N17740, N17739, N17738, N17737, N17736, N17735, N17734, N17733, N17732, N17731, N17730, N17729, N17728, N17727, N17726, N17725, N17724, N17723, N17722, N17721, N17720, N17719, N17718, N17717, N17716, N17715, N17714, N17713, N17712, N17711, N17710, N17709, N17708, N17707, N17706, N17705, N17704, N17703, N17702, N17701, N17700, N17699, N17698, N17697, N17696, N17695, N17694, N17693, N17692, N17691, N17690, N17689, N17688, N17687, N17686, N17685, N17684, N17683, N17682, N17681, N17680, N17679, N17678, N17677, N17676, N17675, N17674, N17673, N17672, N17671, N17670, N17669, N17668, N17667, N17666, N17665, N17664, N17663, N17662, N17661, N17660, N17659, N17658, N17657, N17656, N17655, N17654, N17653, N17652, N17651, N17650, N17649, N17648, N17647, N17646, N17645, N17644, N17643, N17642, N17641, N17640, N17639, N17638, N17637, N17636, N17635, N17634, N17633, N17632, N17631, N17630, N17629, N17628, N17627, N17626, N17625, N17624, N17623, N17622, N17621, N17620, N17619, N17618, N17617, N17616, N17615, N17614, N17613, N17612, N17611, N17610, N17609, N17608, N17607, N17606, N17605, N17604, N17603, N17602, N17601, N17600, N17599, N17598, N17597, N17596, N17595, N17594, N17593, N17592, N17591, N17590, N17589, N17588, N17587, N17586, N17585, N17584, N17583, N17582, N17581, N17580, N17579, N17578, N17577, N17576, N17575, N17574, N17573, N17572, N17571, N17570, N17569, N17568, N17567, N17566, N17565, N17564, N17563, N17562, N17561, N17560, N17559, N17558, N17557, N17556, N17555, N17554, N17553, N17552, N17551, N17550, N17549, N17548, N17547, N17546, N17545, N17544, N17543, N17542, N17541, N17540, N17539, N17538, N17537, N17536, N17535, N17534, N17533, N17532, N17531, N17530, N17529, N17528, N17527, N17526, N17525, N17524, N17523, N17522, N17521, N17520, N17519, N17518, N17517, N17516, N17515, N17514, N17513, N17512, N17511, N17510, N17509, N17508, N17507, N17506, N17505, N17504, N17503, N17502, N17501, N17500, N17499, N17498, N17497, N17496, N17495, N17494, N17493, N17492, N17491, N17490, N17489, N17488, N17487, N17486, N17485, N17484, N17483, N17482, N17481, N17480, N17479, N17478, N17477, N17476, N17475, N17474, N17473, N17472, N17471, N17470, N17469, N17468, N17467, N17466, N17465, N17464, N17463, N17462, N17461, N17460, N17459, N17458, N17457, N17456, N17455, N17454, N17453, N17452, N17451, N17450, N17449, N17448, N17447, N17446, N17445, N17444, N17443, N17442, N17441, N17440, N17439, N17438, N17437, N17436, N17435, N17434, N17433, N17432, N17431, N17430, N17429, N17428, N17427, N17426, N17425, N17424, N17423, N17422, N17421, N17420, N17419, N17418, N17417, N17416, N17415, N17414, N17413, N17412, N17411, N17410, N17409, N17408, N17407, N17406, N17405, N17404, N17403, N17402, N17401, N17400, N17399, N17398, N17397, N17396, N17395, N17394, N17393, N17392, N17391, N17390, N17389, N17388, N17387, N17386, N17385, N17384, N17383, N17382, N17381, N17380, N17379, N17378, N17377, N17376, N17375, N17374, N17373, N17372, N17371, N17370, N17369, N17368, N17367, N17366, N17365, N17364, N17363, N17362, N17361, N17360, N17359, N17358, N17357, N17356, N17355, N17354, N17353, N17352, N17351, N17350, N17349, N17348, N17347, N17346, N17345, N17344, N17343, N17342, N17341, N17340, N17339, N17338, N17337, N17336, N17335, N17334, N17333, N17332, N17331, N17330, N17329, N17328, N17327, N17326, N17325, N17324, N17323, N17322, N17321, N17320, N17319, N17318, N17317, N17316, N17315, N17314, N17313, N17312, N17311, N17310, N17309, N17308, N17307, N17306, N17305, N17304, N17303, N17302, N17301, N17300, N17299, N17298, N17297, N17296, N17295, N17294, N17293, N17292, N17291, N17290, N17289, N17288, N17287, N17286, N17285, N17284, N17283, N17282, N17281, N17280, N17279, N17278, N17277, N17276, N17275, N17274, N17273, N17272, N17271, N17270, N17269, N17268, N17267, N17266, N17265, N17264, N17263, N17262, N17261, N17260, N17259, N17258, N17257, N17256, N17255, N17254, N17253, N17252, N17251, N17250, N17249, N17248, N17247, N17246, N17245, N17244, N17243, N17242, N17241, N17240, N17239, N17238, N17237, N17236, N17235, N17234, N17233, N17232, N17231, N17230, N17229, N17228, N17227, N17226, N17225, N17224, N17223, N17222, N17221, N17220, N17219, N17218, N17217, N17216, N17215, N17214, N17213, N17212, N17211, N17210, N17209, N17208, N17207, N17206, N17205, N17204, N17203, N17202, N17201, N17200, N17199, N17198, N17197, N17196, N17195, N17194, N17193, N17192, N17191, N17190, N17189, N17188, N17187, N17186, N17185, N17184, N17183, N17182, N17181, N17180, N17179, N17178, N17177, N17176, N17175, N17174, N17173, N17172, N17171, N17170, N17169, N17168, N17167, N17166, N17165, N17164, N17163, N17162, N17161, N17160, N17159, N17158, N17157, N17156, N17155, N17154, N17153, N17152, N17151, N17150, N17149, N17148, N17147, N17146, N17145, N17144, N17143, N17142, N17141, N17140, N17139, N17138, N17137, N17136, N17135, N17134, N17133, N17132, N17131, N17130, N17129, N17128, N17127, N17126, N17125, N17124, N17123, N17122, N17121, N17120, N17119, N17118, N17117, N17116, N17115, N17114, N17113, N17112, N17111, N17110, N17109, N17108, N17107, N17106, N17105, N17104, N17103, N17102, N17101, N17100, N17099, N17098, N17097, N17096, N17095, N17094, N17093, N17092, N17091, N17090, N17089, N17088, N17087, N17086, N17085, N17084, N17083, N17082, N17081, N17080, N17079, N17078, N17077, N17076, N17075, N17074, N17073, N17072, N17071, N17070, N17069, N17068, N17067, N17066, N17065, N17064, N17063, N17062, N17061, N17060, N17059, N17058, N17057, N17056, N17055, N17054, N17053, N17052, N17051, N17050, N17049, N17048, N17047, N17046, N17045, N17044, N17043, N17042, N17041, N17040, N17039, N17038, N17037, N17036, N17035, N17034, N17033, N17032, N17031, N17030, N17029, N17028, N17027, N17026, N17025, N17024, N17023, N17022, N17021, N17020, N17019, N17018, N17017, N17016, N17015, N17014, N17013, N17012, N17011, N17010, N17009, N17008, N17007, N17006, N17005, N17004, N17003, N17002, N17001, N17000, N16999, N16998, N16997, N16996, N16995, N16994, N16993, N16992, N16991, N16990, N16989, N16988, N16987, N16986, N16985, N16984, N16983, N16982, N16981, N16980, N16979, N16978, N16977, N16976, N16975, N16974, N16973, N16972, N16971, N16970, N16969, N16968, N16967, N16966, N16965, N16964, N16963, N16962, N16961, N16960, N16959, N16958, N16957, N16956, N16955, N16954, N16953, N16952, N16951, N16950, N16949, N16948, N16947, N16946, N16945, N16944, N16943, N16942, N16941, N16940, N16939, N16938, N16937, N16936, N16935, N16934, N16933, N16932, N16931, N16930, N16929, N16928, N16927, N16926, N16925, N16924, N16923, N16922, N16921, N16920, N16919, N16918, N16917, N16916, N16915, N16914, N16913, N16912, N16911, N16910, N16909, N16908, N16907, N16906, N16905, N16904, N16903, N16902, N16901, N16900, N16899, N16898, N16897, N16896, N16895, N16894, N16893, N16892, N16891, N16890, N16889, N16888, N16887, N16886, N16885, N16884, N16883, N16882, N16881, N16880, N16879, N16878, N16877, N16876, N16875, N16874, N16873, N16872, N16871, N16870, N16869, N16868, N16867, N16866, N16865, N16864, N16863, N16862, N16861, N16860, N16859, N16858, N16857, N16856, N16855, N16854, N16853, N16852, N16851, N16850, N16849, N16848, N16847, N16846, N16845, N16844, N16843, N16842, N16841, N16840, N16839, N16838, N16837, N16836, N16835, N16834, N16833, N16832, N16831, N16830, N16829, N16828, N16827, N16826, N16825, N16824, N16823, N16822, N16821, N16820, N16819, N16818, N16817, N16816, N16815, N16814, N16813, N16812, N16811, N16810, N16809, N16808, N16807, N16806, N16805, N16804, N16803, N16802, N16801, N16800, N16799, N16798, N16797, N16796, N16795, N16794, N16793, N16792, N16791, N16790, N16789, N16788, N16787, N16786, N16785, N16784, N16783, N16782, N16781, N16780, N16779, N16778, N16777, N16776, N16775, N16774, N16773, N16772, N16771, N16770, N16769, N16768, N16767, N16766, N16765, N16764, N16763, N16762, N16761, N16760, N16759, N16758, N16757, N16756, N16755, N16754, N16753, N16752, N16751, N16750, N16749, N16748, N16747, N16746, N16745, N16744, N16743, N16742, N16741, N16740, N16739, N16738, N16737, N16736, N16735, N16734, N16733, N16732, N16731, N16730, N16729, N16728, N16727, N16726, N16725, N16724, N16723, N16722, N16721, N16720, N16719, N16718, N16717, N16716, N16715, N16714, N16713, N16712, N16711, N16710, N16709, N16708, N16707, N16706, N16705, N16704, N16703, N16702, N16701, N16700, N16699, N16698, N16697, N16696, N16695, N16694, N16693, N16692, N16691, N16690, N16689, N16688, N16687, N16686, N16685, N16684, N16683, N16682, N16681, N16680, N16679, N16678, N16677, N16676, N16675, N16674, N16673, N16672, N16671, N16670, N16669, N16668, N16667, N16666, N16665, N16664, N16663, N16662, N16661, N16660, N16659, N16658, N16657, N16656, N16655, N16654, N16653, N16652, N16651, N16650, N16649, N16648, N16647, N16646, N16645, N16644, N16643, N16642, N16641, N16640, N16639, N16638, N16637, N16636, N16635, N16634, N16633, N16632, N16631, N16630, N16629, N16628, N16627, N16626, N16625, N16624, N16623, N16622, N16621, N16620, N16619, N16618, N16617, N16616, N16615, N16614, N16613, N16612, N16611, N16610, N16609, N16608, N16607, N16606, N16605, N16604, N16603, N16602, N16601, N16600, N16599, N16598, N16597, N16596, N16595, N16594, N16593, N16592, N16591, N16590, N16589, N16588, N16587, N16586, N16585, N16584, N16583, N16582, N16581, N16580, N16579, N16578, N16577, N16576, N16575, N16574, N16573, N16572, N16571, N16570, N16569, N16568, N16567, N16566, N16565, N16564, N16563, N16562, N16561, N16560, N16559, N16558, N16557, N16556, N16555, N16554, N16553, N16552, N16551, N16550, N16549, N16548, N16547, N16546, N16545, N16544, N16543, N16542, N16541, N16540, N16539, N16538, N16537, N16536, N16535, N16534, N16533, N16532, N16531, N16530, N16529, N16528, N16527, N16526, N16525, N16524, N16523, N16522, N16521, N16520, N16519, N16518, N16517, N16516, N16515, N16514, N16513, N16512, N16511, N16510, N16509, N16508, N16507, N16506, N16505, N16504, N16503, N16502, N16501, N16500, N16499, N16498, N16497, N16496, N16495, N16494, N16493, N16492, N16491, N16490, N16489, N16488, N16487, N16486, N16485, N16484, N16483, N16482, N16481, N16480, N16479, N16478, N16477, N16476, N16475, N16474, N16473, N16472, N16471, N16470, N16469, N16468, N16467, N16466, N16465, N16464, N16463, N16462, N16461, N16460, N16459, N16458, N16457, N16456, N16455, N16454, N16453, N16452, N16451, N16450, N16449, N16448, N16447, N16446, N16445, N16444, N16443, N16442, N16441, N16440, N16439, N16438, N16437, N16436, N16435, N16434, N16433, N16432, N16431, N16430, N16429, N16428, N16427, N16426, N16425, N16424, N16423, N16422, N16421, N16420, N16419, N16418, N16417, N16416, N16415, N16414, N16413, N16412, N16411, N16410, N16409, N16408, N16407, N16406, N16405, N16404, N16403, N16402, N16401, N16400, N16399, N16398, N16397, N16396, N16395, N16394, N16393, N16392, N16391, N16390, N16389, N16388, N16387, N16386, N16385, N16384, N16383, N16382, N16381, N16380, N16379, N16378, N16377, N16376, N16375, N16374, N16373, N16372, N16371, N16370, N16369, N16368, N16367, N16366, N16365, N16364, N16363, N16362, N16361, N16360, N16359, N16358, N16357, N16356, N16355, N16354, N16353, N16352, N16351, N16350, N16349, N16348, N16347, N16346, N16345, N16344, N16343, N16342, N16341, N16340, N16339, N16338, N16337, N16336, N16335, N16334, N16333, N16332, N16331, N16330, N16329, N16328, N16327, N16326, N16325, N16324, N16323, N16322, N16321, N16320, N16319, N16318, N16317, N16316, N16315, N16314, N16313, N16312, N16311, N16310, N16309, N16308, N16307, N16306, N16305, N16304, N16303, N16302, N16301, N16300, N16299, N16298, N16297, N16296, N16295, N16294, N16293, N16292 } : 1'b0;
  assign N192 = N18372;
  assign N24609 = (N193)? 1'b1 : 
                  (N24625)? N22720 : 1'b0;
  assign N193 = N24617;
  assign N24610 = (N194)? 1'b1 : 
                  (N24690)? N22978 : 1'b0;
  assign N194 = N24618;
  assign N24611 = (N195)? 1'b1 : 
                  (N24755)? N23236 : 1'b0;
  assign N195 = N24619;
  assign N24612 = (N196)? 1'b1 : 
                  (N24820)? N23494 : 1'b0;
  assign N196 = N24620;
  assign N24613 = (N197)? 1'b1 : 
                  (N24885)? N23752 : 1'b0;
  assign N197 = N24621;
  assign N24614 = (N198)? 1'b1 : 
                  (N24950)? N24010 : 1'b0;
  assign N198 = N24622;
  assign N24615 = (N199)? 1'b1 : 
                  (N25015)? N24268 : 1'b0;
  assign N199 = N24623;
  assign N24616 = (N200)? 1'b1 : 
                  (N25080)? N24526 : 1'b0;
  assign N200 = N24624;
  assign { N24689, N24688, N24687, N24686, N24685, N24684, N24683, N24682, N24681, N24680, N24679, N24678, N24677, N24676, N24675, N24674, N24673, N24672, N24671, N24670, N24669, N24668, N24667, N24666, N24665, N24664, N24663, N24662, N24661, N24660, N24659, N24658, N24657, N24656, N24655, N24654, N24653, N24652, N24651, N24650, N24649, N24648, N24647, N24646, N24645, N24644, N24643, N24642, N24641, N24640, N24639, N24638, N24637, N24636, N24635, N24634, N24633, N24632, N24631, N24630, N24629, N24628, N24627, N24626 } = (N193)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24625)? { N22784, N22783, N22782, N22781, N22780, N22779, N22778, N22777, N22776, N22775, N22774, N22773, N22772, N22771, N22770, N22769, N22768, N22767, N22766, N22765, N22764, N22763, N22762, N22761, N22760, N22759, N22758, N22757, N22756, N22755, N22754, N22753, N22752, N22751, N22750, N22749, N22748, N22747, N22746, N22745, N22744, N22743, N22742, N22741, N22740, N22739, N22738, N22737, N22736, N22735, N22734, N22733, N22732, N22731, N22730, N22729, N22728, N22727, N22726, N22725, N22724, N22723, N22722, N22721 } : 1'b0;
  assign { N24754, N24753, N24752, N24751, N24750, N24749, N24748, N24747, N24746, N24745, N24744, N24743, N24742, N24741, N24740, N24739, N24738, N24737, N24736, N24735, N24734, N24733, N24732, N24731, N24730, N24729, N24728, N24727, N24726, N24725, N24724, N24723, N24722, N24721, N24720, N24719, N24718, N24717, N24716, N24715, N24714, N24713, N24712, N24711, N24710, N24709, N24708, N24707, N24706, N24705, N24704, N24703, N24702, N24701, N24700, N24699, N24698, N24697, N24696, N24695, N24694, N24693, N24692, N24691 } = (N194)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24690)? { N23042, N23041, N23040, N23039, N23038, N23037, N23036, N23035, N23034, N23033, N23032, N23031, N23030, N23029, N23028, N23027, N23026, N23025, N23024, N23023, N23022, N23021, N23020, N23019, N23018, N23017, N23016, N23015, N23014, N23013, N23012, N23011, N23010, N23009, N23008, N23007, N23006, N23005, N23004, N23003, N23002, N23001, N23000, N22999, N22998, N22997, N22996, N22995, N22994, N22993, N22992, N22991, N22990, N22989, N22988, N22987, N22986, N22985, N22984, N22983, N22982, N22981, N22980, N22979 } : 1'b0;
  assign { N24819, N24818, N24817, N24816, N24815, N24814, N24813, N24812, N24811, N24810, N24809, N24808, N24807, N24806, N24805, N24804, N24803, N24802, N24801, N24800, N24799, N24798, N24797, N24796, N24795, N24794, N24793, N24792, N24791, N24790, N24789, N24788, N24787, N24786, N24785, N24784, N24783, N24782, N24781, N24780, N24779, N24778, N24777, N24776, N24775, N24774, N24773, N24772, N24771, N24770, N24769, N24768, N24767, N24766, N24765, N24764, N24763, N24762, N24761, N24760, N24759, N24758, N24757, N24756 } = (N195)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24755)? { N23300, N23299, N23298, N23297, N23296, N23295, N23294, N23293, N23292, N23291, N23290, N23289, N23288, N23287, N23286, N23285, N23284, N23283, N23282, N23281, N23280, N23279, N23278, N23277, N23276, N23275, N23274, N23273, N23272, N23271, N23270, N23269, N23268, N23267, N23266, N23265, N23264, N23263, N23262, N23261, N23260, N23259, N23258, N23257, N23256, N23255, N23254, N23253, N23252, N23251, N23250, N23249, N23248, N23247, N23246, N23245, N23244, N23243, N23242, N23241, N23240, N23239, N23238, N23237 } : 1'b0;
  assign { N24884, N24883, N24882, N24881, N24880, N24879, N24878, N24877, N24876, N24875, N24874, N24873, N24872, N24871, N24870, N24869, N24868, N24867, N24866, N24865, N24864, N24863, N24862, N24861, N24860, N24859, N24858, N24857, N24856, N24855, N24854, N24853, N24852, N24851, N24850, N24849, N24848, N24847, N24846, N24845, N24844, N24843, N24842, N24841, N24840, N24839, N24838, N24837, N24836, N24835, N24834, N24833, N24832, N24831, N24830, N24829, N24828, N24827, N24826, N24825, N24824, N24823, N24822, N24821 } = (N196)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24820)? { N23558, N23557, N23556, N23555, N23554, N23553, N23552, N23551, N23550, N23549, N23548, N23547, N23546, N23545, N23544, N23543, N23542, N23541, N23540, N23539, N23538, N23537, N23536, N23535, N23534, N23533, N23532, N23531, N23530, N23529, N23528, N23527, N23526, N23525, N23524, N23523, N23522, N23521, N23520, N23519, N23518, N23517, N23516, N23515, N23514, N23513, N23512, N23511, N23510, N23509, N23508, N23507, N23506, N23505, N23504, N23503, N23502, N23501, N23500, N23499, N23498, N23497, N23496, N23495 } : 1'b0;
  assign { N24949, N24948, N24947, N24946, N24945, N24944, N24943, N24942, N24941, N24940, N24939, N24938, N24937, N24936, N24935, N24934, N24933, N24932, N24931, N24930, N24929, N24928, N24927, N24926, N24925, N24924, N24923, N24922, N24921, N24920, N24919, N24918, N24917, N24916, N24915, N24914, N24913, N24912, N24911, N24910, N24909, N24908, N24907, N24906, N24905, N24904, N24903, N24902, N24901, N24900, N24899, N24898, N24897, N24896, N24895, N24894, N24893, N24892, N24891, N24890, N24889, N24888, N24887, N24886 } = (N197)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24885)? { N23816, N23815, N23814, N23813, N23812, N23811, N23810, N23809, N23808, N23807, N23806, N23805, N23804, N23803, N23802, N23801, N23800, N23799, N23798, N23797, N23796, N23795, N23794, N23793, N23792, N23791, N23790, N23789, N23788, N23787, N23786, N23785, N23784, N23783, N23782, N23781, N23780, N23779, N23778, N23777, N23776, N23775, N23774, N23773, N23772, N23771, N23770, N23769, N23768, N23767, N23766, N23765, N23764, N23763, N23762, N23761, N23760, N23759, N23758, N23757, N23756, N23755, N23754, N23753 } : 1'b0;
  assign { N25014, N25013, N25012, N25011, N25010, N25009, N25008, N25007, N25006, N25005, N25004, N25003, N25002, N25001, N25000, N24999, N24998, N24997, N24996, N24995, N24994, N24993, N24992, N24991, N24990, N24989, N24988, N24987, N24986, N24985, N24984, N24983, N24982, N24981, N24980, N24979, N24978, N24977, N24976, N24975, N24974, N24973, N24972, N24971, N24970, N24969, N24968, N24967, N24966, N24965, N24964, N24963, N24962, N24961, N24960, N24959, N24958, N24957, N24956, N24955, N24954, N24953, N24952, N24951 } = (N198)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24950)? { N24074, N24073, N24072, N24071, N24070, N24069, N24068, N24067, N24066, N24065, N24064, N24063, N24062, N24061, N24060, N24059, N24058, N24057, N24056, N24055, N24054, N24053, N24052, N24051, N24050, N24049, N24048, N24047, N24046, N24045, N24044, N24043, N24042, N24041, N24040, N24039, N24038, N24037, N24036, N24035, N24034, N24033, N24032, N24031, N24030, N24029, N24028, N24027, N24026, N24025, N24024, N24023, N24022, N24021, N24020, N24019, N24018, N24017, N24016, N24015, N24014, N24013, N24012, N24011 } : 1'b0;
  assign { N25079, N25078, N25077, N25076, N25075, N25074, N25073, N25072, N25071, N25070, N25069, N25068, N25067, N25066, N25065, N25064, N25063, N25062, N25061, N25060, N25059, N25058, N25057, N25056, N25055, N25054, N25053, N25052, N25051, N25050, N25049, N25048, N25047, N25046, N25045, N25044, N25043, N25042, N25041, N25040, N25039, N25038, N25037, N25036, N25035, N25034, N25033, N25032, N25031, N25030, N25029, N25028, N25027, N25026, N25025, N25024, N25023, N25022, N25021, N25020, N25019, N25018, N25017, N25016 } = (N199)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25015)? { N24332, N24331, N24330, N24329, N24328, N24327, N24326, N24325, N24324, N24323, N24322, N24321, N24320, N24319, N24318, N24317, N24316, N24315, N24314, N24313, N24312, N24311, N24310, N24309, N24308, N24307, N24306, N24305, N24304, N24303, N24302, N24301, N24300, N24299, N24298, N24297, N24296, N24295, N24294, N24293, N24292, N24291, N24290, N24289, N24288, N24287, N24286, N24285, N24284, N24283, N24282, N24281, N24280, N24279, N24278, N24277, N24276, N24275, N24274, N24273, N24272, N24271, N24270, N24269 } : 1'b0;
  assign { N25144, N25143, N25142, N25141, N25140, N25139, N25138, N25137, N25136, N25135, N25134, N25133, N25132, N25131, N25130, N25129, N25128, N25127, N25126, N25125, N25124, N25123, N25122, N25121, N25120, N25119, N25118, N25117, N25116, N25115, N25114, N25113, N25112, N25111, N25110, N25109, N25108, N25107, N25106, N25105, N25104, N25103, N25102, N25101, N25100, N25099, N25098, N25097, N25096, N25095, N25094, N25093, N25092, N25091, N25090, N25089, N25088, N25087, N25086, N25085, N25084, N25083, N25082, N25081 } = (N200)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25080)? { N24590, N24589, N24588, N24587, N24586, N24585, N24584, N24583, N24582, N24581, N24580, N24579, N24578, N24577, N24576, N24575, N24574, N24573, N24572, N24571, N24570, N24569, N24568, N24567, N24566, N24565, N24564, N24563, N24562, N24561, N24560, N24559, N24558, N24557, N24556, N24555, N24554, N24553, N24552, N24551, N24550, N24549, N24548, N24547, N24546, N24545, N24544, N24543, N24542, N24541, N24540, N24539, N24538, N24537, N24536, N24535, N24534, N24533, N24532, N24531, N24530, N24529, N24528, N24527 } : 1'b0;
  assign { N25208, N25207, N25206, N25205, N25204, N25203, N25202, N25201, N25200, N25199, N25198, N25197, N25196, N25195, N25194, N25193, N25192, N25191, N25190, N25189, N25188, N25187, N25186, N25185, N25184, N25183, N25182, N25181, N25180, N25179, N25178, N25177, N25176, N25175, N25174, N25173, N25172, N25171, N25170, N25169, N25168, N25167, N25166, N25165, N25164, N25163, N25162, N25161, N25160, N25159, N25158, N25157, N25156, N25155, N25154, N25153, N25152, N25151, N25150, N25149, N25148, N25147, N25146, N25145 } = (N193)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24625)? { N22590, N22589, N22588, N22587, N22586, N22585, N22584, N22583, N22582, N22581, N22580, N22579, N22578, N22577, N22576, N22575, N22574, N22573, N22572, N22571, N22570, N22569, N22568, N22567, N22566, N22565, N22564, N22563, N22562, N22561, N22560, N22559, N22558, N22557, N22556, N22555, N22554, N22553, N22552, N22551, N22550, N22549, N22548, N22547, N22546, N22545, N22544, N22543, N22542, N22541, N22540, N22539, N22538, N22537, N22536, N22535, N22534, N22533, N22532, N22531, N22530, N22529, N22528, N22527 } : 1'b0;
  assign { N25272, N25271, N25270, N25269, N25268, N25267, N25266, N25265, N25264, N25263, N25262, N25261, N25260, N25259, N25258, N25257, N25256, N25255, N25254, N25253, N25252, N25251, N25250, N25249, N25248, N25247, N25246, N25245, N25244, N25243, N25242, N25241, N25240, N25239, N25238, N25237, N25236, N25235, N25234, N25233, N25232, N25231, N25230, N25229, N25228, N25227, N25226, N25225, N25224, N25223, N25222, N25221, N25220, N25219, N25218, N25217, N25216, N25215, N25214, N25213, N25212, N25211, N25210, N25209 } = (N194)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24690)? { N22848, N22847, N22846, N22845, N22844, N22843, N22842, N22841, N22840, N22839, N22838, N22837, N22836, N22835, N22834, N22833, N22832, N22831, N22830, N22829, N22828, N22827, N22826, N22825, N22824, N22823, N22822, N22821, N22820, N22819, N22818, N22817, N22816, N22815, N22814, N22813, N22812, N22811, N22810, N22809, N22808, N22807, N22806, N22805, N22804, N22803, N22802, N22801, N22800, N22799, N22798, N22797, N22796, N22795, N22794, N22793, N22792, N22791, N22790, N22789, N22788, N22787, N22786, N22785 } : 1'b0;
  assign { N25336, N25335, N25334, N25333, N25332, N25331, N25330, N25329, N25328, N25327, N25326, N25325, N25324, N25323, N25322, N25321, N25320, N25319, N25318, N25317, N25316, N25315, N25314, N25313, N25312, N25311, N25310, N25309, N25308, N25307, N25306, N25305, N25304, N25303, N25302, N25301, N25300, N25299, N25298, N25297, N25296, N25295, N25294, N25293, N25292, N25291, N25290, N25289, N25288, N25287, N25286, N25285, N25284, N25283, N25282, N25281, N25280, N25279, N25278, N25277, N25276, N25275, N25274, N25273 } = (N195)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24755)? { N23106, N23105, N23104, N23103, N23102, N23101, N23100, N23099, N23098, N23097, N23096, N23095, N23094, N23093, N23092, N23091, N23090, N23089, N23088, N23087, N23086, N23085, N23084, N23083, N23082, N23081, N23080, N23079, N23078, N23077, N23076, N23075, N23074, N23073, N23072, N23071, N23070, N23069, N23068, N23067, N23066, N23065, N23064, N23063, N23062, N23061, N23060, N23059, N23058, N23057, N23056, N23055, N23054, N23053, N23052, N23051, N23050, N23049, N23048, N23047, N23046, N23045, N23044, N23043 } : 1'b0;
  assign { N25400, N25399, N25398, N25397, N25396, N25395, N25394, N25393, N25392, N25391, N25390, N25389, N25388, N25387, N25386, N25385, N25384, N25383, N25382, N25381, N25380, N25379, N25378, N25377, N25376, N25375, N25374, N25373, N25372, N25371, N25370, N25369, N25368, N25367, N25366, N25365, N25364, N25363, N25362, N25361, N25360, N25359, N25358, N25357, N25356, N25355, N25354, N25353, N25352, N25351, N25350, N25349, N25348, N25347, N25346, N25345, N25344, N25343, N25342, N25341, N25340, N25339, N25338, N25337 } = (N196)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24820)? { N23364, N23363, N23362, N23361, N23360, N23359, N23358, N23357, N23356, N23355, N23354, N23353, N23352, N23351, N23350, N23349, N23348, N23347, N23346, N23345, N23344, N23343, N23342, N23341, N23340, N23339, N23338, N23337, N23336, N23335, N23334, N23333, N23332, N23331, N23330, N23329, N23328, N23327, N23326, N23325, N23324, N23323, N23322, N23321, N23320, N23319, N23318, N23317, N23316, N23315, N23314, N23313, N23312, N23311, N23310, N23309, N23308, N23307, N23306, N23305, N23304, N23303, N23302, N23301 } : 1'b0;
  assign { N25464, N25463, N25462, N25461, N25460, N25459, N25458, N25457, N25456, N25455, N25454, N25453, N25452, N25451, N25450, N25449, N25448, N25447, N25446, N25445, N25444, N25443, N25442, N25441, N25440, N25439, N25438, N25437, N25436, N25435, N25434, N25433, N25432, N25431, N25430, N25429, N25428, N25427, N25426, N25425, N25424, N25423, N25422, N25421, N25420, N25419, N25418, N25417, N25416, N25415, N25414, N25413, N25412, N25411, N25410, N25409, N25408, N25407, N25406, N25405, N25404, N25403, N25402, N25401 } = (N197)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24885)? { N23622, N23621, N23620, N23619, N23618, N23617, N23616, N23615, N23614, N23613, N23612, N23611, N23610, N23609, N23608, N23607, N23606, N23605, N23604, N23603, N23602, N23601, N23600, N23599, N23598, N23597, N23596, N23595, N23594, N23593, N23592, N23591, N23590, N23589, N23588, N23587, N23586, N23585, N23584, N23583, N23582, N23581, N23580, N23579, N23578, N23577, N23576, N23575, N23574, N23573, N23572, N23571, N23570, N23569, N23568, N23567, N23566, N23565, N23564, N23563, N23562, N23561, N23560, N23559 } : 1'b0;
  assign { N25528, N25527, N25526, N25525, N25524, N25523, N25522, N25521, N25520, N25519, N25518, N25517, N25516, N25515, N25514, N25513, N25512, N25511, N25510, N25509, N25508, N25507, N25506, N25505, N25504, N25503, N25502, N25501, N25500, N25499, N25498, N25497, N25496, N25495, N25494, N25493, N25492, N25491, N25490, N25489, N25488, N25487, N25486, N25485, N25484, N25483, N25482, N25481, N25480, N25479, N25478, N25477, N25476, N25475, N25474, N25473, N25472, N25471, N25470, N25469, N25468, N25467, N25466, N25465 } = (N198)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24950)? { N23880, N23879, N23878, N23877, N23876, N23875, N23874, N23873, N23872, N23871, N23870, N23869, N23868, N23867, N23866, N23865, N23864, N23863, N23862, N23861, N23860, N23859, N23858, N23857, N23856, N23855, N23854, N23853, N23852, N23851, N23850, N23849, N23848, N23847, N23846, N23845, N23844, N23843, N23842, N23841, N23840, N23839, N23838, N23837, N23836, N23835, N23834, N23833, N23832, N23831, N23830, N23829, N23828, N23827, N23826, N23825, N23824, N23823, N23822, N23821, N23820, N23819, N23818, N23817 } : 1'b0;
  assign { N25592, N25591, N25590, N25589, N25588, N25587, N25586, N25585, N25584, N25583, N25582, N25581, N25580, N25579, N25578, N25577, N25576, N25575, N25574, N25573, N25572, N25571, N25570, N25569, N25568, N25567, N25566, N25565, N25564, N25563, N25562, N25561, N25560, N25559, N25558, N25557, N25556, N25555, N25554, N25553, N25552, N25551, N25550, N25549, N25548, N25547, N25546, N25545, N25544, N25543, N25542, N25541, N25540, N25539, N25538, N25537, N25536, N25535, N25534, N25533, N25532, N25531, N25530, N25529 } = (N199)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25015)? { N24138, N24137, N24136, N24135, N24134, N24133, N24132, N24131, N24130, N24129, N24128, N24127, N24126, N24125, N24124, N24123, N24122, N24121, N24120, N24119, N24118, N24117, N24116, N24115, N24114, N24113, N24112, N24111, N24110, N24109, N24108, N24107, N24106, N24105, N24104, N24103, N24102, N24101, N24100, N24099, N24098, N24097, N24096, N24095, N24094, N24093, N24092, N24091, N24090, N24089, N24088, N24087, N24086, N24085, N24084, N24083, N24082, N24081, N24080, N24079, N24078, N24077, N24076, N24075 } : 1'b0;
  assign { N25656, N25655, N25654, N25653, N25652, N25651, N25650, N25649, N25648, N25647, N25646, N25645, N25644, N25643, N25642, N25641, N25640, N25639, N25638, N25637, N25636, N25635, N25634, N25633, N25632, N25631, N25630, N25629, N25628, N25627, N25626, N25625, N25624, N25623, N25622, N25621, N25620, N25619, N25618, N25617, N25616, N25615, N25614, N25613, N25612, N25611, N25610, N25609, N25608, N25607, N25606, N25605, N25604, N25603, N25602, N25601, N25600, N25599, N25598, N25597, N25596, N25595, N25594, N25593 } = (N200)? resolved_branch_i[69:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25080)? { N24396, N24395, N24394, N24393, N24392, N24391, N24390, N24389, N24388, N24387, N24386, N24385, N24384, N24383, N24382, N24381, N24380, N24379, N24378, N24377, N24376, N24375, N24374, N24373, N24372, N24371, N24370, N24369, N24368, N24367, N24366, N24365, N24364, N24363, N24362, N24361, N24360, N24359, N24358, N24357, N24356, N24355, N24354, N24353, N24352, N24351, N24350, N24349, N24348, N24347, N24346, N24345, N24344, N24343, N24342, N24341, N24340, N24339, N24338, N24337, N24336, N24335, N24334, N24333 } : 1'b0;
  assign { N25790, N25789, N25788, N25787, N25786, N25785, N25784, N25783, N25782, N25781, N25780, N25779, N25778, N25777, N25776, N25775, N25774, N25773, N25772, N25771, N25770, N25769, N25768, N25767, N25766, N25765, N25764, N25763, N25762, N25761, N25760, N25759, N25758, N25757, N25756, N25755, N25754, N25753, N25752, N25751, N25750, N25749, N25748, N25747, N25746, N25745, N25744, N25743, N25742, N25741, N25740, N25739, N25738, N25737, N25736, N25735, N25734, N25733, N25732, N25731, N25730, N25729, N25728, N25727, N25726, N25725, N25724, N25723, N25722, N25721, N25720, N25719, N25718, N25717, N25716, N25715, N25714, N25713, N25712, N25711, N25710, N25709, N25708, N25707, N25706, N25705, N25704, N25703, N25702, N25701, N25700, N25699, N25698, N25697, N25696, N25695, N25694, N25693, N25692, N25691, N25690, N25689, N25688, N25687, N25686, N25685, N25684, N25683, N25682, N25681, N25680, N25679, N25678, N25677, N25676, N25675, N25674, N25673, N25672, N25671, N25670, N25669, N25668, N25667, N25666, N25665, N25664, N25663, N25662 } = (N193)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N24625)? { N22719, N22718, N22717, N22716, N22715, N22714, N22713, N22712, N22711, N22710, N22709, N22708, N22707, N22706, N22705, N22704, N22703, N22702, N22701, N22700, N22699, N22698, N22697, N22696, N22695, N22694, N22693, N22692, N22691, N22690, N22689, N22688, N22687, N22686, N22685, N22684, N22683, N22682, N22681, N22680, N22679, N22678, N22677, N22676, N22675, N22674, N22673, N22672, N22671, N22670, N22669, N22668, N22667, N22666, N22665, N22664, N22663, N22662, N22661, N22660, N22659, N22658, N22657, N22656, N22655, N22654, N22653, N22652, N22651, N22650, N22649, N22648, N22647, N22646, N22645, N22644, N22643, N22642, N22641, N22640, N22639, N22638, N22637, N22636, N22635, N22634, N22633, N22632, N22631, N22630, N22629, N22628, N22627, N22626, N22625, N22624, N22623, N22622, N22621, N22620, N22619, N22618, N22617, N22616, N22615, N22614, N22613, N22612, N22611, N22610, N22609, N22608, N22607, N22606, N22605, N22604, N22603, N22602, N22601, N22600, N22599, N22598, N22597, N22596, N22595, N22594, N22593, N22592, N22591 } : 1'b0;
  assign { N25919, N25918, N25917, N25916, N25915, N25914, N25913, N25912, N25911, N25910, N25909, N25908, N25907, N25906, N25905, N25904, N25903, N25902, N25901, N25900, N25899, N25898, N25897, N25896, N25895, N25894, N25893, N25892, N25891, N25890, N25889, N25888, N25887, N25886, N25885, N25884, N25883, N25882, N25881, N25880, N25879, N25878, N25877, N25876, N25875, N25874, N25873, N25872, N25871, N25870, N25869, N25868, N25867, N25866, N25865, N25864, N25863, N25862, N25861, N25860, N25859, N25858, N25857, N25856, N25855, N25854, N25853, N25852, N25851, N25850, N25849, N25848, N25847, N25846, N25845, N25844, N25843, N25842, N25841, N25840, N25839, N25838, N25837, N25836, N25835, N25834, N25833, N25832, N25831, N25830, N25829, N25828, N25827, N25826, N25825, N25824, N25823, N25822, N25821, N25820, N25819, N25818, N25817, N25816, N25815, N25814, N25813, N25812, N25811, N25810, N25809, N25808, N25807, N25806, N25805, N25804, N25803, N25802, N25801, N25800, N25799, N25798, N25797, N25796, N25795, N25794, N25793, N25792, N25791 } = (N194)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N24690)? { N22977, N22976, N22975, N22974, N22973, N22972, N22971, N22970, N22969, N22968, N22967, N22966, N22965, N22964, N22963, N22962, N22961, N22960, N22959, N22958, N22957, N22956, N22955, N22954, N22953, N22952, N22951, N22950, N22949, N22948, N22947, N22946, N22945, N22944, N22943, N22942, N22941, N22940, N22939, N22938, N22937, N22936, N22935, N22934, N22933, N22932, N22931, N22930, N22929, N22928, N22927, N22926, N22925, N22924, N22923, N22922, N22921, N22920, N22919, N22918, N22917, N22916, N22915, N22914, N22913, N22912, N22911, N22910, N22909, N22908, N22907, N22906, N22905, N22904, N22903, N22902, N22901, N22900, N22899, N22898, N22897, N22896, N22895, N22894, N22893, N22892, N22891, N22890, N22889, N22888, N22887, N22886, N22885, N22884, N22883, N22882, N22881, N22880, N22879, N22878, N22877, N22876, N22875, N22874, N22873, N22872, N22871, N22870, N22869, N22868, N22867, N22866, N22865, N22864, N22863, N22862, N22861, N22860, N22859, N22858, N22857, N22856, N22855, N22854, N22853, N22852, N22851, N22850, N22849 } : 1'b0;
  assign { N26048, N26047, N26046, N26045, N26044, N26043, N26042, N26041, N26040, N26039, N26038, N26037, N26036, N26035, N26034, N26033, N26032, N26031, N26030, N26029, N26028, N26027, N26026, N26025, N26024, N26023, N26022, N26021, N26020, N26019, N26018, N26017, N26016, N26015, N26014, N26013, N26012, N26011, N26010, N26009, N26008, N26007, N26006, N26005, N26004, N26003, N26002, N26001, N26000, N25999, N25998, N25997, N25996, N25995, N25994, N25993, N25992, N25991, N25990, N25989, N25988, N25987, N25986, N25985, N25984, N25983, N25982, N25981, N25980, N25979, N25978, N25977, N25976, N25975, N25974, N25973, N25972, N25971, N25970, N25969, N25968, N25967, N25966, N25965, N25964, N25963, N25962, N25961, N25960, N25959, N25958, N25957, N25956, N25955, N25954, N25953, N25952, N25951, N25950, N25949, N25948, N25947, N25946, N25945, N25944, N25943, N25942, N25941, N25940, N25939, N25938, N25937, N25936, N25935, N25934, N25933, N25932, N25931, N25930, N25929, N25928, N25927, N25926, N25925, N25924, N25923, N25922, N25921, N25920 } = (N195)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N24755)? { N23235, N23234, N23233, N23232, N23231, N23230, N23229, N23228, N23227, N23226, N23225, N23224, N23223, N23222, N23221, N23220, N23219, N23218, N23217, N23216, N23215, N23214, N23213, N23212, N23211, N23210, N23209, N23208, N23207, N23206, N23205, N23204, N23203, N23202, N23201, N23200, N23199, N23198, N23197, N23196, N23195, N23194, N23193, N23192, N23191, N23190, N23189, N23188, N23187, N23186, N23185, N23184, N23183, N23182, N23181, N23180, N23179, N23178, N23177, N23176, N23175, N23174, N23173, N23172, N23171, N23170, N23169, N23168, N23167, N23166, N23165, N23164, N23163, N23162, N23161, N23160, N23159, N23158, N23157, N23156, N23155, N23154, N23153, N23152, N23151, N23150, N23149, N23148, N23147, N23146, N23145, N23144, N23143, N23142, N23141, N23140, N23139, N23138, N23137, N23136, N23135, N23134, N23133, N23132, N23131, N23130, N23129, N23128, N23127, N23126, N23125, N23124, N23123, N23122, N23121, N23120, N23119, N23118, N23117, N23116, N23115, N23114, N23113, N23112, N23111, N23110, N23109, N23108, N23107 } : 1'b0;
  assign { N26177, N26176, N26175, N26174, N26173, N26172, N26171, N26170, N26169, N26168, N26167, N26166, N26165, N26164, N26163, N26162, N26161, N26160, N26159, N26158, N26157, N26156, N26155, N26154, N26153, N26152, N26151, N26150, N26149, N26148, N26147, N26146, N26145, N26144, N26143, N26142, N26141, N26140, N26139, N26138, N26137, N26136, N26135, N26134, N26133, N26132, N26131, N26130, N26129, N26128, N26127, N26126, N26125, N26124, N26123, N26122, N26121, N26120, N26119, N26118, N26117, N26116, N26115, N26114, N26113, N26112, N26111, N26110, N26109, N26108, N26107, N26106, N26105, N26104, N26103, N26102, N26101, N26100, N26099, N26098, N26097, N26096, N26095, N26094, N26093, N26092, N26091, N26090, N26089, N26088, N26087, N26086, N26085, N26084, N26083, N26082, N26081, N26080, N26079, N26078, N26077, N26076, N26075, N26074, N26073, N26072, N26071, N26070, N26069, N26068, N26067, N26066, N26065, N26064, N26063, N26062, N26061, N26060, N26059, N26058, N26057, N26056, N26055, N26054, N26053, N26052, N26051, N26050, N26049 } = (N196)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N24820)? { N23493, N23492, N23491, N23490, N23489, N23488, N23487, N23486, N23485, N23484, N23483, N23482, N23481, N23480, N23479, N23478, N23477, N23476, N23475, N23474, N23473, N23472, N23471, N23470, N23469, N23468, N23467, N23466, N23465, N23464, N23463, N23462, N23461, N23460, N23459, N23458, N23457, N23456, N23455, N23454, N23453, N23452, N23451, N23450, N23449, N23448, N23447, N23446, N23445, N23444, N23443, N23442, N23441, N23440, N23439, N23438, N23437, N23436, N23435, N23434, N23433, N23432, N23431, N23430, N23429, N23428, N23427, N23426, N23425, N23424, N23423, N23422, N23421, N23420, N23419, N23418, N23417, N23416, N23415, N23414, N23413, N23412, N23411, N23410, N23409, N23408, N23407, N23406, N23405, N23404, N23403, N23402, N23401, N23400, N23399, N23398, N23397, N23396, N23395, N23394, N23393, N23392, N23391, N23390, N23389, N23388, N23387, N23386, N23385, N23384, N23383, N23382, N23381, N23380, N23379, N23378, N23377, N23376, N23375, N23374, N23373, N23372, N23371, N23370, N23369, N23368, N23367, N23366, N23365 } : 1'b0;
  assign { N26306, N26305, N26304, N26303, N26302, N26301, N26300, N26299, N26298, N26297, N26296, N26295, N26294, N26293, N26292, N26291, N26290, N26289, N26288, N26287, N26286, N26285, N26284, N26283, N26282, N26281, N26280, N26279, N26278, N26277, N26276, N26275, N26274, N26273, N26272, N26271, N26270, N26269, N26268, N26267, N26266, N26265, N26264, N26263, N26262, N26261, N26260, N26259, N26258, N26257, N26256, N26255, N26254, N26253, N26252, N26251, N26250, N26249, N26248, N26247, N26246, N26245, N26244, N26243, N26242, N26241, N26240, N26239, N26238, N26237, N26236, N26235, N26234, N26233, N26232, N26231, N26230, N26229, N26228, N26227, N26226, N26225, N26224, N26223, N26222, N26221, N26220, N26219, N26218, N26217, N26216, N26215, N26214, N26213, N26212, N26211, N26210, N26209, N26208, N26207, N26206, N26205, N26204, N26203, N26202, N26201, N26200, N26199, N26198, N26197, N26196, N26195, N26194, N26193, N26192, N26191, N26190, N26189, N26188, N26187, N26186, N26185, N26184, N26183, N26182, N26181, N26180, N26179, N26178 } = (N197)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N24885)? { N23751, N23750, N23749, N23748, N23747, N23746, N23745, N23744, N23743, N23742, N23741, N23740, N23739, N23738, N23737, N23736, N23735, N23734, N23733, N23732, N23731, N23730, N23729, N23728, N23727, N23726, N23725, N23724, N23723, N23722, N23721, N23720, N23719, N23718, N23717, N23716, N23715, N23714, N23713, N23712, N23711, N23710, N23709, N23708, N23707, N23706, N23705, N23704, N23703, N23702, N23701, N23700, N23699, N23698, N23697, N23696, N23695, N23694, N23693, N23692, N23691, N23690, N23689, N23688, N23687, N23686, N23685, N23684, N23683, N23682, N23681, N23680, N23679, N23678, N23677, N23676, N23675, N23674, N23673, N23672, N23671, N23670, N23669, N23668, N23667, N23666, N23665, N23664, N23663, N23662, N23661, N23660, N23659, N23658, N23657, N23656, N23655, N23654, N23653, N23652, N23651, N23650, N23649, N23648, N23647, N23646, N23645, N23644, N23643, N23642, N23641, N23640, N23639, N23638, N23637, N23636, N23635, N23634, N23633, N23632, N23631, N23630, N23629, N23628, N23627, N23626, N23625, N23624, N23623 } : 1'b0;
  assign { N26435, N26434, N26433, N26432, N26431, N26430, N26429, N26428, N26427, N26426, N26425, N26424, N26423, N26422, N26421, N26420, N26419, N26418, N26417, N26416, N26415, N26414, N26413, N26412, N26411, N26410, N26409, N26408, N26407, N26406, N26405, N26404, N26403, N26402, N26401, N26400, N26399, N26398, N26397, N26396, N26395, N26394, N26393, N26392, N26391, N26390, N26389, N26388, N26387, N26386, N26385, N26384, N26383, N26382, N26381, N26380, N26379, N26378, N26377, N26376, N26375, N26374, N26373, N26372, N26371, N26370, N26369, N26368, N26367, N26366, N26365, N26364, N26363, N26362, N26361, N26360, N26359, N26358, N26357, N26356, N26355, N26354, N26353, N26352, N26351, N26350, N26349, N26348, N26347, N26346, N26345, N26344, N26343, N26342, N26341, N26340, N26339, N26338, N26337, N26336, N26335, N26334, N26333, N26332, N26331, N26330, N26329, N26328, N26327, N26326, N26325, N26324, N26323, N26322, N26321, N26320, N26319, N26318, N26317, N26316, N26315, N26314, N26313, N26312, N26311, N26310, N26309, N26308, N26307 } = (N198)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N24950)? { N24009, N24008, N24007, N24006, N24005, N24004, N24003, N24002, N24001, N24000, N23999, N23998, N23997, N23996, N23995, N23994, N23993, N23992, N23991, N23990, N23989, N23988, N23987, N23986, N23985, N23984, N23983, N23982, N23981, N23980, N23979, N23978, N23977, N23976, N23975, N23974, N23973, N23972, N23971, N23970, N23969, N23968, N23967, N23966, N23965, N23964, N23963, N23962, N23961, N23960, N23959, N23958, N23957, N23956, N23955, N23954, N23953, N23952, N23951, N23950, N23949, N23948, N23947, N23946, N23945, N23944, N23943, N23942, N23941, N23940, N23939, N23938, N23937, N23936, N23935, N23934, N23933, N23932, N23931, N23930, N23929, N23928, N23927, N23926, N23925, N23924, N23923, N23922, N23921, N23920, N23919, N23918, N23917, N23916, N23915, N23914, N23913, N23912, N23911, N23910, N23909, N23908, N23907, N23906, N23905, N23904, N23903, N23902, N23901, N23900, N23899, N23898, N23897, N23896, N23895, N23894, N23893, N23892, N23891, N23890, N23889, N23888, N23887, N23886, N23885, N23884, N23883, N23882, N23881 } : 1'b0;
  assign { N26564, N26563, N26562, N26561, N26560, N26559, N26558, N26557, N26556, N26555, N26554, N26553, N26552, N26551, N26550, N26549, N26548, N26547, N26546, N26545, N26544, N26543, N26542, N26541, N26540, N26539, N26538, N26537, N26536, N26535, N26534, N26533, N26532, N26531, N26530, N26529, N26528, N26527, N26526, N26525, N26524, N26523, N26522, N26521, N26520, N26519, N26518, N26517, N26516, N26515, N26514, N26513, N26512, N26511, N26510, N26509, N26508, N26507, N26506, N26505, N26504, N26503, N26502, N26501, N26500, N26499, N26498, N26497, N26496, N26495, N26494, N26493, N26492, N26491, N26490, N26489, N26488, N26487, N26486, N26485, N26484, N26483, N26482, N26481, N26480, N26479, N26478, N26477, N26476, N26475, N26474, N26473, N26472, N26471, N26470, N26469, N26468, N26467, N26466, N26465, N26464, N26463, N26462, N26461, N26460, N26459, N26458, N26457, N26456, N26455, N26454, N26453, N26452, N26451, N26450, N26449, N26448, N26447, N26446, N26445, N26444, N26443, N26442, N26441, N26440, N26439, N26438, N26437, N26436 } = (N199)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N25015)? { N24267, N24266, N24265, N24264, N24263, N24262, N24261, N24260, N24259, N24258, N24257, N24256, N24255, N24254, N24253, N24252, N24251, N24250, N24249, N24248, N24247, N24246, N24245, N24244, N24243, N24242, N24241, N24240, N24239, N24238, N24237, N24236, N24235, N24234, N24233, N24232, N24231, N24230, N24229, N24228, N24227, N24226, N24225, N24224, N24223, N24222, N24221, N24220, N24219, N24218, N24217, N24216, N24215, N24214, N24213, N24212, N24211, N24210, N24209, N24208, N24207, N24206, N24205, N24204, N24203, N24202, N24201, N24200, N24199, N24198, N24197, N24196, N24195, N24194, N24193, N24192, N24191, N24190, N24189, N24188, N24187, N24186, N24185, N24184, N24183, N24182, N24181, N24180, N24179, N24178, N24177, N24176, N24175, N24174, N24173, N24172, N24171, N24170, N24169, N24168, N24167, N24166, N24165, N24164, N24163, N24162, N24161, N24160, N24159, N24158, N24157, N24156, N24155, N24154, N24153, N24152, N24151, N24150, N24149, N24148, N24147, N24146, N24145, N24144, N24143, N24142, N24141, N24140, N24139 } : 1'b0;
  assign { N26693, N26692, N26691, N26690, N26689, N26688, N26687, N26686, N26685, N26684, N26683, N26682, N26681, N26680, N26679, N26678, N26677, N26676, N26675, N26674, N26673, N26672, N26671, N26670, N26669, N26668, N26667, N26666, N26665, N26664, N26663, N26662, N26661, N26660, N26659, N26658, N26657, N26656, N26655, N26654, N26653, N26652, N26651, N26650, N26649, N26648, N26647, N26646, N26645, N26644, N26643, N26642, N26641, N26640, N26639, N26638, N26637, N26636, N26635, N26634, N26633, N26632, N26631, N26630, N26629, N26628, N26627, N26626, N26625, N26624, N26623, N26622, N26621, N26620, N26619, N26618, N26617, N26616, N26615, N26614, N26613, N26612, N26611, N26610, N26609, N26608, N26607, N26606, N26605, N26604, N26603, N26602, N26601, N26600, N26599, N26598, N26597, N26596, N26595, N26594, N26593, N26592, N26591, N26590, N26589, N26588, N26587, N26586, N26585, N26584, N26583, N26582, N26581, N26580, N26579, N26578, N26577, N26576, N26575, N26574, N26573, N26572, N26571, N26570, N26569, N26568, N26567, N26566, N26565 } = (N200)? ex_i[515:387] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N25080)? { N24525, N24524, N24523, N24522, N24521, N24520, N24519, N24518, N24517, N24516, N24515, N24514, N24513, N24512, N24511, N24510, N24509, N24508, N24507, N24506, N24505, N24504, N24503, N24502, N24501, N24500, N24499, N24498, N24497, N24496, N24495, N24494, N24493, N24492, N24491, N24490, N24489, N24488, N24487, N24486, N24485, N24484, N24483, N24482, N24481, N24480, N24479, N24478, N24477, N24476, N24475, N24474, N24473, N24472, N24471, N24470, N24469, N24468, N24467, N24466, N24465, N24464, N24463, N24462, N24461, N24460, N24459, N24458, N24457, N24456, N24455, N24454, N24453, N24452, N24451, N24450, N24449, N24448, N24447, N24446, N24445, N24444, N24443, N24442, N24441, N24440, N24439, N24438, N24437, N24436, N24435, N24434, N24433, N24432, N24431, N24430, N24429, N24428, N24427, N24426, N24425, N24424, N24423, N24422, N24421, N24420, N24419, N24418, N24417, N24416, N24415, N24414, N24413, N24412, N24411, N24410, N24409, N24408, N24407, N24406, N24405, N24404, N24403, N24402, N24401, N24400, N24399, N24398, N24397 } : 1'b0;
  assign { N26769, N26768, N26767, N26766, N26765, N26764, N26763, N26762, N26761, N26760, N26759, N26758, N26757, N26756, N26755, N26754, N26753, N26752, N26751, N26750, N26749, N26748, N26747, N26746, N26745, N26744, N26743, N26742, N26741, N26740, N26739, N26738, N26737, N26736, N26735, N26734, N26733, N26732, N26731, N26730, N26729, N26728, N26727, N26726, N26725, N26724, N26723, N26722, N26721, N26720, N26719, N26718, N26717, N26716, N26715, N26714, N26713, N26712, N26711, N26710, N26709, N26708, N26707, N26706 } = (N193)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24625)? { N22719, N22718, N22717, N22716, N22715, N22714, N22713, N22712, N22711, N22710, N22709, N22708, N22707, N22706, N22705, N22704, N22703, N22702, N22701, N22700, N22699, N22698, N22697, N22696, N22695, N22694, N22693, N22692, N22691, N22690, N22689, N22688, N22687, N22686, N22685, N22684, N22683, N22682, N22681, N22680, N22679, N22678, N22677, N22676, N22675, N22674, N22673, N22672, N22671, N22670, N22669, N22668, N22667, N22666, N22665, N22664, N22663, N22662, N22661, N22660, N22659, N22658, N22657, N22656 } : 1'b0;
  assign { N26833, N26832, N26831, N26830, N26829, N26828, N26827, N26826, N26825, N26824, N26823, N26822, N26821, N26820, N26819, N26818, N26817, N26816, N26815, N26814, N26813, N26812, N26811, N26810, N26809, N26808, N26807, N26806, N26805, N26804, N26803, N26802, N26801, N26800, N26799, N26798, N26797, N26796, N26795, N26794, N26793, N26792, N26791, N26790, N26789, N26788, N26787, N26786, N26785, N26784, N26783, N26782, N26781, N26780, N26779, N26778, N26777, N26776, N26775, N26774, N26773, N26772, N26771, N26770 } = (N194)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24690)? { N22977, N22976, N22975, N22974, N22973, N22972, N22971, N22970, N22969, N22968, N22967, N22966, N22965, N22964, N22963, N22962, N22961, N22960, N22959, N22958, N22957, N22956, N22955, N22954, N22953, N22952, N22951, N22950, N22949, N22948, N22947, N22946, N22945, N22944, N22943, N22942, N22941, N22940, N22939, N22938, N22937, N22936, N22935, N22934, N22933, N22932, N22931, N22930, N22929, N22928, N22927, N22926, N22925, N22924, N22923, N22922, N22921, N22920, N22919, N22918, N22917, N22916, N22915, N22914 } : 1'b0;
  assign { N26897, N26896, N26895, N26894, N26893, N26892, N26891, N26890, N26889, N26888, N26887, N26886, N26885, N26884, N26883, N26882, N26881, N26880, N26879, N26878, N26877, N26876, N26875, N26874, N26873, N26872, N26871, N26870, N26869, N26868, N26867, N26866, N26865, N26864, N26863, N26862, N26861, N26860, N26859, N26858, N26857, N26856, N26855, N26854, N26853, N26852, N26851, N26850, N26849, N26848, N26847, N26846, N26845, N26844, N26843, N26842, N26841, N26840, N26839, N26838, N26837, N26836, N26835, N26834 } = (N195)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24755)? { N23235, N23234, N23233, N23232, N23231, N23230, N23229, N23228, N23227, N23226, N23225, N23224, N23223, N23222, N23221, N23220, N23219, N23218, N23217, N23216, N23215, N23214, N23213, N23212, N23211, N23210, N23209, N23208, N23207, N23206, N23205, N23204, N23203, N23202, N23201, N23200, N23199, N23198, N23197, N23196, N23195, N23194, N23193, N23192, N23191, N23190, N23189, N23188, N23187, N23186, N23185, N23184, N23183, N23182, N23181, N23180, N23179, N23178, N23177, N23176, N23175, N23174, N23173, N23172 } : 1'b0;
  assign { N26961, N26960, N26959, N26958, N26957, N26956, N26955, N26954, N26953, N26952, N26951, N26950, N26949, N26948, N26947, N26946, N26945, N26944, N26943, N26942, N26941, N26940, N26939, N26938, N26937, N26936, N26935, N26934, N26933, N26932, N26931, N26930, N26929, N26928, N26927, N26926, N26925, N26924, N26923, N26922, N26921, N26920, N26919, N26918, N26917, N26916, N26915, N26914, N26913, N26912, N26911, N26910, N26909, N26908, N26907, N26906, N26905, N26904, N26903, N26902, N26901, N26900, N26899, N26898 } = (N196)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24820)? { N23493, N23492, N23491, N23490, N23489, N23488, N23487, N23486, N23485, N23484, N23483, N23482, N23481, N23480, N23479, N23478, N23477, N23476, N23475, N23474, N23473, N23472, N23471, N23470, N23469, N23468, N23467, N23466, N23465, N23464, N23463, N23462, N23461, N23460, N23459, N23458, N23457, N23456, N23455, N23454, N23453, N23452, N23451, N23450, N23449, N23448, N23447, N23446, N23445, N23444, N23443, N23442, N23441, N23440, N23439, N23438, N23437, N23436, N23435, N23434, N23433, N23432, N23431, N23430 } : 1'b0;
  assign { N27025, N27024, N27023, N27022, N27021, N27020, N27019, N27018, N27017, N27016, N27015, N27014, N27013, N27012, N27011, N27010, N27009, N27008, N27007, N27006, N27005, N27004, N27003, N27002, N27001, N27000, N26999, N26998, N26997, N26996, N26995, N26994, N26993, N26992, N26991, N26990, N26989, N26988, N26987, N26986, N26985, N26984, N26983, N26982, N26981, N26980, N26979, N26978, N26977, N26976, N26975, N26974, N26973, N26972, N26971, N26970, N26969, N26968, N26967, N26966, N26965, N26964, N26963, N26962 } = (N197)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24885)? { N23751, N23750, N23749, N23748, N23747, N23746, N23745, N23744, N23743, N23742, N23741, N23740, N23739, N23738, N23737, N23736, N23735, N23734, N23733, N23732, N23731, N23730, N23729, N23728, N23727, N23726, N23725, N23724, N23723, N23722, N23721, N23720, N23719, N23718, N23717, N23716, N23715, N23714, N23713, N23712, N23711, N23710, N23709, N23708, N23707, N23706, N23705, N23704, N23703, N23702, N23701, N23700, N23699, N23698, N23697, N23696, N23695, N23694, N23693, N23692, N23691, N23690, N23689, N23688 } : 1'b0;
  assign { N27089, N27088, N27087, N27086, N27085, N27084, N27083, N27082, N27081, N27080, N27079, N27078, N27077, N27076, N27075, N27074, N27073, N27072, N27071, N27070, N27069, N27068, N27067, N27066, N27065, N27064, N27063, N27062, N27061, N27060, N27059, N27058, N27057, N27056, N27055, N27054, N27053, N27052, N27051, N27050, N27049, N27048, N27047, N27046, N27045, N27044, N27043, N27042, N27041, N27040, N27039, N27038, N27037, N27036, N27035, N27034, N27033, N27032, N27031, N27030, N27029, N27028, N27027, N27026 } = (N198)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24950)? { N24009, N24008, N24007, N24006, N24005, N24004, N24003, N24002, N24001, N24000, N23999, N23998, N23997, N23996, N23995, N23994, N23993, N23992, N23991, N23990, N23989, N23988, N23987, N23986, N23985, N23984, N23983, N23982, N23981, N23980, N23979, N23978, N23977, N23976, N23975, N23974, N23973, N23972, N23971, N23970, N23969, N23968, N23967, N23966, N23965, N23964, N23963, N23962, N23961, N23960, N23959, N23958, N23957, N23956, N23955, N23954, N23953, N23952, N23951, N23950, N23949, N23948, N23947, N23946 } : 1'b0;
  assign { N27153, N27152, N27151, N27150, N27149, N27148, N27147, N27146, N27145, N27144, N27143, N27142, N27141, N27140, N27139, N27138, N27137, N27136, N27135, N27134, N27133, N27132, N27131, N27130, N27129, N27128, N27127, N27126, N27125, N27124, N27123, N27122, N27121, N27120, N27119, N27118, N27117, N27116, N27115, N27114, N27113, N27112, N27111, N27110, N27109, N27108, N27107, N27106, N27105, N27104, N27103, N27102, N27101, N27100, N27099, N27098, N27097, N27096, N27095, N27094, N27093, N27092, N27091, N27090 } = (N199)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25015)? { N24267, N24266, N24265, N24264, N24263, N24262, N24261, N24260, N24259, N24258, N24257, N24256, N24255, N24254, N24253, N24252, N24251, N24250, N24249, N24248, N24247, N24246, N24245, N24244, N24243, N24242, N24241, N24240, N24239, N24238, N24237, N24236, N24235, N24234, N24233, N24232, N24231, N24230, N24229, N24228, N24227, N24226, N24225, N24224, N24223, N24222, N24221, N24220, N24219, N24218, N24217, N24216, N24215, N24214, N24213, N24212, N24211, N24210, N24209, N24208, N24207, N24206, N24205, N24204 } : 1'b0;
  assign { N27217, N27216, N27215, N27214, N27213, N27212, N27211, N27210, N27209, N27208, N27207, N27206, N27205, N27204, N27203, N27202, N27201, N27200, N27199, N27198, N27197, N27196, N27195, N27194, N27193, N27192, N27191, N27190, N27189, N27188, N27187, N27186, N27185, N27184, N27183, N27182, N27181, N27180, N27179, N27178, N27177, N27176, N27175, N27174, N27173, N27172, N27171, N27170, N27169, N27168, N27167, N27166, N27165, N27164, N27163, N27162, N27161, N27160, N27159, N27158, N27157, N27156, N27155, N27154 } = (N200)? ex_i[515:452] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25080)? { N24525, N24524, N24523, N24522, N24521, N24520, N24519, N24518, N24517, N24516, N24515, N24514, N24513, N24512, N24511, N24510, N24509, N24508, N24507, N24506, N24505, N24504, N24503, N24502, N24501, N24500, N24499, N24498, N24497, N24496, N24495, N24494, N24493, N24492, N24491, N24490, N24489, N24488, N24487, N24486, N24485, N24484, N24483, N24482, N24481, N24480, N24479, N24478, N24477, N24476, N24475, N24474, N24473, N24472, N24471, N24470, N24469, N24468, N24467, N24466, N24465, N24464, N24463, N24462 } : 1'b0;
  assign { N27729, N27728, N27727, N27726, N27725, N27724, N27723, N27722, N27721, N27720, N27719, N27718, N27717, N27716, N27715, N27714, N27713, N27712, N27711, N27710, N27709, N27708, N27707, N27706, N27705, N27704, N27703, N27702, N27701, N27700, N27699, N27698, N27697, N27696, N27695, N27694, N27693, N27692, N27691, N27690, N27689, N27688, N27687, N27686, N27685, N27684, N27683, N27682, N27681, N27680, N27679, N27678, N27677, N27676, N27675, N27674, N27673, N27672, N27671, N27670, N27669, N27668, N27667, N27666, N27665, N27664, N27663, N27662, N27661, N27660, N27659, N27658, N27657, N27656, N27655, N27654, N27653, N27652, N27651, N27650, N27649, N27648, N27647, N27646, N27645, N27644, N27643, N27642, N27641, N27640, N27639, N27638, N27637, N27636, N27635, N27634, N27633, N27632, N27631, N27630, N27629, N27628, N27627, N27626, N27625, N27624, N27623, N27622, N27621, N27620, N27619, N27618, N27617, N27616, N27615, N27614, N27613, N27612, N27611, N27610, N27609, N27608, N27607, N27606, N27605, N27604, N27603, N27602, N27601, N27600, N27599, N27598, N27597, N27596, N27595, N27594, N27593, N27592, N27591, N27590, N27589, N27588, N27587, N27586, N27585, N27584, N27583, N27582, N27581, N27580, N27579, N27578, N27577, N27576, N27575, N27574, N27573, N27572, N27571, N27570, N27569, N27568, N27567, N27566, N27565, N27564, N27563, N27562, N27561, N27560, N27559, N27558, N27557, N27556, N27555, N27554, N27553, N27552, N27551, N27550, N27549, N27548, N27547, N27546, N27545, N27544, N27543, N27542, N27541, N27540, N27539, N27538, N27537, N27536, N27535, N27534, N27533, N27532, N27531, N27530, N27529, N27528, N27527, N27526, N27525, N27524, N27523, N27522, N27521, N27520, N27519, N27518, N27517, N27516, N27515, N27514, N27513, N27512, N27511, N27510, N27509, N27508, N27507, N27506, N27505, N27504, N27503, N27502, N27501, N27500, N27499, N27498, N27497, N27496, N27495, N27494, N27493, N27492, N27491, N27490, N27489, N27488, N27487, N27486, N27485, N27484, N27483, N27482, N27481, N27480, N27479, N27478, N27477, N27476, N27475, N27474, N27473, N27472, N27471, N27470, N27469, N27468, N27467, N27466, N27465, N27464, N27463, N27462, N27461, N27460, N27459, N27458, N27457, N27456, N27455, N27454, N27453, N27452, N27451, N27450, N27449, N27448, N27447, N27446, N27445, N27444, N27443, N27442, N27441, N27440, N27439, N27438, N27437, N27436, N27435, N27434, N27433, N27432, N27431, N27430, N27429, N27428, N27427, N27426, N27425, N27424, N27423, N27422, N27421, N27420, N27419, N27418, N27417, N27416, N27415, N27414, N27413, N27412, N27411, N27410, N27409, N27408, N27407, N27406, N27405, N27404, N27403, N27402, N27401, N27400, N27399, N27398, N27397, N27396, N27395, N27394, N27393, N27392, N27391, N27390, N27389, N27388, N27387, N27386, N27385, N27384, N27383, N27382, N27381, N27380, N27379, N27378, N27377, N27376, N27375, N27374, N27373, N27372, N27371, N27370, N27369, N27368, N27367, N27366, N27365, N27364, N27363, N27362, N27361, N27360, N27359, N27358, N27357, N27356, N27355, N27354, N27353, N27352, N27351, N27350, N27349, N27348, N27347, N27346, N27345, N27344, N27343, N27342, N27341, N27340, N27339, N27338, N27337, N27336, N27335, N27334, N27333, N27332, N27331, N27330, N27329, N27328, N27327, N27326, N27325, N27324, N27323, N27322, N27321, N27320, N27319, N27318, N27317, N27316, N27315, N27314, N27313, N27312, N27311, N27310, N27309, N27308, N27307, N27306, N27305, N27304, N27303, N27302, N27301, N27300, N27299, N27298, N27297, N27296, N27295, N27294, N27293, N27292, N27291, N27290, N27289, N27288, N27287, N27286, N27285, N27284, N27283, N27282, N27281, N27280, N27279, N27278, N27277, N27276, N27275, N27274, N27273, N27272, N27271, N27270, N27269, N27268, N27267, N27266, N27265, N27264, N27263, N27262, N27261, N27260, N27259, N27258, N27257, N27256, N27255, N27254, N27253, N27252, N27251, N27250, N27249, N27248, N27247, N27246, N27245, N27244, N27243, N27242, N27241, N27240, N27239, N27238, N27237, N27236, N27235, N27234, N27233, N27232, N27231, N27230, N27229, N27228, N27227, N27226, N27225, N27224, N27223, N27222, N27221, N27220, N27219, N27218 } = (N201)? { N27217, N27216, N27215, N27214, N27213, N27212, N27211, N27210, N27209, N27208, N27207, N27206, N27205, N27204, N27203, N27202, N27201, N27200, N27199, N27198, N27197, N27196, N27195, N27194, N27193, N27192, N27191, N27190, N27189, N27188, N27187, N27186, N27185, N27184, N27183, N27182, N27181, N27180, N27179, N27178, N27177, N27176, N27175, N27174, N27173, N27172, N27171, N27170, N27169, N27168, N27167, N27166, N27165, N27164, N27163, N27162, N27161, N27160, N27159, N27158, N27157, N27156, N27155, N27154, N27153, N27152, N27151, N27150, N27149, N27148, N27147, N27146, N27145, N27144, N27143, N27142, N27141, N27140, N27139, N27138, N27137, N27136, N27135, N27134, N27133, N27132, N27131, N27130, N27129, N27128, N27127, N27126, N27125, N27124, N27123, N27122, N27121, N27120, N27119, N27118, N27117, N27116, N27115, N27114, N27113, N27112, N27111, N27110, N27109, N27108, N27107, N27106, N27105, N27104, N27103, N27102, N27101, N27100, N27099, N27098, N27097, N27096, N27095, N27094, N27093, N27092, N27091, N27090, N27089, N27088, N27087, N27086, N27085, N27084, N27083, N27082, N27081, N27080, N27079, N27078, N27077, N27076, N27075, N27074, N27073, N27072, N27071, N27070, N27069, N27068, N27067, N27066, N27065, N27064, N27063, N27062, N27061, N27060, N27059, N27058, N27057, N27056, N27055, N27054, N27053, N27052, N27051, N27050, N27049, N27048, N27047, N27046, N27045, N27044, N27043, N27042, N27041, N27040, N27039, N27038, N27037, N27036, N27035, N27034, N27033, N27032, N27031, N27030, N27029, N27028, N27027, N27026, N27025, N27024, N27023, N27022, N27021, N27020, N27019, N27018, N27017, N27016, N27015, N27014, N27013, N27012, N27011, N27010, N27009, N27008, N27007, N27006, N27005, N27004, N27003, N27002, N27001, N27000, N26999, N26998, N26997, N26996, N26995, N26994, N26993, N26992, N26991, N26990, N26989, N26988, N26987, N26986, N26985, N26984, N26983, N26982, N26981, N26980, N26979, N26978, N26977, N26976, N26975, N26974, N26973, N26972, N26971, N26970, N26969, N26968, N26967, N26966, N26965, N26964, N26963, N26962, N26961, N26960, N26959, N26958, N26957, N26956, N26955, N26954, N26953, N26952, N26951, N26950, N26949, N26948, N26947, N26946, N26945, N26944, N26943, N26942, N26941, N26940, N26939, N26938, N26937, N26936, N26935, N26934, N26933, N26932, N26931, N26930, N26929, N26928, N26927, N26926, N26925, N26924, N26923, N26922, N26921, N26920, N26919, N26918, N26917, N26916, N26915, N26914, N26913, N26912, N26911, N26910, N26909, N26908, N26907, N26906, N26905, N26904, N26903, N26902, N26901, N26900, N26899, N26898, N26897, N26896, N26895, N26894, N26893, N26892, N26891, N26890, N26889, N26888, N26887, N26886, N26885, N26884, N26883, N26882, N26881, N26880, N26879, N26878, N26877, N26876, N26875, N26874, N26873, N26872, N26871, N26870, N26869, N26868, N26867, N26866, N26865, N26864, N26863, N26862, N26861, N26860, N26859, N26858, N26857, N26856, N26855, N26854, N26853, N26852, N26851, N26850, N26849, N26848, N26847, N26846, N26845, N26844, N26843, N26842, N26841, N26840, N26839, N26838, N26837, N26836, N26835, N26834, N26833, N26832, N26831, N26830, N26829, N26828, N26827, N26826, N26825, N26824, N26823, N26822, N26821, N26820, N26819, N26818, N26817, N26816, N26815, N26814, N26813, N26812, N26811, N26810, N26809, N26808, N26807, N26806, N26805, N26804, N26803, N26802, N26801, N26800, N26799, N26798, N26797, N26796, N26795, N26794, N26793, N26792, N26791, N26790, N26789, N26788, N26787, N26786, N26785, N26784, N26783, N26782, N26781, N26780, N26779, N26778, N26777, N26776, N26775, N26774, N26773, N26772, N26771, N26770, N26769, N26768, N26767, N26766, N26765, N26764, N26763, N26762, N26761, N26760, N26759, N26758, N26757, N26756, N26755, N26754, N26753, N26752, N26751, N26750, N26749, N26748, N26747, N26746, N26745, N26744, N26743, N26742, N26741, N26740, N26739, N26738, N26737, N26736, N26735, N26734, N26733, N26732, N26731, N26730, N26729, N26728, N26727, N26726, N26725, N26724, N26723, N26722, N26721, N26720, N26719, N26718, N26717, N26716, N26715, N26714, N26713, N26712, N26711, N26710, N26709, N26708, N26707, N26706 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N202)? { N24525, N24524, N24523, N24522, N24521, N24520, N24519, N24518, N24517, N24516, N24515, N24514, N24513, N24512, N24511, N24510, N24509, N24508, N24507, N24506, N24505, N24504, N24503, N24502, N24501, N24500, N24499, N24498, N24497, N24496, N24495, N24494, N24493, N24492, N24491, N24490, N24489, N24488, N24487, N24486, N24485, N24484, N24483, N24482, N24481, N24480, N24479, N24478, N24477, N24476, N24475, N24474, N24473, N24472, N24471, N24470, N24469, N24468, N24467, N24466, N24465, N24464, N24463, N24462, N24267, N24266, N24265, N24264, N24263, N24262, N24261, N24260, N24259, N24258, N24257, N24256, N24255, N24254, N24253, N24252, N24251, N24250, N24249, N24248, N24247, N24246, N24245, N24244, N24243, N24242, N24241, N24240, N24239, N24238, N24237, N24236, N24235, N24234, N24233, N24232, N24231, N24230, N24229, N24228, N24227, N24226, N24225, N24224, N24223, N24222, N24221, N24220, N24219, N24218, N24217, N24216, N24215, N24214, N24213, N24212, N24211, N24210, N24209, N24208, N24207, N24206, N24205, N24204, N24009, N24008, N24007, N24006, N24005, N24004, N24003, N24002, N24001, N24000, N23999, N23998, N23997, N23996, N23995, N23994, N23993, N23992, N23991, N23990, N23989, N23988, N23987, N23986, N23985, N23984, N23983, N23982, N23981, N23980, N23979, N23978, N23977, N23976, N23975, N23974, N23973, N23972, N23971, N23970, N23969, N23968, N23967, N23966, N23965, N23964, N23963, N23962, N23961, N23960, N23959, N23958, N23957, N23956, N23955, N23954, N23953, N23952, N23951, N23950, N23949, N23948, N23947, N23946, N23751, N23750, N23749, N23748, N23747, N23746, N23745, N23744, N23743, N23742, N23741, N23740, N23739, N23738, N23737, N23736, N23735, N23734, N23733, N23732, N23731, N23730, N23729, N23728, N23727, N23726, N23725, N23724, N23723, N23722, N23721, N23720, N23719, N23718, N23717, N23716, N23715, N23714, N23713, N23712, N23711, N23710, N23709, N23708, N23707, N23706, N23705, N23704, N23703, N23702, N23701, N23700, N23699, N23698, N23697, N23696, N23695, N23694, N23693, N23692, N23691, N23690, N23689, N23688, N23493, N23492, N23491, N23490, N23489, N23488, N23487, N23486, N23485, N23484, N23483, N23482, N23481, N23480, N23479, N23478, N23477, N23476, N23475, N23474, N23473, N23472, N23471, N23470, N23469, N23468, N23467, N23466, N23465, N23464, N23463, N23462, N23461, N23460, N23459, N23458, N23457, N23456, N23455, N23454, N23453, N23452, N23451, N23450, N23449, N23448, N23447, N23446, N23445, N23444, N23443, N23442, N23441, N23440, N23439, N23438, N23437, N23436, N23435, N23434, N23433, N23432, N23431, N23430, N23235, N23234, N23233, N23232, N23231, N23230, N23229, N23228, N23227, N23226, N23225, N23224, N23223, N23222, N23221, N23220, N23219, N23218, N23217, N23216, N23215, N23214, N23213, N23212, N23211, N23210, N23209, N23208, N23207, N23206, N23205, N23204, N23203, N23202, N23201, N23200, N23199, N23198, N23197, N23196, N23195, N23194, N23193, N23192, N23191, N23190, N23189, N23188, N23187, N23186, N23185, N23184, N23183, N23182, N23181, N23180, N23179, N23178, N23177, N23176, N23175, N23174, N23173, N23172, N22977, N22976, N22975, N22974, N22973, N22972, N22971, N22970, N22969, N22968, N22967, N22966, N22965, N22964, N22963, N22962, N22961, N22960, N22959, N22958, N22957, N22956, N22955, N22954, N22953, N22952, N22951, N22950, N22949, N22948, N22947, N22946, N22945, N22944, N22943, N22942, N22941, N22940, N22939, N22938, N22937, N22936, N22935, N22934, N22933, N22932, N22931, N22930, N22929, N22928, N22927, N22926, N22925, N22924, N22923, N22922, N22921, N22920, N22919, N22918, N22917, N22916, N22915, N22914, N22719, N22718, N22717, N22716, N22715, N22714, N22713, N22712, N22711, N22710, N22709, N22708, N22707, N22706, N22705, N22704, N22703, N22702, N22701, N22700, N22699, N22698, N22697, N22696, N22695, N22694, N22693, N22692, N22691, N22690, N22689, N22688, N22687, N22686, N22685, N22684, N22683, N22682, N22681, N22680, N22679, N22678, N22677, N22676, N22675, N22674, N22673, N22672, N22671, N22670, N22669, N22668, N22667, N22666, N22665, N22664, N22663, N22662, N22661, N22660, N22659, N22658, N22657, N22656 } : 1'b0;
  assign N201 = N26704;
  assign N202 = N26705;
  assign { N28761, N28760, N28759, N28758, N28757, N28756, N28755, N28754, N28753, N28752, N28751, N28750, N28749, N28748, N28747, N28746, N28745, N28744, N28743, N28742, N28741, N28740, N28739, N28738, N28737, N28736, N28735, N28734, N28733, N28732, N28731, N28730, N28729, N28728, N28727, N28726, N28725, N28724, N28723, N28722, N28721, N28720, N28719, N28718, N28717, N28716, N28715, N28714, N28713, N28712, N28711, N28710, N28709, N28708, N28707, N28706, N28705, N28704, N28703, N28702, N28701, N28700, N28699, N28698, N28697, N28696, N28695, N28694, N28693, N28692, N28691, N28690, N28689, N28688, N28687, N28686, N28685, N28684, N28683, N28682, N28681, N28680, N28679, N28678, N28677, N28676, N28675, N28674, N28673, N28672, N28671, N28670, N28669, N28668, N28667, N28666, N28665, N28664, N28663, N28662, N28661, N28660, N28659, N28658, N28657, N28656, N28655, N28654, N28653, N28652, N28651, N28650, N28649, N28648, N28647, N28646, N28645, N28644, N28643, N28642, N28641, N28640, N28639, N28638, N28637, N28636, N28635, N28634, N28633, N28632, N28631, N28630, N28629, N28628, N28627, N28626, N28625, N28624, N28623, N28622, N28621, N28620, N28619, N28618, N28617, N28616, N28615, N28614, N28613, N28612, N28611, N28610, N28609, N28608, N28607, N28606, N28605, N28604, N28603, N28602, N28601, N28600, N28599, N28598, N28597, N28596, N28595, N28594, N28593, N28592, N28591, N28590, N28589, N28588, N28587, N28586, N28585, N28584, N28583, N28582, N28581, N28580, N28579, N28578, N28577, N28576, N28575, N28574, N28573, N28572, N28571, N28570, N28569, N28568, N28567, N28566, N28565, N28564, N28563, N28562, N28561, N28560, N28559, N28558, N28557, N28556, N28555, N28554, N28553, N28552, N28551, N28550, N28549, N28548, N28547, N28546, N28545, N28544, N28543, N28542, N28541, N28540, N28539, N28538, N28537, N28536, N28535, N28534, N28533, N28532, N28531, N28530, N28529, N28528, N28527, N28526, N28525, N28524, N28523, N28522, N28521, N28520, N28519, N28518, N28517, N28516, N28515, N28514, N28513, N28512, N28511, N28510, N28509, N28508, N28507, N28506, N28505, N28504, N28503, N28502, N28501, N28500, N28499, N28498, N28497, N28496, N28495, N28494, N28493, N28492, N28491, N28490, N28489, N28488, N28487, N28486, N28485, N28484, N28483, N28482, N28481, N28480, N28479, N28478, N28477, N28476, N28475, N28474, N28473, N28472, N28471, N28470, N28469, N28468, N28467, N28466, N28465, N28464, N28463, N28462, N28461, N28460, N28459, N28458, N28457, N28456, N28455, N28454, N28453, N28452, N28451, N28450, N28449, N28448, N28447, N28446, N28445, N28444, N28443, N28442, N28441, N28440, N28439, N28438, N28437, N28436, N28435, N28434, N28433, N28432, N28431, N28430, N28429, N28428, N28427, N28426, N28425, N28424, N28423, N28422, N28421, N28420, N28419, N28418, N28417, N28416, N28415, N28414, N28413, N28412, N28411, N28410, N28409, N28408, N28407, N28406, N28405, N28404, N28403, N28402, N28401, N28400, N28399, N28398, N28397, N28396, N28395, N28394, N28393, N28392, N28391, N28390, N28389, N28388, N28387, N28386, N28385, N28384, N28383, N28382, N28381, N28380, N28379, N28378, N28377, N28376, N28375, N28374, N28373, N28372, N28371, N28370, N28369, N28368, N28367, N28366, N28365, N28364, N28363, N28362, N28361, N28360, N28359, N28358, N28357, N28356, N28355, N28354, N28353, N28352, N28351, N28350, N28349, N28348, N28347, N28346, N28345, N28344, N28343, N28342, N28341, N28340, N28339, N28338, N28337, N28336, N28335, N28334, N28333, N28332, N28331, N28330, N28329, N28328, N28327, N28326, N28325, N28324, N28323, N28322, N28321, N28320, N28319, N28318, N28317, N28316, N28315, N28314, N28313, N28312, N28311, N28310, N28309, N28308, N28307, N28306, N28305, N28304, N28303, N28302, N28301, N28300, N28299, N28298, N28297, N28296, N28295, N28294, N28293, N28292, N28291, N28290, N28289, N28288, N28287, N28286, N28285, N28284, N28283, N28282, N28281, N28280, N28279, N28278, N28277, N28276, N28275, N28274, N28273, N28272, N28271, N28270, N28269, N28268, N28267, N28266, N28265, N28264, N28263, N28262, N28261, N28260, N28259, N28258, N28257, N28256, N28255, N28254, N28253, N28252, N28251, N28250, N28249, N28248, N28247, N28246, N28245, N28244, N28243, N28242, N28241, N28240, N28239, N28238, N28237, N28236, N28235, N28234, N28233, N28232, N28231, N28230, N28229, N28228, N28227, N28226, N28225, N28224, N28223, N28222, N28221, N28220, N28219, N28218, N28217, N28216, N28215, N28214, N28213, N28212, N28211, N28210, N28209, N28208, N28207, N28206, N28205, N28204, N28203, N28202, N28201, N28200, N28199, N28198, N28197, N28196, N28195, N28194, N28193, N28192, N28191, N28190, N28189, N28188, N28187, N28186, N28185, N28184, N28183, N28182, N28181, N28180, N28179, N28178, N28177, N28176, N28175, N28174, N28173, N28172, N28171, N28170, N28169, N28168, N28167, N28166, N28165, N28164, N28163, N28162, N28161, N28160, N28159, N28158, N28157, N28156, N28155, N28154, N28153, N28152, N28151, N28150, N28149, N28148, N28147, N28146, N28145, N28144, N28143, N28142, N28141, N28140, N28139, N28138, N28137, N28136, N28135, N28134, N28133, N28132, N28131, N28130, N28129, N28128, N28127, N28126, N28125, N28124, N28123, N28122, N28121, N28120, N28119, N28118, N28117, N28116, N28115, N28114, N28113, N28112, N28111, N28110, N28109, N28108, N28107, N28106, N28105, N28104, N28103, N28102, N28101, N28100, N28099, N28098, N28097, N28096, N28095, N28094, N28093, N28092, N28091, N28090, N28089, N28088, N28087, N28086, N28085, N28084, N28083, N28082, N28081, N28080, N28079, N28078, N28077, N28076, N28075, N28074, N28073, N28072, N28071, N28070, N28069, N28068, N28067, N28066, N28065, N28064, N28063, N28062, N28061, N28060, N28059, N28058, N28057, N28056, N28055, N28054, N28053, N28052, N28051, N28050, N28049, N28048, N28047, N28046, N28045, N28044, N28043, N28042, N28041, N28040, N28039, N28038, N28037, N28036, N28035, N28034, N28033, N28032, N28031, N28030, N28029, N28028, N28027, N28026, N28025, N28024, N28023, N28022, N28021, N28020, N28019, N28018, N28017, N28016, N28015, N28014, N28013, N28012, N28011, N28010, N28009, N28008, N28007, N28006, N28005, N28004, N28003, N28002, N28001, N28000, N27999, N27998, N27997, N27996, N27995, N27994, N27993, N27992, N27991, N27990, N27989, N27988, N27987, N27986, N27985, N27984, N27983, N27982, N27981, N27980, N27979, N27978, N27977, N27976, N27975, N27974, N27973, N27972, N27971, N27970, N27969, N27968, N27967, N27966, N27965, N27964, N27963, N27962, N27961, N27960, N27959, N27958, N27957, N27956, N27955, N27954, N27953, N27952, N27951, N27950, N27949, N27948, N27947, N27946, N27945, N27944, N27943, N27942, N27941, N27940, N27939, N27938, N27937, N27936, N27935, N27934, N27933, N27932, N27931, N27930, N27929, N27928, N27927, N27926, N27925, N27924, N27923, N27922, N27921, N27920, N27919, N27918, N27917, N27916, N27915, N27914, N27913, N27912, N27911, N27910, N27909, N27908, N27907, N27906, N27905, N27904, N27903, N27902, N27901, N27900, N27899, N27898, N27897, N27896, N27895, N27894, N27893, N27892, N27891, N27890, N27889, N27888, N27887, N27886, N27885, N27884, N27883, N27882, N27881, N27880, N27879, N27878, N27877, N27876, N27875, N27874, N27873, N27872, N27871, N27870, N27869, N27868, N27867, N27866, N27865, N27864, N27863, N27862, N27861, N27860, N27859, N27858, N27857, N27856, N27855, N27854, N27853, N27852, N27851, N27850, N27849, N27848, N27847, N27846, N27845, N27844, N27843, N27842, N27841, N27840, N27839, N27838, N27837, N27836, N27835, N27834, N27833, N27832, N27831, N27830, N27829, N27828, N27827, N27826, N27825, N27824, N27823, N27822, N27821, N27820, N27819, N27818, N27817, N27816, N27815, N27814, N27813, N27812, N27811, N27810, N27809, N27808, N27807, N27806, N27805, N27804, N27803, N27802, N27801, N27800, N27799, N27798, N27797, N27796, N27795, N27794, N27793, N27792, N27791, N27790, N27789, N27788, N27787, N27786, N27785, N27784, N27783, N27782, N27781, N27780, N27779, N27778, N27777, N27776, N27775, N27774, N27773, N27772, N27771, N27770, N27769, N27768, N27767, N27766, N27765, N27764, N27763, N27762, N27761, N27760, N27759, N27758, N27757, N27756, N27755, N27754, N27753, N27752, N27751, N27750, N27749, N27748, N27747, N27746, N27745, N27744, N27743, N27742, N27741, N27740, N27739, N27738, N27737, N27736, N27735, N27734, N27733, N27732, N27731, N27730 } = (N203)? { N26693, N26692, N26691, N26690, N26689, N26688, N26687, N26686, N26685, N26684, N26683, N26682, N26681, N26680, N26679, N26678, N26677, N26676, N26675, N26674, N26673, N26672, N26671, N26670, N26669, N26668, N26667, N26666, N26665, N26664, N26663, N26662, N26661, N26660, N26659, N26658, N26657, N26656, N26655, N26654, N26653, N26652, N26651, N26650, N26649, N26648, N26647, N26646, N26645, N26644, N26643, N26642, N26641, N26640, N26639, N26638, N26637, N26636, N26635, N26634, N26633, N26632, N26631, N26630, N26629, N26628, N26627, N26626, N26625, N26624, N26623, N26622, N26621, N26620, N26619, N26618, N26617, N26616, N26615, N26614, N26613, N26612, N26611, N26610, N26609, N26608, N26607, N26606, N26605, N26604, N26603, N26602, N26601, N26600, N26599, N26598, N26597, N26596, N26595, N26594, N26593, N26592, N26591, N26590, N26589, N26588, N26587, N26586, N26585, N26584, N26583, N26582, N26581, N26580, N26579, N26578, N26577, N26576, N26575, N26574, N26573, N26572, N26571, N26570, N26569, N26568, N26567, N26566, N26565, N26564, N26563, N26562, N26561, N26560, N26559, N26558, N26557, N26556, N26555, N26554, N26553, N26552, N26551, N26550, N26549, N26548, N26547, N26546, N26545, N26544, N26543, N26542, N26541, N26540, N26539, N26538, N26537, N26536, N26535, N26534, N26533, N26532, N26531, N26530, N26529, N26528, N26527, N26526, N26525, N26524, N26523, N26522, N26521, N26520, N26519, N26518, N26517, N26516, N26515, N26514, N26513, N26512, N26511, N26510, N26509, N26508, N26507, N26506, N26505, N26504, N26503, N26502, N26501, N26500, N26499, N26498, N26497, N26496, N26495, N26494, N26493, N26492, N26491, N26490, N26489, N26488, N26487, N26486, N26485, N26484, N26483, N26482, N26481, N26480, N26479, N26478, N26477, N26476, N26475, N26474, N26473, N26472, N26471, N26470, N26469, N26468, N26467, N26466, N26465, N26464, N26463, N26462, N26461, N26460, N26459, N26458, N26457, N26456, N26455, N26454, N26453, N26452, N26451, N26450, N26449, N26448, N26447, N26446, N26445, N26444, N26443, N26442, N26441, N26440, N26439, N26438, N26437, N26436, N26435, N26434, N26433, N26432, N26431, N26430, N26429, N26428, N26427, N26426, N26425, N26424, N26423, N26422, N26421, N26420, N26419, N26418, N26417, N26416, N26415, N26414, N26413, N26412, N26411, N26410, N26409, N26408, N26407, N26406, N26405, N26404, N26403, N26402, N26401, N26400, N26399, N26398, N26397, N26396, N26395, N26394, N26393, N26392, N26391, N26390, N26389, N26388, N26387, N26386, N26385, N26384, N26383, N26382, N26381, N26380, N26379, N26378, N26377, N26376, N26375, N26374, N26373, N26372, N26371, N26370, N26369, N26368, N26367, N26366, N26365, N26364, N26363, N26362, N26361, N26360, N26359, N26358, N26357, N26356, N26355, N26354, N26353, N26352, N26351, N26350, N26349, N26348, N26347, N26346, N26345, N26344, N26343, N26342, N26341, N26340, N26339, N26338, N26337, N26336, N26335, N26334, N26333, N26332, N26331, N26330, N26329, N26328, N26327, N26326, N26325, N26324, N26323, N26322, N26321, N26320, N26319, N26318, N26317, N26316, N26315, N26314, N26313, N26312, N26311, N26310, N26309, N26308, N26307, N26306, N26305, N26304, N26303, N26302, N26301, N26300, N26299, N26298, N26297, N26296, N26295, N26294, N26293, N26292, N26291, N26290, N26289, N26288, N26287, N26286, N26285, N26284, N26283, N26282, N26281, N26280, N26279, N26278, N26277, N26276, N26275, N26274, N26273, N26272, N26271, N26270, N26269, N26268, N26267, N26266, N26265, N26264, N26263, N26262, N26261, N26260, N26259, N26258, N26257, N26256, N26255, N26254, N26253, N26252, N26251, N26250, N26249, N26248, N26247, N26246, N26245, N26244, N26243, N26242, N26241, N26240, N26239, N26238, N26237, N26236, N26235, N26234, N26233, N26232, N26231, N26230, N26229, N26228, N26227, N26226, N26225, N26224, N26223, N26222, N26221, N26220, N26219, N26218, N26217, N26216, N26215, N26214, N26213, N26212, N26211, N26210, N26209, N26208, N26207, N26206, N26205, N26204, N26203, N26202, N26201, N26200, N26199, N26198, N26197, N26196, N26195, N26194, N26193, N26192, N26191, N26190, N26189, N26188, N26187, N26186, N26185, N26184, N26183, N26182, N26181, N26180, N26179, N26178, N26177, N26176, N26175, N26174, N26173, N26172, N26171, N26170, N26169, N26168, N26167, N26166, N26165, N26164, N26163, N26162, N26161, N26160, N26159, N26158, N26157, N26156, N26155, N26154, N26153, N26152, N26151, N26150, N26149, N26148, N26147, N26146, N26145, N26144, N26143, N26142, N26141, N26140, N26139, N26138, N26137, N26136, N26135, N26134, N26133, N26132, N26131, N26130, N26129, N26128, N26127, N26126, N26125, N26124, N26123, N26122, N26121, N26120, N26119, N26118, N26117, N26116, N26115, N26114, N26113, N26112, N26111, N26110, N26109, N26108, N26107, N26106, N26105, N26104, N26103, N26102, N26101, N26100, N26099, N26098, N26097, N26096, N26095, N26094, N26093, N26092, N26091, N26090, N26089, N26088, N26087, N26086, N26085, N26084, N26083, N26082, N26081, N26080, N26079, N26078, N26077, N26076, N26075, N26074, N26073, N26072, N26071, N26070, N26069, N26068, N26067, N26066, N26065, N26064, N26063, N26062, N26061, N26060, N26059, N26058, N26057, N26056, N26055, N26054, N26053, N26052, N26051, N26050, N26049, N26048, N26047, N26046, N26045, N26044, N26043, N26042, N26041, N26040, N26039, N26038, N26037, N26036, N26035, N26034, N26033, N26032, N26031, N26030, N26029, N26028, N26027, N26026, N26025, N26024, N26023, N26022, N26021, N26020, N26019, N26018, N26017, N26016, N26015, N26014, N26013, N26012, N26011, N26010, N26009, N26008, N26007, N26006, N26005, N26004, N26003, N26002, N26001, N26000, N25999, N25998, N25997, N25996, N25995, N25994, N25993, N25992, N25991, N25990, N25989, N25988, N25987, N25986, N25985, N25984, N25983, N25982, N25981, N25980, N25979, N25978, N25977, N25976, N25975, N25974, N25973, N25972, N25971, N25970, N25969, N25968, N25967, N25966, N25965, N25964, N25963, N25962, N25961, N25960, N25959, N25958, N25957, N25956, N25955, N25954, N25953, N25952, N25951, N25950, N25949, N25948, N25947, N25946, N25945, N25944, N25943, N25942, N25941, N25940, N25939, N25938, N25937, N25936, N25935, N25934, N25933, N25932, N25931, N25930, N25929, N25928, N25927, N25926, N25925, N25924, N25923, N25922, N25921, N25920, N25919, N25918, N25917, N25916, N25915, N25914, N25913, N25912, N25911, N25910, N25909, N25908, N25907, N25906, N25905, N25904, N25903, N25902, N25901, N25900, N25899, N25898, N25897, N25896, N25895, N25894, N25893, N25892, N25891, N25890, N25889, N25888, N25887, N25886, N25885, N25884, N25883, N25882, N25881, N25880, N25879, N25878, N25877, N25876, N25875, N25874, N25873, N25872, N25871, N25870, N25869, N25868, N25867, N25866, N25865, N25864, N25863, N25862, N25861, N25860, N25859, N25858, N25857, N25856, N25855, N25854, N25853, N25852, N25851, N25850, N25849, N25848, N25847, N25846, N25845, N25844, N25843, N25842, N25841, N25840, N25839, N25838, N25837, N25836, N25835, N25834, N25833, N25832, N25831, N25830, N25829, N25828, N25827, N25826, N25825, N25824, N25823, N25822, N25821, N25820, N25819, N25818, N25817, N25816, N25815, N25814, N25813, N25812, N25811, N25810, N25809, N25808, N25807, N25806, N25805, N25804, N25803, N25802, N25801, N25800, N25799, N25798, N25797, N25796, N25795, N25794, N25793, N25792, N25791, N25790, N25789, N25788, N25787, N25786, N25785, N25784, N25783, N25782, N25781, N25780, N25779, N25778, N25777, N25776, N25775, N25774, N25773, N25772, N25771, N25770, N25769, N25768, N25767, N25766, N25765, N25764, N25763, N25762, N25761, N25760, N25759, N25758, N25757, N25756, N25755, N25754, N25753, N25752, N25751, N25750, N25749, N25748, N25747, N25746, N25745, N25744, N25743, N25742, N25741, N25740, N25739, N25738, N25737, N25736, N25735, N25734, N25733, N25732, N25731, N25730, N25729, N25728, N25727, N25726, N25725, N25724, N25723, N25722, N25721, N25720, N25719, N25718, N25717, N25716, N25715, N25714, N25713, N25712, N25711, N25710, N25709, N25708, N25707, N25706, N25705, N25704, N25703, N25702, N25701, N25700, N25699, N25698, N25697, N25696, N25695, N25694, N25693, N25692, N25691, N25690, N25689, N25688, N25687, N25686, N25685, N25684, N25683, N25682, N25681, N25680, N25679, N25678, N25677, N25676, N25675, N25674, N25673, N25672, N25671, N25670, N25669, N25668, N25667, N25666, N25665, N25664, N25663, N25662 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25661)? { N27729, N27728, N27727, N27726, N27725, N27724, N27723, N27722, N27721, N27720, N27719, N27718, N27717, N27716, N27715, N27714, N27713, N27712, N27711, N27710, N27709, N27708, N27707, N27706, N27705, N27704, N27703, N27702, N27701, N27700, N27699, N27698, N27697, N27696, N27695, N27694, N27693, N27692, N27691, N27690, N27689, N27688, N27687, N27686, N27685, N27684, N27683, N27682, N27681, N27680, N27679, N27678, N27677, N27676, N27675, N27674, N27673, N27672, N27671, N27670, N27669, N27668, N27667, N27666, N24461, N24460, N24459, N24458, N24457, N24456, N24455, N24454, N24453, N24452, N24451, N24450, N24449, N24448, N24447, N24446, N24445, N24444, N24443, N24442, N24441, N24440, N24439, N24438, N24437, N24436, N24435, N24434, N24433, N24432, N24431, N24430, N24429, N24428, N24427, N24426, N24425, N24424, N24423, N24422, N24421, N24420, N24419, N24418, N24417, N24416, N24415, N24414, N24413, N24412, N24411, N24410, N24409, N24408, N24407, N24406, N24405, N24404, N24403, N24402, N24401, N24400, N24399, N24398, N24397, N27665, N27664, N27663, N27662, N27661, N27660, N27659, N27658, N27657, N27656, N27655, N27654, N27653, N27652, N27651, N27650, N27649, N27648, N27647, N27646, N27645, N27644, N27643, N27642, N27641, N27640, N27639, N27638, N27637, N27636, N27635, N27634, N27633, N27632, N27631, N27630, N27629, N27628, N27627, N27626, N27625, N27624, N27623, N27622, N27621, N27620, N27619, N27618, N27617, N27616, N27615, N27614, N27613, N27612, N27611, N27610, N27609, N27608, N27607, N27606, N27605, N27604, N27603, N27602, N24203, N24202, N24201, N24200, N24199, N24198, N24197, N24196, N24195, N24194, N24193, N24192, N24191, N24190, N24189, N24188, N24187, N24186, N24185, N24184, N24183, N24182, N24181, N24180, N24179, N24178, N24177, N24176, N24175, N24174, N24173, N24172, N24171, N24170, N24169, N24168, N24167, N24166, N24165, N24164, N24163, N24162, N24161, N24160, N24159, N24158, N24157, N24156, N24155, N24154, N24153, N24152, N24151, N24150, N24149, N24148, N24147, N24146, N24145, N24144, N24143, N24142, N24141, N24140, N24139, N27601, N27600, N27599, N27598, N27597, N27596, N27595, N27594, N27593, N27592, N27591, N27590, N27589, N27588, N27587, N27586, N27585, N27584, N27583, N27582, N27581, N27580, N27579, N27578, N27577, N27576, N27575, N27574, N27573, N27572, N27571, N27570, N27569, N27568, N27567, N27566, N27565, N27564, N27563, N27562, N27561, N27560, N27559, N27558, N27557, N27556, N27555, N27554, N27553, N27552, N27551, N27550, N27549, N27548, N27547, N27546, N27545, N27544, N27543, N27542, N27541, N27540, N27539, N27538, N23945, N23944, N23943, N23942, N23941, N23940, N23939, N23938, N23937, N23936, N23935, N23934, N23933, N23932, N23931, N23930, N23929, N23928, N23927, N23926, N23925, N23924, N23923, N23922, N23921, N23920, N23919, N23918, N23917, N23916, N23915, N23914, N23913, N23912, N23911, N23910, N23909, N23908, N23907, N23906, N23905, N23904, N23903, N23902, N23901, N23900, N23899, N23898, N23897, N23896, N23895, N23894, N23893, N23892, N23891, N23890, N23889, N23888, N23887, N23886, N23885, N23884, N23883, N23882, N23881, N27537, N27536, N27535, N27534, N27533, N27532, N27531, N27530, N27529, N27528, N27527, N27526, N27525, N27524, N27523, N27522, N27521, N27520, N27519, N27518, N27517, N27516, N27515, N27514, N27513, N27512, N27511, N27510, N27509, N27508, N27507, N27506, N27505, N27504, N27503, N27502, N27501, N27500, N27499, N27498, N27497, N27496, N27495, N27494, N27493, N27492, N27491, N27490, N27489, N27488, N27487, N27486, N27485, N27484, N27483, N27482, N27481, N27480, N27479, N27478, N27477, N27476, N27475, N27474, N23687, N23686, N23685, N23684, N23683, N23682, N23681, N23680, N23679, N23678, N23677, N23676, N23675, N23674, N23673, N23672, N23671, N23670, N23669, N23668, N23667, N23666, N23665, N23664, N23663, N23662, N23661, N23660, N23659, N23658, N23657, N23656, N23655, N23654, N23653, N23652, N23651, N23650, N23649, N23648, N23647, N23646, N23645, N23644, N23643, N23642, N23641, N23640, N23639, N23638, N23637, N23636, N23635, N23634, N23633, N23632, N23631, N23630, N23629, N23628, N23627, N23626, N23625, N23624, N23623, N27473, N27472, N27471, N27470, N27469, N27468, N27467, N27466, N27465, N27464, N27463, N27462, N27461, N27460, N27459, N27458, N27457, N27456, N27455, N27454, N27453, N27452, N27451, N27450, N27449, N27448, N27447, N27446, N27445, N27444, N27443, N27442, N27441, N27440, N27439, N27438, N27437, N27436, N27435, N27434, N27433, N27432, N27431, N27430, N27429, N27428, N27427, N27426, N27425, N27424, N27423, N27422, N27421, N27420, N27419, N27418, N27417, N27416, N27415, N27414, N27413, N27412, N27411, N27410, N23429, N23428, N23427, N23426, N23425, N23424, N23423, N23422, N23421, N23420, N23419, N23418, N23417, N23416, N23415, N23414, N23413, N23412, N23411, N23410, N23409, N23408, N23407, N23406, N23405, N23404, N23403, N23402, N23401, N23400, N23399, N23398, N23397, N23396, N23395, N23394, N23393, N23392, N23391, N23390, N23389, N23388, N23387, N23386, N23385, N23384, N23383, N23382, N23381, N23380, N23379, N23378, N23377, N23376, N23375, N23374, N23373, N23372, N23371, N23370, N23369, N23368, N23367, N23366, N23365, N27409, N27408, N27407, N27406, N27405, N27404, N27403, N27402, N27401, N27400, N27399, N27398, N27397, N27396, N27395, N27394, N27393, N27392, N27391, N27390, N27389, N27388, N27387, N27386, N27385, N27384, N27383, N27382, N27381, N27380, N27379, N27378, N27377, N27376, N27375, N27374, N27373, N27372, N27371, N27370, N27369, N27368, N27367, N27366, N27365, N27364, N27363, N27362, N27361, N27360, N27359, N27358, N27357, N27356, N27355, N27354, N27353, N27352, N27351, N27350, N27349, N27348, N27347, N27346, N23171, N23170, N23169, N23168, N23167, N23166, N23165, N23164, N23163, N23162, N23161, N23160, N23159, N23158, N23157, N23156, N23155, N23154, N23153, N23152, N23151, N23150, N23149, N23148, N23147, N23146, N23145, N23144, N23143, N23142, N23141, N23140, N23139, N23138, N23137, N23136, N23135, N23134, N23133, N23132, N23131, N23130, N23129, N23128, N23127, N23126, N23125, N23124, N23123, N23122, N23121, N23120, N23119, N23118, N23117, N23116, N23115, N23114, N23113, N23112, N23111, N23110, N23109, N23108, N23107, N27345, N27344, N27343, N27342, N27341, N27340, N27339, N27338, N27337, N27336, N27335, N27334, N27333, N27332, N27331, N27330, N27329, N27328, N27327, N27326, N27325, N27324, N27323, N27322, N27321, N27320, N27319, N27318, N27317, N27316, N27315, N27314, N27313, N27312, N27311, N27310, N27309, N27308, N27307, N27306, N27305, N27304, N27303, N27302, N27301, N27300, N27299, N27298, N27297, N27296, N27295, N27294, N27293, N27292, N27291, N27290, N27289, N27288, N27287, N27286, N27285, N27284, N27283, N27282, N22913, N22912, N22911, N22910, N22909, N22908, N22907, N22906, N22905, N22904, N22903, N22902, N22901, N22900, N22899, N22898, N22897, N22896, N22895, N22894, N22893, N22892, N22891, N22890, N22889, N22888, N22887, N22886, N22885, N22884, N22883, N22882, N22881, N22880, N22879, N22878, N22877, N22876, N22875, N22874, N22873, N22872, N22871, N22870, N22869, N22868, N22867, N22866, N22865, N22864, N22863, N22862, N22861, N22860, N22859, N22858, N22857, N22856, N22855, N22854, N22853, N22852, N22851, N22850, N22849, N27281, N27280, N27279, N27278, N27277, N27276, N27275, N27274, N27273, N27272, N27271, N27270, N27269, N27268, N27267, N27266, N27265, N27264, N27263, N27262, N27261, N27260, N27259, N27258, N27257, N27256, N27255, N27254, N27253, N27252, N27251, N27250, N27249, N27248, N27247, N27246, N27245, N27244, N27243, N27242, N27241, N27240, N27239, N27238, N27237, N27236, N27235, N27234, N27233, N27232, N27231, N27230, N27229, N27228, N27227, N27226, N27225, N27224, N27223, N27222, N27221, N27220, N27219, N27218, N22655, N22654, N22653, N22652, N22651, N22650, N22649, N22648, N22647, N22646, N22645, N22644, N22643, N22642, N22641, N22640, N22639, N22638, N22637, N22636, N22635, N22634, N22633, N22632, N22631, N22630, N22629, N22628, N22627, N22626, N22625, N22624, N22623, N22622, N22621, N22620, N22619, N22618, N22617, N22616, N22615, N22614, N22613, N22612, N22611, N22610, N22609, N22608, N22607, N22606, N22605, N22604, N22603, N22602, N22601, N22600, N22599, N22598, N22597, N22596, N22595, N22594, N22593, N22592, N22591 } : 1'b0;
  assign N203 = ex_i[387];
  assign { mem_n[2806:2743], N28777, mem_n[2738:2611], N28776, mem_n[2608:2545], mem_n[2443:2380], N28775, mem_n[2375:2248], N28774, mem_n[2245:2182], mem_n[2080:2017], N28773, mem_n[2012:1885], N28772, mem_n[1882:1819], mem_n[1717:1654], N28771, mem_n[1649:1522], N28770, mem_n[1519:1456], mem_n[1354:1291], N28769, mem_n[1286:1159], N28768, mem_n[1156:1093], mem_n[991:928], N28767, mem_n[923:796], N28766, mem_n[793:730], mem_n[628:565], N28765, mem_n[560:433], N28764, mem_n[430:367], mem_n[265:202], N28763, mem_n[197:70], N28762, mem_n[67:4] } = (N204)? { N25144, N25143, N25142, N25141, N25140, N25139, N25138, N25137, N25136, N25135, N25134, N25133, N25132, N25131, N25130, N25129, N25128, N25127, N25126, N25125, N25124, N25123, N25122, N25121, N25120, N25119, N25118, N25117, N25116, N25115, N25114, N25113, N25112, N25111, N25110, N25109, N25108, N25107, N25106, N25105, N25104, N25103, N25102, N25101, N25100, N25099, N25098, N25097, N25096, N25095, N25094, N25093, N25092, N25091, N25090, N25089, N25088, N25087, N25086, N25085, N25084, N25083, N25082, N25081, N24616, N28761, N28760, N28759, N28758, N28757, N28756, N28755, N28754, N28753, N28752, N28751, N28750, N28749, N28748, N28747, N28746, N28745, N28744, N28743, N28742, N28741, N28740, N28739, N28738, N28737, N28736, N28735, N28734, N28733, N28732, N28731, N28730, N28729, N28728, N28727, N28726, N28725, N28724, N28723, N28722, N28721, N28720, N28719, N28718, N28717, N28716, N28715, N28714, N28713, N28712, N28711, N28710, N28709, N28708, N28707, N28706, N28705, N28704, N28703, N28702, N28701, N28700, N28699, N28698, N28697, N28696, N28695, N28694, N28693, N28692, N28691, N28690, N28689, N28688, N28687, N28686, N28685, N28684, N28683, N28682, N28681, N28680, N28679, N28678, N28677, N28676, N28675, N28674, N28673, N28672, N28671, N28670, N28669, N28668, N28667, N28666, N28665, N28664, N28663, N28662, N28661, N28660, N28659, N28658, N28657, N28656, N28655, N28654, N28653, N28652, N28651, N28650, N28649, N28648, N28647, N28646, N28645, N28644, N28643, N28642, N28641, N28640, N28639, N28638, N28637, N28636, N28635, N28634, N28633, N25656, N25655, N25654, N25653, N25652, N25651, N25650, N25649, N25648, N25647, N25646, N25645, N25644, N25643, N25642, N25641, N25640, N25639, N25638, N25637, N25636, N25635, N25634, N25633, N25632, N25631, N25630, N25629, N25628, N25627, N25626, N25625, N25624, N25623, N25622, N25621, N25620, N25619, N25618, N25617, N25616, N25615, N25614, N25613, N25612, N25611, N25610, N25609, N25608, N25607, N25606, N25605, N25604, N25603, N25602, N25601, N25600, N25599, N25598, N25597, N25596, N25595, N25594, N25593, N25079, N25078, N25077, N25076, N25075, N25074, N25073, N25072, N25071, N25070, N25069, N25068, N25067, N25066, N25065, N25064, N25063, N25062, N25061, N25060, N25059, N25058, N25057, N25056, N25055, N25054, N25053, N25052, N25051, N25050, N25049, N25048, N25047, N25046, N25045, N25044, N25043, N25042, N25041, N25040, N25039, N25038, N25037, N25036, N25035, N25034, N25033, N25032, N25031, N25030, N25029, N25028, N25027, N25026, N25025, N25024, N25023, N25022, N25021, N25020, N25019, N25018, N25017, N25016, N24615, N28632, N28631, N28630, N28629, N28628, N28627, N28626, N28625, N28624, N28623, N28622, N28621, N28620, N28619, N28618, N28617, N28616, N28615, N28614, N28613, N28612, N28611, N28610, N28609, N28608, N28607, N28606, N28605, N28604, N28603, N28602, N28601, N28600, N28599, N28598, N28597, N28596, N28595, N28594, N28593, N28592, N28591, N28590, N28589, N28588, N28587, N28586, N28585, N28584, N28583, N28582, N28581, N28580, N28579, N28578, N28577, N28576, N28575, N28574, N28573, N28572, N28571, N28570, N28569, N28568, N28567, N28566, N28565, N28564, N28563, N28562, N28561, N28560, N28559, N28558, N28557, N28556, N28555, N28554, N28553, N28552, N28551, N28550, N28549, N28548, N28547, N28546, N28545, N28544, N28543, N28542, N28541, N28540, N28539, N28538, N28537, N28536, N28535, N28534, N28533, N28532, N28531, N28530, N28529, N28528, N28527, N28526, N28525, N28524, N28523, N28522, N28521, N28520, N28519, N28518, N28517, N28516, N28515, N28514, N28513, N28512, N28511, N28510, N28509, N28508, N28507, N28506, N28505, N28504, N25592, N25591, N25590, N25589, N25588, N25587, N25586, N25585, N25584, N25583, N25582, N25581, N25580, N25579, N25578, N25577, N25576, N25575, N25574, N25573, N25572, N25571, N25570, N25569, N25568, N25567, N25566, N25565, N25564, N25563, N25562, N25561, N25560, N25559, N25558, N25557, N25556, N25555, N25554, N25553, N25552, N25551, N25550, N25549, N25548, N25547, N25546, N25545, N25544, N25543, N25542, N25541, N25540, N25539, N25538, N25537, N25536, N25535, N25534, N25533, N25532, N25531, N25530, N25529, N25014, N25013, N25012, N25011, N25010, N25009, N25008, N25007, N25006, N25005, N25004, N25003, N25002, N25001, N25000, N24999, N24998, N24997, N24996, N24995, N24994, N24993, N24992, N24991, N24990, N24989, N24988, N24987, N24986, N24985, N24984, N24983, N24982, N24981, N24980, N24979, N24978, N24977, N24976, N24975, N24974, N24973, N24972, N24971, N24970, N24969, N24968, N24967, N24966, N24965, N24964, N24963, N24962, N24961, N24960, N24959, N24958, N24957, N24956, N24955, N24954, N24953, N24952, N24951, N24614, N28503, N28502, N28501, N28500, N28499, N28498, N28497, N28496, N28495, N28494, N28493, N28492, N28491, N28490, N28489, N28488, N28487, N28486, N28485, N28484, N28483, N28482, N28481, N28480, N28479, N28478, N28477, N28476, N28475, N28474, N28473, N28472, N28471, N28470, N28469, N28468, N28467, N28466, N28465, N28464, N28463, N28462, N28461, N28460, N28459, N28458, N28457, N28456, N28455, N28454, N28453, N28452, N28451, N28450, N28449, N28448, N28447, N28446, N28445, N28444, N28443, N28442, N28441, N28440, N28439, N28438, N28437, N28436, N28435, N28434, N28433, N28432, N28431, N28430, N28429, N28428, N28427, N28426, N28425, N28424, N28423, N28422, N28421, N28420, N28419, N28418, N28417, N28416, N28415, N28414, N28413, N28412, N28411, N28410, N28409, N28408, N28407, N28406, N28405, N28404, N28403, N28402, N28401, N28400, N28399, N28398, N28397, N28396, N28395, N28394, N28393, N28392, N28391, N28390, N28389, N28388, N28387, N28386, N28385, N28384, N28383, N28382, N28381, N28380, N28379, N28378, N28377, N28376, N28375, N25528, N25527, N25526, N25525, N25524, N25523, N25522, N25521, N25520, N25519, N25518, N25517, N25516, N25515, N25514, N25513, N25512, N25511, N25510, N25509, N25508, N25507, N25506, N25505, N25504, N25503, N25502, N25501, N25500, N25499, N25498, N25497, N25496, N25495, N25494, N25493, N25492, N25491, N25490, N25489, N25488, N25487, N25486, N25485, N25484, N25483, N25482, N25481, N25480, N25479, N25478, N25477, N25476, N25475, N25474, N25473, N25472, N25471, N25470, N25469, N25468, N25467, N25466, N25465, N24949, N24948, N24947, N24946, N24945, N24944, N24943, N24942, N24941, N24940, N24939, N24938, N24937, N24936, N24935, N24934, N24933, N24932, N24931, N24930, N24929, N24928, N24927, N24926, N24925, N24924, N24923, N24922, N24921, N24920, N24919, N24918, N24917, N24916, N24915, N24914, N24913, N24912, N24911, N24910, N24909, N24908, N24907, N24906, N24905, N24904, N24903, N24902, N24901, N24900, N24899, N24898, N24897, N24896, N24895, N24894, N24893, N24892, N24891, N24890, N24889, N24888, N24887, N24886, N24613, N28374, N28373, N28372, N28371, N28370, N28369, N28368, N28367, N28366, N28365, N28364, N28363, N28362, N28361, N28360, N28359, N28358, N28357, N28356, N28355, N28354, N28353, N28352, N28351, N28350, N28349, N28348, N28347, N28346, N28345, N28344, N28343, N28342, N28341, N28340, N28339, N28338, N28337, N28336, N28335, N28334, N28333, N28332, N28331, N28330, N28329, N28328, N28327, N28326, N28325, N28324, N28323, N28322, N28321, N28320, N28319, N28318, N28317, N28316, N28315, N28314, N28313, N28312, N28311, N28310, N28309, N28308, N28307, N28306, N28305, N28304, N28303, N28302, N28301, N28300, N28299, N28298, N28297, N28296, N28295, N28294, N28293, N28292, N28291, N28290, N28289, N28288, N28287, N28286, N28285, N28284, N28283, N28282, N28281, N28280, N28279, N28278, N28277, N28276, N28275, N28274, N28273, N28272, N28271, N28270, N28269, N28268, N28267, N28266, N28265, N28264, N28263, N28262, N28261, N28260, N28259, N28258, N28257, N28256, N28255, N28254, N28253, N28252, N28251, N28250, N28249, N28248, N28247, N28246, N25464, N25463, N25462, N25461, N25460, N25459, N25458, N25457, N25456, N25455, N25454, N25453, N25452, N25451, N25450, N25449, N25448, N25447, N25446, N25445, N25444, N25443, N25442, N25441, N25440, N25439, N25438, N25437, N25436, N25435, N25434, N25433, N25432, N25431, N25430, N25429, N25428, N25427, N25426, N25425, N25424, N25423, N25422, N25421, N25420, N25419, N25418, N25417, N25416, N25415, N25414, N25413, N25412, N25411, N25410, N25409, N25408, N25407, N25406, N25405, N25404, N25403, N25402, N25401, N24884, N24883, N24882, N24881, N24880, N24879, N24878, N24877, N24876, N24875, N24874, N24873, N24872, N24871, N24870, N24869, N24868, N24867, N24866, N24865, N24864, N24863, N24862, N24861, N24860, N24859, N24858, N24857, N24856, N24855, N24854, N24853, N24852, N24851, N24850, N24849, N24848, N24847, N24846, N24845, N24844, N24843, N24842, N24841, N24840, N24839, N24838, N24837, N24836, N24835, N24834, N24833, N24832, N24831, N24830, N24829, N24828, N24827, N24826, N24825, N24824, N24823, N24822, N24821, N24612, N28245, N28244, N28243, N28242, N28241, N28240, N28239, N28238, N28237, N28236, N28235, N28234, N28233, N28232, N28231, N28230, N28229, N28228, N28227, N28226, N28225, N28224, N28223, N28222, N28221, N28220, N28219, N28218, N28217, N28216, N28215, N28214, N28213, N28212, N28211, N28210, N28209, N28208, N28207, N28206, N28205, N28204, N28203, N28202, N28201, N28200, N28199, N28198, N28197, N28196, N28195, N28194, N28193, N28192, N28191, N28190, N28189, N28188, N28187, N28186, N28185, N28184, N28183, N28182, N28181, N28180, N28179, N28178, N28177, N28176, N28175, N28174, N28173, N28172, N28171, N28170, N28169, N28168, N28167, N28166, N28165, N28164, N28163, N28162, N28161, N28160, N28159, N28158, N28157, N28156, N28155, N28154, N28153, N28152, N28151, N28150, N28149, N28148, N28147, N28146, N28145, N28144, N28143, N28142, N28141, N28140, N28139, N28138, N28137, N28136, N28135, N28134, N28133, N28132, N28131, N28130, N28129, N28128, N28127, N28126, N28125, N28124, N28123, N28122, N28121, N28120, N28119, N28118, N28117, N25400, N25399, N25398, N25397, N25396, N25395, N25394, N25393, N25392, N25391, N25390, N25389, N25388, N25387, N25386, N25385, N25384, N25383, N25382, N25381, N25380, N25379, N25378, N25377, N25376, N25375, N25374, N25373, N25372, N25371, N25370, N25369, N25368, N25367, N25366, N25365, N25364, N25363, N25362, N25361, N25360, N25359, N25358, N25357, N25356, N25355, N25354, N25353, N25352, N25351, N25350, N25349, N25348, N25347, N25346, N25345, N25344, N25343, N25342, N25341, N25340, N25339, N25338, N25337, N24819, N24818, N24817, N24816, N24815, N24814, N24813, N24812, N24811, N24810, N24809, N24808, N24807, N24806, N24805, N24804, N24803, N24802, N24801, N24800, N24799, N24798, N24797, N24796, N24795, N24794, N24793, N24792, N24791, N24790, N24789, N24788, N24787, N24786, N24785, N24784, N24783, N24782, N24781, N24780, N24779, N24778, N24777, N24776, N24775, N24774, N24773, N24772, N24771, N24770, N24769, N24768, N24767, N24766, N24765, N24764, N24763, N24762, N24761, N24760, N24759, N24758, N24757, N24756, N24611, N28116, N28115, N28114, N28113, N28112, N28111, N28110, N28109, N28108, N28107, N28106, N28105, N28104, N28103, N28102, N28101, N28100, N28099, N28098, N28097, N28096, N28095, N28094, N28093, N28092, N28091, N28090, N28089, N28088, N28087, N28086, N28085, N28084, N28083, N28082, N28081, N28080, N28079, N28078, N28077, N28076, N28075, N28074, N28073, N28072, N28071, N28070, N28069, N28068, N28067, N28066, N28065, N28064, N28063, N28062, N28061, N28060, N28059, N28058, N28057, N28056, N28055, N28054, N28053, N28052, N28051, N28050, N28049, N28048, N28047, N28046, N28045, N28044, N28043, N28042, N28041, N28040, N28039, N28038, N28037, N28036, N28035, N28034, N28033, N28032, N28031, N28030, N28029, N28028, N28027, N28026, N28025, N28024, N28023, N28022, N28021, N28020, N28019, N28018, N28017, N28016, N28015, N28014, N28013, N28012, N28011, N28010, N28009, N28008, N28007, N28006, N28005, N28004, N28003, N28002, N28001, N28000, N27999, N27998, N27997, N27996, N27995, N27994, N27993, N27992, N27991, N27990, N27989, N27988, N25336, N25335, N25334, N25333, N25332, N25331, N25330, N25329, N25328, N25327, N25326, N25325, N25324, N25323, N25322, N25321, N25320, N25319, N25318, N25317, N25316, N25315, N25314, N25313, N25312, N25311, N25310, N25309, N25308, N25307, N25306, N25305, N25304, N25303, N25302, N25301, N25300, N25299, N25298, N25297, N25296, N25295, N25294, N25293, N25292, N25291, N25290, N25289, N25288, N25287, N25286, N25285, N25284, N25283, N25282, N25281, N25280, N25279, N25278, N25277, N25276, N25275, N25274, N25273, N24754, N24753, N24752, N24751, N24750, N24749, N24748, N24747, N24746, N24745, N24744, N24743, N24742, N24741, N24740, N24739, N24738, N24737, N24736, N24735, N24734, N24733, N24732, N24731, N24730, N24729, N24728, N24727, N24726, N24725, N24724, N24723, N24722, N24721, N24720, N24719, N24718, N24717, N24716, N24715, N24714, N24713, N24712, N24711, N24710, N24709, N24708, N24707, N24706, N24705, N24704, N24703, N24702, N24701, N24700, N24699, N24698, N24697, N24696, N24695, N24694, N24693, N24692, N24691, N24610, N27987, N27986, N27985, N27984, N27983, N27982, N27981, N27980, N27979, N27978, N27977, N27976, N27975, N27974, N27973, N27972, N27971, N27970, N27969, N27968, N27967, N27966, N27965, N27964, N27963, N27962, N27961, N27960, N27959, N27958, N27957, N27956, N27955, N27954, N27953, N27952, N27951, N27950, N27949, N27948, N27947, N27946, N27945, N27944, N27943, N27942, N27941, N27940, N27939, N27938, N27937, N27936, N27935, N27934, N27933, N27932, N27931, N27930, N27929, N27928, N27927, N27926, N27925, N27924, N27923, N27922, N27921, N27920, N27919, N27918, N27917, N27916, N27915, N27914, N27913, N27912, N27911, N27910, N27909, N27908, N27907, N27906, N27905, N27904, N27903, N27902, N27901, N27900, N27899, N27898, N27897, N27896, N27895, N27894, N27893, N27892, N27891, N27890, N27889, N27888, N27887, N27886, N27885, N27884, N27883, N27882, N27881, N27880, N27879, N27878, N27877, N27876, N27875, N27874, N27873, N27872, N27871, N27870, N27869, N27868, N27867, N27866, N27865, N27864, N27863, N27862, N27861, N27860, N27859, N25272, N25271, N25270, N25269, N25268, N25267, N25266, N25265, N25264, N25263, N25262, N25261, N25260, N25259, N25258, N25257, N25256, N25255, N25254, N25253, N25252, N25251, N25250, N25249, N25248, N25247, N25246, N25245, N25244, N25243, N25242, N25241, N25240, N25239, N25238, N25237, N25236, N25235, N25234, N25233, N25232, N25231, N25230, N25229, N25228, N25227, N25226, N25225, N25224, N25223, N25222, N25221, N25220, N25219, N25218, N25217, N25216, N25215, N25214, N25213, N25212, N25211, N25210, N25209, N24689, N24688, N24687, N24686, N24685, N24684, N24683, N24682, N24681, N24680, N24679, N24678, N24677, N24676, N24675, N24674, N24673, N24672, N24671, N24670, N24669, N24668, N24667, N24666, N24665, N24664, N24663, N24662, N24661, N24660, N24659, N24658, N24657, N24656, N24655, N24654, N24653, N24652, N24651, N24650, N24649, N24648, N24647, N24646, N24645, N24644, N24643, N24642, N24641, N24640, N24639, N24638, N24637, N24636, N24635, N24634, N24633, N24632, N24631, N24630, N24629, N24628, N24627, N24626, N24609, N27858, N27857, N27856, N27855, N27854, N27853, N27852, N27851, N27850, N27849, N27848, N27847, N27846, N27845, N27844, N27843, N27842, N27841, N27840, N27839, N27838, N27837, N27836, N27835, N27834, N27833, N27832, N27831, N27830, N27829, N27828, N27827, N27826, N27825, N27824, N27823, N27822, N27821, N27820, N27819, N27818, N27817, N27816, N27815, N27814, N27813, N27812, N27811, N27810, N27809, N27808, N27807, N27806, N27805, N27804, N27803, N27802, N27801, N27800, N27799, N27798, N27797, N27796, N27795, N27794, N27793, N27792, N27791, N27790, N27789, N27788, N27787, N27786, N27785, N27784, N27783, N27782, N27781, N27780, N27779, N27778, N27777, N27776, N27775, N27774, N27773, N27772, N27771, N27770, N27769, N27768, N27767, N27766, N27765, N27764, N27763, N27762, N27761, N27760, N27759, N27758, N27757, N27756, N27755, N27754, N27753, N27752, N27751, N27750, N27749, N27748, N27747, N27746, N27745, N27744, N27743, N27742, N27741, N27740, N27739, N27738, N27737, N27736, N27735, N27734, N27733, N27732, N27731, N27730, N25208, N25207, N25206, N25205, N25204, N25203, N25202, N25201, N25200, N25199, N25198, N25197, N25196, N25195, N25194, N25193, N25192, N25191, N25190, N25189, N25188, N25187, N25186, N25185, N25184, N25183, N25182, N25181, N25180, N25179, N25178, N25177, N25176, N25175, N25174, N25173, N25172, N25171, N25170, N25169, N25168, N25167, N25166, N25165, N25164, N25163, N25162, N25161, N25160, N25159, N25158, N25157, N25156, N25155, N25154, N25153, N25152, N25151, N25150, N25149, N25148, N25147, N25146, N25145 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N24608)? { N24590, N24589, N24588, N24587, N24586, N24585, N24584, N24583, N24582, N24581, N24580, N24579, N24578, N24577, N24576, N24575, N24574, N24573, N24572, N24571, N24570, N24569, N24568, N24567, N24566, N24565, N24564, N24563, N24562, N24561, N24560, N24559, N24558, N24557, N24556, N24555, N24554, N24553, N24552, N24551, N24550, N24549, N24548, N24547, N24546, N24545, N24544, N24543, N24542, N24541, N24540, N24539, N24538, N24537, N24536, N24535, N24534, N24533, N24532, N24531, N24530, N24529, N24528, N24527, N24526, N24525, N24524, N24523, N24522, N24521, N24520, N24519, N24518, N24517, N24516, N24515, N24514, N24513, N24512, N24511, N24510, N24509, N24508, N24507, N24506, N24505, N24504, N24503, N24502, N24501, N24500, N24499, N24498, N24497, N24496, N24495, N24494, N24493, N24492, N24491, N24490, N24489, N24488, N24487, N24486, N24485, N24484, N24483, N24482, N24481, N24480, N24479, N24478, N24477, N24476, N24475, N24474, N24473, N24472, N24471, N24470, N24469, N24468, N24467, N24466, N24465, N24464, N24463, N24462, N24461, N24460, N24459, N24458, N24457, N24456, N24455, N24454, N24453, N24452, N24451, N24450, N24449, N24448, N24447, N24446, N24445, N24444, N24443, N24442, N24441, N24440, N24439, N24438, N24437, N24436, N24435, N24434, N24433, N24432, N24431, N24430, N24429, N24428, N24427, N24426, N24425, N24424, N24423, N24422, N24421, N24420, N24419, N24418, N24417, N24416, N24415, N24414, N24413, N24412, N24411, N24410, N24409, N24408, N24407, N24406, N24405, N24404, N24403, N24402, N24401, N24400, N24399, N24398, N24397, N24396, N24395, N24394, N24393, N24392, N24391, N24390, N24389, N24388, N24387, N24386, N24385, N24384, N24383, N24382, N24381, N24380, N24379, N24378, N24377, N24376, N24375, N24374, N24373, N24372, N24371, N24370, N24369, N24368, N24367, N24366, N24365, N24364, N24363, N24362, N24361, N24360, N24359, N24358, N24357, N24356, N24355, N24354, N24353, N24352, N24351, N24350, N24349, N24348, N24347, N24346, N24345, N24344, N24343, N24342, N24341, N24340, N24339, N24338, N24337, N24336, N24335, N24334, N24333, N24332, N24331, N24330, N24329, N24328, N24327, N24326, N24325, N24324, N24323, N24322, N24321, N24320, N24319, N24318, N24317, N24316, N24315, N24314, N24313, N24312, N24311, N24310, N24309, N24308, N24307, N24306, N24305, N24304, N24303, N24302, N24301, N24300, N24299, N24298, N24297, N24296, N24295, N24294, N24293, N24292, N24291, N24290, N24289, N24288, N24287, N24286, N24285, N24284, N24283, N24282, N24281, N24280, N24279, N24278, N24277, N24276, N24275, N24274, N24273, N24272, N24271, N24270, N24269, N24268, N24267, N24266, N24265, N24264, N24263, N24262, N24261, N24260, N24259, N24258, N24257, N24256, N24255, N24254, N24253, N24252, N24251, N24250, N24249, N24248, N24247, N24246, N24245, N24244, N24243, N24242, N24241, N24240, N24239, N24238, N24237, N24236, N24235, N24234, N24233, N24232, N24231, N24230, N24229, N24228, N24227, N24226, N24225, N24224, N24223, N24222, N24221, N24220, N24219, N24218, N24217, N24216, N24215, N24214, N24213, N24212, N24211, N24210, N24209, N24208, N24207, N24206, N24205, N24204, N24203, N24202, N24201, N24200, N24199, N24198, N24197, N24196, N24195, N24194, N24193, N24192, N24191, N24190, N24189, N24188, N24187, N24186, N24185, N24184, N24183, N24182, N24181, N24180, N24179, N24178, N24177, N24176, N24175, N24174, N24173, N24172, N24171, N24170, N24169, N24168, N24167, N24166, N24165, N24164, N24163, N24162, N24161, N24160, N24159, N24158, N24157, N24156, N24155, N24154, N24153, N24152, N24151, N24150, N24149, N24148, N24147, N24146, N24145, N24144, N24143, N24142, N24141, N24140, N24139, N24138, N24137, N24136, N24135, N24134, N24133, N24132, N24131, N24130, N24129, N24128, N24127, N24126, N24125, N24124, N24123, N24122, N24121, N24120, N24119, N24118, N24117, N24116, N24115, N24114, N24113, N24112, N24111, N24110, N24109, N24108, N24107, N24106, N24105, N24104, N24103, N24102, N24101, N24100, N24099, N24098, N24097, N24096, N24095, N24094, N24093, N24092, N24091, N24090, N24089, N24088, N24087, N24086, N24085, N24084, N24083, N24082, N24081, N24080, N24079, N24078, N24077, N24076, N24075, N24074, N24073, N24072, N24071, N24070, N24069, N24068, N24067, N24066, N24065, N24064, N24063, N24062, N24061, N24060, N24059, N24058, N24057, N24056, N24055, N24054, N24053, N24052, N24051, N24050, N24049, N24048, N24047, N24046, N24045, N24044, N24043, N24042, N24041, N24040, N24039, N24038, N24037, N24036, N24035, N24034, N24033, N24032, N24031, N24030, N24029, N24028, N24027, N24026, N24025, N24024, N24023, N24022, N24021, N24020, N24019, N24018, N24017, N24016, N24015, N24014, N24013, N24012, N24011, N24010, N24009, N24008, N24007, N24006, N24005, N24004, N24003, N24002, N24001, N24000, N23999, N23998, N23997, N23996, N23995, N23994, N23993, N23992, N23991, N23990, N23989, N23988, N23987, N23986, N23985, N23984, N23983, N23982, N23981, N23980, N23979, N23978, N23977, N23976, N23975, N23974, N23973, N23972, N23971, N23970, N23969, N23968, N23967, N23966, N23965, N23964, N23963, N23962, N23961, N23960, N23959, N23958, N23957, N23956, N23955, N23954, N23953, N23952, N23951, N23950, N23949, N23948, N23947, N23946, N23945, N23944, N23943, N23942, N23941, N23940, N23939, N23938, N23937, N23936, N23935, N23934, N23933, N23932, N23931, N23930, N23929, N23928, N23927, N23926, N23925, N23924, N23923, N23922, N23921, N23920, N23919, N23918, N23917, N23916, N23915, N23914, N23913, N23912, N23911, N23910, N23909, N23908, N23907, N23906, N23905, N23904, N23903, N23902, N23901, N23900, N23899, N23898, N23897, N23896, N23895, N23894, N23893, N23892, N23891, N23890, N23889, N23888, N23887, N23886, N23885, N23884, N23883, N23882, N23881, N23880, N23879, N23878, N23877, N23876, N23875, N23874, N23873, N23872, N23871, N23870, N23869, N23868, N23867, N23866, N23865, N23864, N23863, N23862, N23861, N23860, N23859, N23858, N23857, N23856, N23855, N23854, N23853, N23852, N23851, N23850, N23849, N23848, N23847, N23846, N23845, N23844, N23843, N23842, N23841, N23840, N23839, N23838, N23837, N23836, N23835, N23834, N23833, N23832, N23831, N23830, N23829, N23828, N23827, N23826, N23825, N23824, N23823, N23822, N23821, N23820, N23819, N23818, N23817, N23816, N23815, N23814, N23813, N23812, N23811, N23810, N23809, N23808, N23807, N23806, N23805, N23804, N23803, N23802, N23801, N23800, N23799, N23798, N23797, N23796, N23795, N23794, N23793, N23792, N23791, N23790, N23789, N23788, N23787, N23786, N23785, N23784, N23783, N23782, N23781, N23780, N23779, N23778, N23777, N23776, N23775, N23774, N23773, N23772, N23771, N23770, N23769, N23768, N23767, N23766, N23765, N23764, N23763, N23762, N23761, N23760, N23759, N23758, N23757, N23756, N23755, N23754, N23753, N23752, N23751, N23750, N23749, N23748, N23747, N23746, N23745, N23744, N23743, N23742, N23741, N23740, N23739, N23738, N23737, N23736, N23735, N23734, N23733, N23732, N23731, N23730, N23729, N23728, N23727, N23726, N23725, N23724, N23723, N23722, N23721, N23720, N23719, N23718, N23717, N23716, N23715, N23714, N23713, N23712, N23711, N23710, N23709, N23708, N23707, N23706, N23705, N23704, N23703, N23702, N23701, N23700, N23699, N23698, N23697, N23696, N23695, N23694, N23693, N23692, N23691, N23690, N23689, N23688, N23687, N23686, N23685, N23684, N23683, N23682, N23681, N23680, N23679, N23678, N23677, N23676, N23675, N23674, N23673, N23672, N23671, N23670, N23669, N23668, N23667, N23666, N23665, N23664, N23663, N23662, N23661, N23660, N23659, N23658, N23657, N23656, N23655, N23654, N23653, N23652, N23651, N23650, N23649, N23648, N23647, N23646, N23645, N23644, N23643, N23642, N23641, N23640, N23639, N23638, N23637, N23636, N23635, N23634, N23633, N23632, N23631, N23630, N23629, N23628, N23627, N23626, N23625, N23624, N23623, N23622, N23621, N23620, N23619, N23618, N23617, N23616, N23615, N23614, N23613, N23612, N23611, N23610, N23609, N23608, N23607, N23606, N23605, N23604, N23603, N23602, N23601, N23600, N23599, N23598, N23597, N23596, N23595, N23594, N23593, N23592, N23591, N23590, N23589, N23588, N23587, N23586, N23585, N23584, N23583, N23582, N23581, N23580, N23579, N23578, N23577, N23576, N23575, N23574, N23573, N23572, N23571, N23570, N23569, N23568, N23567, N23566, N23565, N23564, N23563, N23562, N23561, N23560, N23559, N23558, N23557, N23556, N23555, N23554, N23553, N23552, N23551, N23550, N23549, N23548, N23547, N23546, N23545, N23544, N23543, N23542, N23541, N23540, N23539, N23538, N23537, N23536, N23535, N23534, N23533, N23532, N23531, N23530, N23529, N23528, N23527, N23526, N23525, N23524, N23523, N23522, N23521, N23520, N23519, N23518, N23517, N23516, N23515, N23514, N23513, N23512, N23511, N23510, N23509, N23508, N23507, N23506, N23505, N23504, N23503, N23502, N23501, N23500, N23499, N23498, N23497, N23496, N23495, N23494, N23493, N23492, N23491, N23490, N23489, N23488, N23487, N23486, N23485, N23484, N23483, N23482, N23481, N23480, N23479, N23478, N23477, N23476, N23475, N23474, N23473, N23472, N23471, N23470, N23469, N23468, N23467, N23466, N23465, N23464, N23463, N23462, N23461, N23460, N23459, N23458, N23457, N23456, N23455, N23454, N23453, N23452, N23451, N23450, N23449, N23448, N23447, N23446, N23445, N23444, N23443, N23442, N23441, N23440, N23439, N23438, N23437, N23436, N23435, N23434, N23433, N23432, N23431, N23430, N23429, N23428, N23427, N23426, N23425, N23424, N23423, N23422, N23421, N23420, N23419, N23418, N23417, N23416, N23415, N23414, N23413, N23412, N23411, N23410, N23409, N23408, N23407, N23406, N23405, N23404, N23403, N23402, N23401, N23400, N23399, N23398, N23397, N23396, N23395, N23394, N23393, N23392, N23391, N23390, N23389, N23388, N23387, N23386, N23385, N23384, N23383, N23382, N23381, N23380, N23379, N23378, N23377, N23376, N23375, N23374, N23373, N23372, N23371, N23370, N23369, N23368, N23367, N23366, N23365, N23364, N23363, N23362, N23361, N23360, N23359, N23358, N23357, N23356, N23355, N23354, N23353, N23352, N23351, N23350, N23349, N23348, N23347, N23346, N23345, N23344, N23343, N23342, N23341, N23340, N23339, N23338, N23337, N23336, N23335, N23334, N23333, N23332, N23331, N23330, N23329, N23328, N23327, N23326, N23325, N23324, N23323, N23322, N23321, N23320, N23319, N23318, N23317, N23316, N23315, N23314, N23313, N23312, N23311, N23310, N23309, N23308, N23307, N23306, N23305, N23304, N23303, N23302, N23301, N23300, N23299, N23298, N23297, N23296, N23295, N23294, N23293, N23292, N23291, N23290, N23289, N23288, N23287, N23286, N23285, N23284, N23283, N23282, N23281, N23280, N23279, N23278, N23277, N23276, N23275, N23274, N23273, N23272, N23271, N23270, N23269, N23268, N23267, N23266, N23265, N23264, N23263, N23262, N23261, N23260, N23259, N23258, N23257, N23256, N23255, N23254, N23253, N23252, N23251, N23250, N23249, N23248, N23247, N23246, N23245, N23244, N23243, N23242, N23241, N23240, N23239, N23238, N23237, N23236, N23235, N23234, N23233, N23232, N23231, N23230, N23229, N23228, N23227, N23226, N23225, N23224, N23223, N23222, N23221, N23220, N23219, N23218, N23217, N23216, N23215, N23214, N23213, N23212, N23211, N23210, N23209, N23208, N23207, N23206, N23205, N23204, N23203, N23202, N23201, N23200, N23199, N23198, N23197, N23196, N23195, N23194, N23193, N23192, N23191, N23190, N23189, N23188, N23187, N23186, N23185, N23184, N23183, N23182, N23181, N23180, N23179, N23178, N23177, N23176, N23175, N23174, N23173, N23172, N23171, N23170, N23169, N23168, N23167, N23166, N23165, N23164, N23163, N23162, N23161, N23160, N23159, N23158, N23157, N23156, N23155, N23154, N23153, N23152, N23151, N23150, N23149, N23148, N23147, N23146, N23145, N23144, N23143, N23142, N23141, N23140, N23139, N23138, N23137, N23136, N23135, N23134, N23133, N23132, N23131, N23130, N23129, N23128, N23127, N23126, N23125, N23124, N23123, N23122, N23121, N23120, N23119, N23118, N23117, N23116, N23115, N23114, N23113, N23112, N23111, N23110, N23109, N23108, N23107, N23106, N23105, N23104, N23103, N23102, N23101, N23100, N23099, N23098, N23097, N23096, N23095, N23094, N23093, N23092, N23091, N23090, N23089, N23088, N23087, N23086, N23085, N23084, N23083, N23082, N23081, N23080, N23079, N23078, N23077, N23076, N23075, N23074, N23073, N23072, N23071, N23070, N23069, N23068, N23067, N23066, N23065, N23064, N23063, N23062, N23061, N23060, N23059, N23058, N23057, N23056, N23055, N23054, N23053, N23052, N23051, N23050, N23049, N23048, N23047, N23046, N23045, N23044, N23043, N23042, N23041, N23040, N23039, N23038, N23037, N23036, N23035, N23034, N23033, N23032, N23031, N23030, N23029, N23028, N23027, N23026, N23025, N23024, N23023, N23022, N23021, N23020, N23019, N23018, N23017, N23016, N23015, N23014, N23013, N23012, N23011, N23010, N23009, N23008, N23007, N23006, N23005, N23004, N23003, N23002, N23001, N23000, N22999, N22998, N22997, N22996, N22995, N22994, N22993, N22992, N22991, N22990, N22989, N22988, N22987, N22986, N22985, N22984, N22983, N22982, N22981, N22980, N22979, N22978, N22977, N22976, N22975, N22974, N22973, N22972, N22971, N22970, N22969, N22968, N22967, N22966, N22965, N22964, N22963, N22962, N22961, N22960, N22959, N22958, N22957, N22956, N22955, N22954, N22953, N22952, N22951, N22950, N22949, N22948, N22947, N22946, N22945, N22944, N22943, N22942, N22941, N22940, N22939, N22938, N22937, N22936, N22935, N22934, N22933, N22932, N22931, N22930, N22929, N22928, N22927, N22926, N22925, N22924, N22923, N22922, N22921, N22920, N22919, N22918, N22917, N22916, N22915, N22914, N22913, N22912, N22911, N22910, N22909, N22908, N22907, N22906, N22905, N22904, N22903, N22902, N22901, N22900, N22899, N22898, N22897, N22896, N22895, N22894, N22893, N22892, N22891, N22890, N22889, N22888, N22887, N22886, N22885, N22884, N22883, N22882, N22881, N22880, N22879, N22878, N22877, N22876, N22875, N22874, N22873, N22872, N22871, N22870, N22869, N22868, N22867, N22866, N22865, N22864, N22863, N22862, N22861, N22860, N22859, N22858, N22857, N22856, N22855, N22854, N22853, N22852, N22851, N22850, N22849, N22848, N22847, N22846, N22845, N22844, N22843, N22842, N22841, N22840, N22839, N22838, N22837, N22836, N22835, N22834, N22833, N22832, N22831, N22830, N22829, N22828, N22827, N22826, N22825, N22824, N22823, N22822, N22821, N22820, N22819, N22818, N22817, N22816, N22815, N22814, N22813, N22812, N22811, N22810, N22809, N22808, N22807, N22806, N22805, N22804, N22803, N22802, N22801, N22800, N22799, N22798, N22797, N22796, N22795, N22794, N22793, N22792, N22791, N22790, N22789, N22788, N22787, N22786, N22785, N22784, N22783, N22782, N22781, N22780, N22779, N22778, N22777, N22776, N22775, N22774, N22773, N22772, N22771, N22770, N22769, N22768, N22767, N22766, N22765, N22764, N22763, N22762, N22761, N22760, N22759, N22758, N22757, N22756, N22755, N22754, N22753, N22752, N22751, N22750, N22749, N22748, N22747, N22746, N22745, N22744, N22743, N22742, N22741, N22740, N22739, N22738, N22737, N22736, N22735, N22734, N22733, N22732, N22731, N22730, N22729, N22728, N22727, N22726, N22725, N22724, N22723, N22722, N22721, N22720, N22719, N22718, N22717, N22716, N22715, N22714, N22713, N22712, N22711, N22710, N22709, N22708, N22707, N22706, N22705, N22704, N22703, N22702, N22701, N22700, N22699, N22698, N22697, N22696, N22695, N22694, N22693, N22692, N22691, N22690, N22689, N22688, N22687, N22686, N22685, N22684, N22683, N22682, N22681, N22680, N22679, N22678, N22677, N22676, N22675, N22674, N22673, N22672, N22671, N22670, N22669, N22668, N22667, N22666, N22665, N22664, N22663, N22662, N22661, N22660, N22659, N22658, N22657, N22656, N22655, N22654, N22653, N22652, N22651, N22650, N22649, N22648, N22647, N22646, N22645, N22644, N22643, N22642, N22641, N22640, N22639, N22638, N22637, N22636, N22635, N22634, N22633, N22632, N22631, N22630, N22629, N22628, N22627, N22626, N22625, N22624, N22623, N22622, N22621, N22620, N22619, N22618, N22617, N22616, N22615, N22614, N22613, N22612, N22611, N22610, N22609, N22608, N22607, N22606, N22605, N22604, N22603, N22602, N22601, N22600, N22599, N22598, N22597, N22596, N22595, N22594, N22593, N22592, N22591, N22590, N22589, N22588, N22587, N22586, N22585, N22584, N22583, N22582, N22581, N22580, N22579, N22578, N22577, N22576, N22575, N22574, N22573, N22572, N22571, N22570, N22569, N22568, N22567, N22566, N22565, N22564, N22563, N22562, N22561, N22560, N22559, N22558, N22557, N22556, N22555, N22554, N22553, N22552, N22551, N22550, N22549, N22548, N22547, N22546, N22545, N22544, N22543, N22542, N22541, N22540, N22539, N22538, N22537, N22536, N22535, N22534, N22533, N22532, N22531, N22530, N22529, N22528, N22527 } : 1'b0;
  assign N204 = N24607;
  assign N28789 = (N205)? 1'b0 : 
                  (N28788)? N4072 : 1'b0;
  assign N205 = N28780;
  assign N28791 = (N206)? 1'b0 : 
                  (N28790)? N4331 : 1'b0;
  assign N206 = N28781;
  assign N28793 = (N207)? 1'b0 : 
                  (N28792)? N4590 : 1'b0;
  assign N207 = N28782;
  assign N28795 = (N208)? 1'b0 : 
                  (N28794)? N4849 : 1'b0;
  assign N208 = N28783;
  assign N28797 = (N209)? 1'b0 : 
                  (N28796)? N5108 : 1'b0;
  assign N209 = N28784;
  assign N28799 = (N210)? 1'b0 : 
                  (N28798)? N5367 : 1'b0;
  assign N210 = N28785;
  assign N28801 = (N211)? 1'b0 : 
                  (N28800)? N5626 : 1'b0;
  assign N211 = N28786;
  assign N28803 = (N212)? 1'b0 : 
                  (N28802)? N5885 : 1'b0;
  assign N212 = N28787;
  assign N28813 = (N213)? 1'b0 : 
                  (N28812)? N28763 : 1'b0;
  assign N213 = N28804;
  assign N28815 = (N214)? 1'b0 : 
                  (N28814)? N28765 : 1'b0;
  assign N214 = N28805;
  assign N28817 = (N215)? 1'b0 : 
                  (N28816)? N28767 : 1'b0;
  assign N215 = N28806;
  assign N28819 = (N216)? 1'b0 : 
                  (N28818)? N28769 : 1'b0;
  assign N216 = N28807;
  assign N28821 = (N217)? 1'b0 : 
                  (N28820)? N28771 : 1'b0;
  assign N217 = N28808;
  assign N28823 = (N218)? 1'b0 : 
                  (N28822)? N28773 : 1'b0;
  assign N218 = N28809;
  assign N28825 = (N219)? 1'b0 : 
                  (N28824)? N28775 : 1'b0;
  assign N219 = N28810;
  assign N28827 = (N220)? 1'b0 : 
                  (N28826)? N28777 : 1'b0;
  assign N220 = N28811;
  assign { N28849, N28848, N28847, N28846, N28845, N28844, N28843, N28842, N28841, N28840, N28839, N28838, N28837, N28836, N28835, N28834 } = (N221)? { N28803, N28827, N28801, N28825, N28799, N28823, N28797, N28821, N28795, N28819, N28793, N28817, N28791, N28815, N28789, N28813 } : 
                                                                                                                                              (N28778)? { N5885, N28777, N5626, N28775, N5367, N28773, N5108, N28771, N4849, N28769, N4590, N28767, N4331, N28765, N4072, N28763 } : 1'b0;
  assign N221 = commit_ack_i[0];
  assign { N28852, N28851, N28850 } = (N221)? { N28830, N28829, N28828 } : 
                                      (N28778)? commit_pointer_q : 1'b0;
  assign N28867 = (N222)? 1'b0 : 
                  (N28866)? N28835 : 1'b0;
  assign N222 = N28858;
  assign N28869 = (N223)? 1'b0 : 
                  (N28868)? N28837 : 1'b0;
  assign N223 = N28859;
  assign N28871 = (N224)? 1'b0 : 
                  (N28870)? N28839 : 1'b0;
  assign N224 = N28860;
  assign N28873 = (N225)? 1'b0 : 
                  (N28872)? N28841 : 1'b0;
  assign N225 = N28861;
  assign N28875 = (N226)? 1'b0 : 
                  (N28874)? N28843 : 1'b0;
  assign N226 = N28862;
  assign N28877 = (N227)? 1'b0 : 
                  (N28876)? N28845 : 1'b0;
  assign N227 = N28863;
  assign N28879 = (N228)? 1'b0 : 
                  (N28878)? N28847 : 1'b0;
  assign N228 = N28864;
  assign N28881 = (N229)? 1'b0 : 
                  (N28880)? N28849 : 1'b0;
  assign N229 = N28865;
  assign N28894 = (N230)? 1'b0 : 
                  (N28893)? N28834 : 1'b0;
  assign N230 = N28885;
  assign N28896 = (N231)? 1'b0 : 
                  (N28895)? N28836 : 1'b0;
  assign N231 = N28886;
  assign N28898 = (N232)? 1'b0 : 
                  (N28897)? N28838 : 1'b0;
  assign N232 = N28887;
  assign N28900 = (N233)? 1'b0 : 
                  (N28899)? N28840 : 1'b0;
  assign N233 = N28888;
  assign N28902 = (N234)? 1'b0 : 
                  (N28901)? N28842 : 1'b0;
  assign N234 = N28889;
  assign N28904 = (N235)? 1'b0 : 
                  (N28903)? N28844 : 1'b0;
  assign N235 = N28890;
  assign N28906 = (N236)? 1'b0 : 
                  (N28905)? N28846 : 1'b0;
  assign N236 = N28891;
  assign N28908 = (N237)? 1'b0 : 
                  (N28907)? N28848 : 1'b0;
  assign N237 = N28892;
  assign { N28930, N28929, N28928, N28927, N28926, N28925, N28924, N28923, N28922, N28921, N28920, N28919, N28918, N28917, N28916, N28915 } = (N238)? { N28881, N28908, N28879, N28906, N28877, N28904, N28875, N28902, N28873, N28900, N28871, N28898, N28869, N28896, N28867, N28894 } : 
                                                                                                                                              (N28853)? { N28849, N28848, N28847, N28846, N28845, N28844, N28843, N28842, N28841, N28840, N28839, N28838, N28837, N28836, N28835, N28834 } : 1'b0;
  assign N238 = commit_ack_i[1];
  assign { N28933, N28932, N28931 } = (N238)? { N28911, N28910, N28909 } : 
                                      (N28853)? { N28852, N28851, N28850 } : 1'b0;
  assign issue_pointer_n = (N239)? { 1'b0, 1'b0, 1'b0 } : 
                           (N240)? { N3810, N3809, N3808 } : 1'b0;
  assign N239 = flush_i;
  assign N240 = N28934;
  assign commit_pointer_n = (N239)? { 1'b0, 1'b0, 1'b0 } : 
                            (N240)? { N28933, N28932, N28931 } : 1'b0;
  assign { mem_n[2903:2903], mem_n[2742:2742], mem_n[2610:2610], mem_n[2540:2540], mem_n[2379:2379], mem_n[2247:2247], mem_n[2177:2177], mem_n[2016:2016], mem_n[1884:1884], mem_n[1814:1814], mem_n[1653:1653], mem_n[1521:1521], mem_n[1451:1451], mem_n[1290:1290], mem_n[1158:1158], mem_n[1088:1088], mem_n[927:927], mem_n[795:795], mem_n[725:725], mem_n[564:564], mem_n[432:432], mem_n[362:362], mem_n[201:201], mem_n[69:69] } = (N239)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                            (N240)? { N28930, N28929, N28776, N28928, N28927, N28774, N28926, N28925, N28772, N28924, N28923, N28770, N28922, N28921, N28768, N28920, N28919, N28766, N28918, N28917, N28764, N28916, N28915, N28762 } : 1'b0;
  assign issue_cnt_n = (N239)? { 1'b0, 1'b0, 1'b0 } : 
                       (N240)? { N28914, N28913, N28912 } : 1'b0;
  assign { N29003, N29002, N29001, N29000 } = (N241)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N28999)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N241 = N28936;
  assign { N29008, N29007, N29006, N29005 } = (N242)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29004)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N242 = N28937;
  assign { N29013, N29012, N29011, N29010 } = (N243)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29009)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N243 = N28938;
  assign { N29018, N29017, N29016, N29015 } = (N244)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29014)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N244 = N28939;
  assign { N29023, N29022, N29021, N29020 } = (N245)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29019)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N245 = N28940;
  assign { N29028, N29027, N29026, N29025 } = (N246)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29024)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N246 = N28941;
  assign { N29033, N29032, N29031, N29030 } = (N247)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29029)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N247 = N28942;
  assign { N29038, N29037, N29036, N29035 } = (N248)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29034)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N248 = N28943;
  assign { N29043, N29042, N29041, N29040 } = (N249)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29039)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N249 = N28944;
  assign { N29048, N29047, N29046, N29045 } = (N250)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29044)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N250 = N28945;
  assign { N29053, N29052, N29051, N29050 } = (N251)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29049)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N251 = N28946;
  assign { N29058, N29057, N29056, N29055 } = (N252)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29054)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N252 = N28947;
  assign { N29063, N29062, N29061, N29060 } = (N253)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29059)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N253 = N28948;
  assign { N29068, N29067, N29066, N29065 } = (N254)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29064)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N254 = N28949;
  assign { N29073, N29072, N29071, N29070 } = (N255)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29069)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N255 = N28950;
  assign { N29078, N29077, N29076, N29075 } = (N256)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29074)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N256 = N28951;
  assign { N29083, N29082, N29081, N29080 } = (N257)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29079)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N257 = N28952;
  assign { N29088, N29087, N29086, N29085 } = (N258)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29084)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N258 = N28953;
  assign { N29093, N29092, N29091, N29090 } = (N259)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29089)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N259 = N28954;
  assign { N29098, N29097, N29096, N29095 } = (N260)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29094)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N260 = N28955;
  assign { N29103, N29102, N29101, N29100 } = (N261)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29099)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N261 = N28956;
  assign { N29108, N29107, N29106, N29105 } = (N262)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29104)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N262 = N28957;
  assign { N29113, N29112, N29111, N29110 } = (N263)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29109)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N263 = N28958;
  assign { N29118, N29117, N29116, N29115 } = (N264)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29114)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N264 = N28959;
  assign { N29123, N29122, N29121, N29120 } = (N265)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29119)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N265 = N28960;
  assign { N29128, N29127, N29126, N29125 } = (N266)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29124)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N266 = N28961;
  assign { N29133, N29132, N29131, N29130 } = (N267)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29129)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N267 = N28962;
  assign { N29138, N29137, N29136, N29135 } = (N268)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29134)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N268 = N28963;
  assign { N29143, N29142, N29141, N29140 } = (N269)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29139)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N269 = N28964;
  assign { N29148, N29147, N29146, N29145 } = (N270)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29144)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N270 = N28965;
  assign { N29153, N29152, N29151, N29150 } = (N271)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29149)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N271 = N28966;
  assign { N29158, N29157, N29156, N29155 } = (N272)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29154)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N272 = N28967;
  assign { N29163, N29162, N29161, N29160 } = (N273)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29159)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N273 = N28968;
  assign { N29168, N29167, N29166, N29165 } = (N274)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29164)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N274 = N28969;
  assign { N29173, N29172, N29171, N29170 } = (N275)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29169)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N275 = N28970;
  assign { N29178, N29177, N29176, N29175 } = (N276)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29174)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N276 = N28971;
  assign { N29183, N29182, N29181, N29180 } = (N277)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29179)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N277 = N28972;
  assign { N29188, N29187, N29186, N29185 } = (N278)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29184)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N278 = N28973;
  assign { N29193, N29192, N29191, N29190 } = (N279)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29189)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N279 = N28974;
  assign { N29198, N29197, N29196, N29195 } = (N280)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29194)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N280 = N28975;
  assign { N29203, N29202, N29201, N29200 } = (N281)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29199)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N281 = N28976;
  assign { N29208, N29207, N29206, N29205 } = (N282)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29204)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N282 = N28977;
  assign { N29213, N29212, N29211, N29210 } = (N283)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29209)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N283 = N28978;
  assign { N29218, N29217, N29216, N29215 } = (N284)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29214)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N284 = N28979;
  assign { N29223, N29222, N29221, N29220 } = (N285)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29219)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N285 = N28980;
  assign { N29228, N29227, N29226, N29225 } = (N286)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29224)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N286 = N28981;
  assign { N29233, N29232, N29231, N29230 } = (N287)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29229)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N287 = N28982;
  assign { N29238, N29237, N29236, N29235 } = (N288)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29234)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N288 = N28983;
  assign { N29243, N29242, N29241, N29240 } = (N289)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29239)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N289 = N28984;
  assign { N29248, N29247, N29246, N29245 } = (N290)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29244)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N290 = N28985;
  assign { N29253, N29252, N29251, N29250 } = (N291)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29249)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N291 = N28986;
  assign { N29258, N29257, N29256, N29255 } = (N292)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29254)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N292 = N28987;
  assign { N29263, N29262, N29261, N29260 } = (N293)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29259)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N293 = N28988;
  assign { N29268, N29267, N29266, N29265 } = (N294)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29264)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N294 = N28989;
  assign { N29273, N29272, N29271, N29270 } = (N295)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29269)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N295 = N28990;
  assign { N29278, N29277, N29276, N29275 } = (N296)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29274)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N296 = N28991;
  assign { N29283, N29282, N29281, N29280 } = (N297)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29279)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N297 = N28992;
  assign { N29288, N29287, N29286, N29285 } = (N298)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29284)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N298 = N28993;
  assign { N29293, N29292, N29291, N29290 } = (N299)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29289)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N299 = N28994;
  assign { N29298, N29297, N29296, N29295 } = (N300)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29294)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N300 = N28995;
  assign { N29303, N29302, N29301, N29300 } = (N301)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29299)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N301 = N28996;
  assign { N29308, N29307, N29306, N29305 } = (N302)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29304)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N302 = N28997;
  assign { N29313, N29312, N29311, N29310 } = (N303)? { mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294] } : 
                                              (N29309)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N303 = N28998;
  assign { N29565, N29564, N29563, N29562, N29561, N29560, N29559, N29558, N29557, N29556, N29555, N29554, N29553, N29552, N29551, N29550, N29549, N29548, N29547, N29546, N29545, N29544, N29543, N29542, N29541, N29540, N29539, N29538, N29537, N29536, N29535, N29534, N29533, N29532, N29531, N29530, N29529, N29528, N29527, N29526, N29525, N29524, N29523, N29522, N29521, N29520, N29519, N29518, N29517, N29516, N29515, N29514, N29513, N29512, N29511, N29510, N29509, N29508, N29507, N29506, N29505, N29504, N29503, N29502, N29501, N29500, N29499, N29498, N29497, N29496, N29495, N29494, N29493, N29492, N29491, N29490, N29489, N29488, N29487, N29486, N29485, N29484, N29483, N29482, N29481, N29480, N29479, N29478, N29477, N29476, N29475, N29474, N29473, N29472, N29471, N29470, N29469, N29468, N29467, N29466, N29465, N29464, N29463, N29462, N29461, N29460, N29459, N29458, N29457, N29456, N29455, N29454, N29453, N29452, N29451, N29450, N29449, N29448, N29447, N29446, N29445, N29444, N29443, N29442, N29441, N29440, N29439, N29438, N29437, N29436, N29435, N29434, N29433, N29432, N29431, N29430, N29429, N29428, N29427, N29426, N29425, N29424, N29423, N29422, N29421, N29420, N29419, N29418, N29417, N29416, N29415, N29414, N29413, N29412, N29411, N29410, N29409, N29408, N29407, N29406, N29405, N29404, N29403, N29402, N29401, N29400, N29399, N29398, N29397, N29396, N29395, N29394, N29393, N29392, N29391, N29390, N29389, N29388, N29387, N29386, N29385, N29384, N29383, N29382, N29381, N29380, N29379, N29378, N29377, N29376, N29375, N29374, N29373, N29372, N29371, N29370, N29369, N29368, N29367, N29366, N29365, N29364, N29363, N29362, N29361, N29360, N29359, N29358, N29357, N29356, N29355, N29354, N29353, N29352, N29351, N29350, N29349, N29348, N29347, N29346, N29345, N29344, N29343, N29342, N29341, N29340, N29339, N29338, N29337, N29336, N29335, N29334, N29333, N29332, N29331, N29330, N29329, N29328, N29327, N29326, N29325, N29324, N29323, N29322, N29321, N29320, N29319, N29318, N29317, N29316, N29315, N29314 } = (N304)? { N29310, N29311, N29312, N29313, N29305, N29306, N29307, N29308, N29300, N29301, N29302, N29303, N29295, N29296, N29297, N29298, N29290, N29291, N29292, N29293, N29285, N29286, N29287, N29288, N29280, N29281, N29282, N29283, N29275, N29276, N29277, N29278, N29270, N29271, N29272, N29273, N29265, N29266, N29267, N29268, N29260, N29261, N29262, N29263, N29255, N29256, N29257, N29258, N29250, N29251, N29252, N29253, N29245, N29246, N29247, N29248, N29240, N29241, N29242, N29243, N29235, N29236, N29237, N29238, N29230, N29231, N29232, N29233, N29225, N29226, N29227, N29228, N29220, N29221, N29222, N29223, N29215, N29216, N29217, N29218, N29210, N29211, N29212, N29213, N29205, N29206, N29207, N29208, N29200, N29201, N29202, N29203, N29195, N29196, N29197, N29198, N29190, N29191, N29192, N29193, N29185, N29186, N29187, N29188, N29180, N29181, N29182, N29183, N29175, N29176, N29177, N29178, N29170, N29171, N29172, N29173, N29165, N29166, N29167, N29168, N29160, N29161, N29162, N29163, N29155, N29156, N29157, N29158, N29150, N29151, N29152, N29153, N29145, N29146, N29147, N29148, N29140, N29141, N29142, N29143, N29135, N29136, N29137, N29138, N29130, N29131, N29132, N29133, N29125, N29126, N29127, N29128, N29120, N29121, N29122, N29123, N29115, N29116, N29117, N29118, N29110, N29111, N29112, N29113, N29105, N29106, N29107, N29108, N29100, N29101, N29102, N29103, N29095, N29096, N29097, N29098, N29090, N29091, N29092, N29093, N29085, N29086, N29087, N29088, N29080, N29081, N29082, N29083, N29075, N29076, N29077, N29078, N29070, N29071, N29072, N29073, N29065, N29066, N29067, N29068, N29060, N29061, N29062, N29063, N29055, N29056, N29057, N29058, N29050, N29051, N29052, N29053, N29045, N29046, N29047, N29048, N29040, N29041, N29042, N29043, N29035, N29036, N29037, N29038, N29030, N29031, N29032, N29033, N29025, N29026, N29027, N29028, N29020, N29021, N29022, N29023, N29015, N29016, N29017, N29018, N29010, N29011, N29012, N29013, N29005, N29006, N29007, N29008, N29000, N29001, N29002, N29003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N28935)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N304 = mem_q[362];
  assign { N29634, N29633, N29632, N29631 } = (N305)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29630)? { N29314, N29315, N29316, N29317 } : 1'b0;
  assign N305 = N29567;
  assign { N29639, N29638, N29637, N29636 } = (N306)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29635)? { N29318, N29319, N29320, N29321 } : 1'b0;
  assign N306 = N29568;
  assign { N29644, N29643, N29642, N29641 } = (N307)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29640)? { N29322, N29323, N29324, N29325 } : 1'b0;
  assign N307 = N29569;
  assign { N29649, N29648, N29647, N29646 } = (N308)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29645)? { N29326, N29327, N29328, N29329 } : 1'b0;
  assign N308 = N29570;
  assign { N29654, N29653, N29652, N29651 } = (N309)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29650)? { N29330, N29331, N29332, N29333 } : 1'b0;
  assign N309 = N29571;
  assign { N29659, N29658, N29657, N29656 } = (N310)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29655)? { N29334, N29335, N29336, N29337 } : 1'b0;
  assign N310 = N29572;
  assign { N29664, N29663, N29662, N29661 } = (N311)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29660)? { N29338, N29339, N29340, N29341 } : 1'b0;
  assign N311 = N29573;
  assign { N29669, N29668, N29667, N29666 } = (N312)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29665)? { N29342, N29343, N29344, N29345 } : 1'b0;
  assign N312 = N29574;
  assign { N29674, N29673, N29672, N29671 } = (N313)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29670)? { N29346, N29347, N29348, N29349 } : 1'b0;
  assign N313 = N29575;
  assign { N29679, N29678, N29677, N29676 } = (N314)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29675)? { N29350, N29351, N29352, N29353 } : 1'b0;
  assign N314 = N29576;
  assign { N29684, N29683, N29682, N29681 } = (N315)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29680)? { N29354, N29355, N29356, N29357 } : 1'b0;
  assign N315 = N29577;
  assign { N29689, N29688, N29687, N29686 } = (N316)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29685)? { N29358, N29359, N29360, N29361 } : 1'b0;
  assign N316 = N29578;
  assign { N29694, N29693, N29692, N29691 } = (N317)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29690)? { N29362, N29363, N29364, N29365 } : 1'b0;
  assign N317 = N29579;
  assign { N29699, N29698, N29697, N29696 } = (N318)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29695)? { N29366, N29367, N29368, N29369 } : 1'b0;
  assign N318 = N29580;
  assign { N29704, N29703, N29702, N29701 } = (N319)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29700)? { N29370, N29371, N29372, N29373 } : 1'b0;
  assign N319 = N29581;
  assign { N29709, N29708, N29707, N29706 } = (N320)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29705)? { N29374, N29375, N29376, N29377 } : 1'b0;
  assign N320 = N29582;
  assign { N29714, N29713, N29712, N29711 } = (N321)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29710)? { N29378, N29379, N29380, N29381 } : 1'b0;
  assign N321 = N29583;
  assign { N29719, N29718, N29717, N29716 } = (N322)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29715)? { N29382, N29383, N29384, N29385 } : 1'b0;
  assign N322 = N29584;
  assign { N29724, N29723, N29722, N29721 } = (N323)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29720)? { N29386, N29387, N29388, N29389 } : 1'b0;
  assign N323 = N29585;
  assign { N29729, N29728, N29727, N29726 } = (N324)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29725)? { N29390, N29391, N29392, N29393 } : 1'b0;
  assign N324 = N29586;
  assign { N29734, N29733, N29732, N29731 } = (N325)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29730)? { N29394, N29395, N29396, N29397 } : 1'b0;
  assign N325 = N29587;
  assign { N29739, N29738, N29737, N29736 } = (N326)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29735)? { N29398, N29399, N29400, N29401 } : 1'b0;
  assign N326 = N29588;
  assign { N29744, N29743, N29742, N29741 } = (N327)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29740)? { N29402, N29403, N29404, N29405 } : 1'b0;
  assign N327 = N29589;
  assign { N29749, N29748, N29747, N29746 } = (N328)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29745)? { N29406, N29407, N29408, N29409 } : 1'b0;
  assign N328 = N29590;
  assign { N29754, N29753, N29752, N29751 } = (N329)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29750)? { N29410, N29411, N29412, N29413 } : 1'b0;
  assign N329 = N29591;
  assign { N29759, N29758, N29757, N29756 } = (N330)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29755)? { N29414, N29415, N29416, N29417 } : 1'b0;
  assign N330 = N29592;
  assign { N29764, N29763, N29762, N29761 } = (N331)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29760)? { N29418, N29419, N29420, N29421 } : 1'b0;
  assign N331 = N29593;
  assign { N29769, N29768, N29767, N29766 } = (N332)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29765)? { N29422, N29423, N29424, N29425 } : 1'b0;
  assign N332 = N29594;
  assign { N29774, N29773, N29772, N29771 } = (N333)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29770)? { N29426, N29427, N29428, N29429 } : 1'b0;
  assign N333 = N29595;
  assign { N29779, N29778, N29777, N29776 } = (N334)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29775)? { N29430, N29431, N29432, N29433 } : 1'b0;
  assign N334 = N29596;
  assign { N29784, N29783, N29782, N29781 } = (N335)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29780)? { N29434, N29435, N29436, N29437 } : 1'b0;
  assign N335 = N29597;
  assign { N29789, N29788, N29787, N29786 } = (N336)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29785)? { N29438, N29439, N29440, N29441 } : 1'b0;
  assign N336 = N29598;
  assign { N29794, N29793, N29792, N29791 } = (N337)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29790)? { N29442, N29443, N29444, N29445 } : 1'b0;
  assign N337 = N29599;
  assign { N29799, N29798, N29797, N29796 } = (N338)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29795)? { N29446, N29447, N29448, N29449 } : 1'b0;
  assign N338 = N29600;
  assign { N29804, N29803, N29802, N29801 } = (N339)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29800)? { N29450, N29451, N29452, N29453 } : 1'b0;
  assign N339 = N29601;
  assign { N29809, N29808, N29807, N29806 } = (N340)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29805)? { N29454, N29455, N29456, N29457 } : 1'b0;
  assign N340 = N29602;
  assign { N29814, N29813, N29812, N29811 } = (N341)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29810)? { N29458, N29459, N29460, N29461 } : 1'b0;
  assign N341 = N29603;
  assign { N29819, N29818, N29817, N29816 } = (N342)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29815)? { N29462, N29463, N29464, N29465 } : 1'b0;
  assign N342 = N29604;
  assign { N29824, N29823, N29822, N29821 } = (N343)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29820)? { N29466, N29467, N29468, N29469 } : 1'b0;
  assign N343 = N29605;
  assign { N29829, N29828, N29827, N29826 } = (N344)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29825)? { N29470, N29471, N29472, N29473 } : 1'b0;
  assign N344 = N29606;
  assign { N29834, N29833, N29832, N29831 } = (N345)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29830)? { N29474, N29475, N29476, N29477 } : 1'b0;
  assign N345 = N29607;
  assign { N29839, N29838, N29837, N29836 } = (N346)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29835)? { N29478, N29479, N29480, N29481 } : 1'b0;
  assign N346 = N29608;
  assign { N29844, N29843, N29842, N29841 } = (N347)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29840)? { N29482, N29483, N29484, N29485 } : 1'b0;
  assign N347 = N29609;
  assign { N29849, N29848, N29847, N29846 } = (N348)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29845)? { N29486, N29487, N29488, N29489 } : 1'b0;
  assign N348 = N29610;
  assign { N29854, N29853, N29852, N29851 } = (N349)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29850)? { N29490, N29491, N29492, N29493 } : 1'b0;
  assign N349 = N29611;
  assign { N29859, N29858, N29857, N29856 } = (N350)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29855)? { N29494, N29495, N29496, N29497 } : 1'b0;
  assign N350 = N29612;
  assign { N29864, N29863, N29862, N29861 } = (N351)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29860)? { N29498, N29499, N29500, N29501 } : 1'b0;
  assign N351 = N29613;
  assign { N29869, N29868, N29867, N29866 } = (N352)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29865)? { N29502, N29503, N29504, N29505 } : 1'b0;
  assign N352 = N29614;
  assign { N29874, N29873, N29872, N29871 } = (N353)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29870)? { N29506, N29507, N29508, N29509 } : 1'b0;
  assign N353 = N29615;
  assign { N29879, N29878, N29877, N29876 } = (N354)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29875)? { N29510, N29511, N29512, N29513 } : 1'b0;
  assign N354 = N29616;
  assign { N29884, N29883, N29882, N29881 } = (N355)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29880)? { N29514, N29515, N29516, N29517 } : 1'b0;
  assign N355 = N29617;
  assign { N29889, N29888, N29887, N29886 } = (N356)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29885)? { N29518, N29519, N29520, N29521 } : 1'b0;
  assign N356 = N29618;
  assign { N29894, N29893, N29892, N29891 } = (N357)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29890)? { N29522, N29523, N29524, N29525 } : 1'b0;
  assign N357 = N29619;
  assign { N29899, N29898, N29897, N29896 } = (N358)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29895)? { N29526, N29527, N29528, N29529 } : 1'b0;
  assign N358 = N29620;
  assign { N29904, N29903, N29902, N29901 } = (N359)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29900)? { N29530, N29531, N29532, N29533 } : 1'b0;
  assign N359 = N29621;
  assign { N29909, N29908, N29907, N29906 } = (N360)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29905)? { N29534, N29535, N29536, N29537 } : 1'b0;
  assign N360 = N29622;
  assign { N29914, N29913, N29912, N29911 } = (N361)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29910)? { N29538, N29539, N29540, N29541 } : 1'b0;
  assign N361 = N29623;
  assign { N29919, N29918, N29917, N29916 } = (N362)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29915)? { N29542, N29543, N29544, N29545 } : 1'b0;
  assign N362 = N29624;
  assign { N29924, N29923, N29922, N29921 } = (N363)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29920)? { N29546, N29547, N29548, N29549 } : 1'b0;
  assign N363 = N29625;
  assign { N29929, N29928, N29927, N29926 } = (N364)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29925)? { N29550, N29551, N29552, N29553 } : 1'b0;
  assign N364 = N29626;
  assign { N29934, N29933, N29932, N29931 } = (N365)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29930)? { N29554, N29555, N29556, N29557 } : 1'b0;
  assign N365 = N29627;
  assign { N29939, N29938, N29937, N29936 } = (N366)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29935)? { N29558, N29559, N29560, N29561 } : 1'b0;
  assign N366 = N29628;
  assign { N29944, N29943, N29942, N29941 } = (N367)? { mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657] } : 
                                              (N29940)? { N29562, N29563, N29564, N29565 } : 1'b0;
  assign N367 = N29629;
  assign { N30196, N30195, N30194, N30193, N30192, N30191, N30190, N30189, N30188, N30187, N30186, N30185, N30184, N30183, N30182, N30181, N30180, N30179, N30178, N30177, N30176, N30175, N30174, N30173, N30172, N30171, N30170, N30169, N30168, N30167, N30166, N30165, N30164, N30163, N30162, N30161, N30160, N30159, N30158, N30157, N30156, N30155, N30154, N30153, N30152, N30151, N30150, N30149, N30148, N30147, N30146, N30145, N30144, N30143, N30142, N30141, N30140, N30139, N30138, N30137, N30136, N30135, N30134, N30133, N30132, N30131, N30130, N30129, N30128, N30127, N30126, N30125, N30124, N30123, N30122, N30121, N30120, N30119, N30118, N30117, N30116, N30115, N30114, N30113, N30112, N30111, N30110, N30109, N30108, N30107, N30106, N30105, N30104, N30103, N30102, N30101, N30100, N30099, N30098, N30097, N30096, N30095, N30094, N30093, N30092, N30091, N30090, N30089, N30088, N30087, N30086, N30085, N30084, N30083, N30082, N30081, N30080, N30079, N30078, N30077, N30076, N30075, N30074, N30073, N30072, N30071, N30070, N30069, N30068, N30067, N30066, N30065, N30064, N30063, N30062, N30061, N30060, N30059, N30058, N30057, N30056, N30055, N30054, N30053, N30052, N30051, N30050, N30049, N30048, N30047, N30046, N30045, N30044, N30043, N30042, N30041, N30040, N30039, N30038, N30037, N30036, N30035, N30034, N30033, N30032, N30031, N30030, N30029, N30028, N30027, N30026, N30025, N30024, N30023, N30022, N30021, N30020, N30019, N30018, N30017, N30016, N30015, N30014, N30013, N30012, N30011, N30010, N30009, N30008, N30007, N30006, N30005, N30004, N30003, N30002, N30001, N30000, N29999, N29998, N29997, N29996, N29995, N29994, N29993, N29992, N29991, N29990, N29989, N29988, N29987, N29986, N29985, N29984, N29983, N29982, N29981, N29980, N29979, N29978, N29977, N29976, N29975, N29974, N29973, N29972, N29971, N29970, N29969, N29968, N29967, N29966, N29965, N29964, N29963, N29962, N29961, N29960, N29959, N29958, N29957, N29956, N29955, N29954, N29953, N29952, N29951, N29950, N29949, N29948, N29947, N29946, N29945 } = (N368)? { N29941, N29942, N29943, N29944, N29936, N29937, N29938, N29939, N29931, N29932, N29933, N29934, N29926, N29927, N29928, N29929, N29921, N29922, N29923, N29924, N29916, N29917, N29918, N29919, N29911, N29912, N29913, N29914, N29906, N29907, N29908, N29909, N29901, N29902, N29903, N29904, N29896, N29897, N29898, N29899, N29891, N29892, N29893, N29894, N29886, N29887, N29888, N29889, N29881, N29882, N29883, N29884, N29876, N29877, N29878, N29879, N29871, N29872, N29873, N29874, N29866, N29867, N29868, N29869, N29861, N29862, N29863, N29864, N29856, N29857, N29858, N29859, N29851, N29852, N29853, N29854, N29846, N29847, N29848, N29849, N29841, N29842, N29843, N29844, N29836, N29837, N29838, N29839, N29831, N29832, N29833, N29834, N29826, N29827, N29828, N29829, N29821, N29822, N29823, N29824, N29816, N29817, N29818, N29819, N29811, N29812, N29813, N29814, N29806, N29807, N29808, N29809, N29801, N29802, N29803, N29804, N29796, N29797, N29798, N29799, N29791, N29792, N29793, N29794, N29786, N29787, N29788, N29789, N29781, N29782, N29783, N29784, N29776, N29777, N29778, N29779, N29771, N29772, N29773, N29774, N29766, N29767, N29768, N29769, N29761, N29762, N29763, N29764, N29756, N29757, N29758, N29759, N29751, N29752, N29753, N29754, N29746, N29747, N29748, N29749, N29741, N29742, N29743, N29744, N29736, N29737, N29738, N29739, N29731, N29732, N29733, N29734, N29726, N29727, N29728, N29729, N29721, N29722, N29723, N29724, N29716, N29717, N29718, N29719, N29711, N29712, N29713, N29714, N29706, N29707, N29708, N29709, N29701, N29702, N29703, N29704, N29696, N29697, N29698, N29699, N29691, N29692, N29693, N29694, N29686, N29687, N29688, N29689, N29681, N29682, N29683, N29684, N29676, N29677, N29678, N29679, N29671, N29672, N29673, N29674, N29666, N29667, N29668, N29669, N29661, N29662, N29663, N29664, N29656, N29657, N29658, N29659, N29651, N29652, N29653, N29654, N29646, N29647, N29648, N29649, N29641, N29642, N29643, N29644, N29636, N29637, N29638, N29639, N29631, N29632, N29633, N29634 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N29566)? { N29565, N29564, N29563, N29562, N29561, N29560, N29559, N29558, N29557, N29556, N29555, N29554, N29553, N29552, N29551, N29550, N29549, N29548, N29547, N29546, N29545, N29544, N29543, N29542, N29541, N29540, N29539, N29538, N29537, N29536, N29535, N29534, N29533, N29532, N29531, N29530, N29529, N29528, N29527, N29526, N29525, N29524, N29523, N29522, N29521, N29520, N29519, N29518, N29517, N29516, N29515, N29514, N29513, N29512, N29511, N29510, N29509, N29508, N29507, N29506, N29505, N29504, N29503, N29502, N29501, N29500, N29499, N29498, N29497, N29496, N29495, N29494, N29493, N29492, N29491, N29490, N29489, N29488, N29487, N29486, N29485, N29484, N29483, N29482, N29481, N29480, N29479, N29478, N29477, N29476, N29475, N29474, N29473, N29472, N29471, N29470, N29469, N29468, N29467, N29466, N29465, N29464, N29463, N29462, N29461, N29460, N29459, N29458, N29457, N29456, N29455, N29454, N29453, N29452, N29451, N29450, N29449, N29448, N29447, N29446, N29445, N29444, N29443, N29442, N29441, N29440, N29439, N29438, N29437, N29436, N29435, N29434, N29433, N29432, N29431, N29430, N29429, N29428, N29427, N29426, N29425, N29424, N29423, N29422, N29421, N29420, N29419, N29418, N29417, N29416, N29415, N29414, N29413, N29412, N29411, N29410, N29409, N29408, N29407, N29406, N29405, N29404, N29403, N29402, N29401, N29400, N29399, N29398, N29397, N29396, N29395, N29394, N29393, N29392, N29391, N29390, N29389, N29388, N29387, N29386, N29385, N29384, N29383, N29382, N29381, N29380, N29379, N29378, N29377, N29376, N29375, N29374, N29373, N29372, N29371, N29370, N29369, N29368, N29367, N29366, N29365, N29364, N29363, N29362, N29361, N29360, N29359, N29358, N29357, N29356, N29355, N29354, N29353, N29352, N29351, N29350, N29349, N29348, N29347, N29346, N29345, N29344, N29343, N29342, N29341, N29340, N29339, N29338, N29337, N29336, N29335, N29334, N29333, N29332, N29331, N29330, N29329, N29328, N29327, N29326, N29325, N29324, N29323, N29322, N29321, N29320, N29319, N29318, N29317, N29316, N29315, N29314 } : 1'b0;
  assign N368 = mem_q[725];
  assign { N30265, N30264, N30263, N30262 } = (N369)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30261)? { N29945, N29946, N29947, N29948 } : 1'b0;
  assign N369 = N30198;
  assign { N30270, N30269, N30268, N30267 } = (N370)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30266)? { N29949, N29950, N29951, N29952 } : 1'b0;
  assign N370 = N30199;
  assign { N30275, N30274, N30273, N30272 } = (N371)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30271)? { N29953, N29954, N29955, N29956 } : 1'b0;
  assign N371 = N30200;
  assign { N30280, N30279, N30278, N30277 } = (N372)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30276)? { N29957, N29958, N29959, N29960 } : 1'b0;
  assign N372 = N30201;
  assign { N30285, N30284, N30283, N30282 } = (N373)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30281)? { N29961, N29962, N29963, N29964 } : 1'b0;
  assign N373 = N30202;
  assign { N30290, N30289, N30288, N30287 } = (N374)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30286)? { N29965, N29966, N29967, N29968 } : 1'b0;
  assign N374 = N30203;
  assign { N30295, N30294, N30293, N30292 } = (N375)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30291)? { N29969, N29970, N29971, N29972 } : 1'b0;
  assign N375 = N30204;
  assign { N30300, N30299, N30298, N30297 } = (N376)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30296)? { N29973, N29974, N29975, N29976 } : 1'b0;
  assign N376 = N30205;
  assign { N30305, N30304, N30303, N30302 } = (N377)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30301)? { N29977, N29978, N29979, N29980 } : 1'b0;
  assign N377 = N30206;
  assign { N30310, N30309, N30308, N30307 } = (N378)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30306)? { N29981, N29982, N29983, N29984 } : 1'b0;
  assign N378 = N30207;
  assign { N30315, N30314, N30313, N30312 } = (N379)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30311)? { N29985, N29986, N29987, N29988 } : 1'b0;
  assign N379 = N30208;
  assign { N30320, N30319, N30318, N30317 } = (N380)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30316)? { N29989, N29990, N29991, N29992 } : 1'b0;
  assign N380 = N30209;
  assign { N30325, N30324, N30323, N30322 } = (N381)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30321)? { N29993, N29994, N29995, N29996 } : 1'b0;
  assign N381 = N30210;
  assign { N30330, N30329, N30328, N30327 } = (N382)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30326)? { N29997, N29998, N29999, N30000 } : 1'b0;
  assign N382 = N30211;
  assign { N30335, N30334, N30333, N30332 } = (N383)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30331)? { N30001, N30002, N30003, N30004 } : 1'b0;
  assign N383 = N30212;
  assign { N30340, N30339, N30338, N30337 } = (N384)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30336)? { N30005, N30006, N30007, N30008 } : 1'b0;
  assign N384 = N30213;
  assign { N30345, N30344, N30343, N30342 } = (N385)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30341)? { N30009, N30010, N30011, N30012 } : 1'b0;
  assign N385 = N30214;
  assign { N30350, N30349, N30348, N30347 } = (N386)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30346)? { N30013, N30014, N30015, N30016 } : 1'b0;
  assign N386 = N30215;
  assign { N30355, N30354, N30353, N30352 } = (N387)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30351)? { N30017, N30018, N30019, N30020 } : 1'b0;
  assign N387 = N30216;
  assign { N30360, N30359, N30358, N30357 } = (N388)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30356)? { N30021, N30022, N30023, N30024 } : 1'b0;
  assign N388 = N30217;
  assign { N30365, N30364, N30363, N30362 } = (N389)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30361)? { N30025, N30026, N30027, N30028 } : 1'b0;
  assign N389 = N30218;
  assign { N30370, N30369, N30368, N30367 } = (N390)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30366)? { N30029, N30030, N30031, N30032 } : 1'b0;
  assign N390 = N30219;
  assign { N30375, N30374, N30373, N30372 } = (N391)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30371)? { N30033, N30034, N30035, N30036 } : 1'b0;
  assign N391 = N30220;
  assign { N30380, N30379, N30378, N30377 } = (N392)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30376)? { N30037, N30038, N30039, N30040 } : 1'b0;
  assign N392 = N30221;
  assign { N30385, N30384, N30383, N30382 } = (N393)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30381)? { N30041, N30042, N30043, N30044 } : 1'b0;
  assign N393 = N30222;
  assign { N30390, N30389, N30388, N30387 } = (N394)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30386)? { N30045, N30046, N30047, N30048 } : 1'b0;
  assign N394 = N30223;
  assign { N30395, N30394, N30393, N30392 } = (N395)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30391)? { N30049, N30050, N30051, N30052 } : 1'b0;
  assign N395 = N30224;
  assign { N30400, N30399, N30398, N30397 } = (N396)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30396)? { N30053, N30054, N30055, N30056 } : 1'b0;
  assign N396 = N30225;
  assign { N30405, N30404, N30403, N30402 } = (N397)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30401)? { N30057, N30058, N30059, N30060 } : 1'b0;
  assign N397 = N30226;
  assign { N30410, N30409, N30408, N30407 } = (N398)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30406)? { N30061, N30062, N30063, N30064 } : 1'b0;
  assign N398 = N30227;
  assign { N30415, N30414, N30413, N30412 } = (N399)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30411)? { N30065, N30066, N30067, N30068 } : 1'b0;
  assign N399 = N30228;
  assign { N30420, N30419, N30418, N30417 } = (N400)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30416)? { N30069, N30070, N30071, N30072 } : 1'b0;
  assign N400 = N30229;
  assign { N30425, N30424, N30423, N30422 } = (N401)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30421)? { N30073, N30074, N30075, N30076 } : 1'b0;
  assign N401 = N30230;
  assign { N30430, N30429, N30428, N30427 } = (N402)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30426)? { N30077, N30078, N30079, N30080 } : 1'b0;
  assign N402 = N30231;
  assign { N30435, N30434, N30433, N30432 } = (N403)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30431)? { N30081, N30082, N30083, N30084 } : 1'b0;
  assign N403 = N30232;
  assign { N30440, N30439, N30438, N30437 } = (N404)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30436)? { N30085, N30086, N30087, N30088 } : 1'b0;
  assign N404 = N30233;
  assign { N30445, N30444, N30443, N30442 } = (N405)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30441)? { N30089, N30090, N30091, N30092 } : 1'b0;
  assign N405 = N30234;
  assign { N30450, N30449, N30448, N30447 } = (N406)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30446)? { N30093, N30094, N30095, N30096 } : 1'b0;
  assign N406 = N30235;
  assign { N30455, N30454, N30453, N30452 } = (N407)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30451)? { N30097, N30098, N30099, N30100 } : 1'b0;
  assign N407 = N30236;
  assign { N30460, N30459, N30458, N30457 } = (N408)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30456)? { N30101, N30102, N30103, N30104 } : 1'b0;
  assign N408 = N30237;
  assign { N30465, N30464, N30463, N30462 } = (N409)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30461)? { N30105, N30106, N30107, N30108 } : 1'b0;
  assign N409 = N30238;
  assign { N30470, N30469, N30468, N30467 } = (N410)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30466)? { N30109, N30110, N30111, N30112 } : 1'b0;
  assign N410 = N30239;
  assign { N30475, N30474, N30473, N30472 } = (N411)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30471)? { N30113, N30114, N30115, N30116 } : 1'b0;
  assign N411 = N30240;
  assign { N30480, N30479, N30478, N30477 } = (N412)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30476)? { N30117, N30118, N30119, N30120 } : 1'b0;
  assign N412 = N30241;
  assign { N30485, N30484, N30483, N30482 } = (N413)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30481)? { N30121, N30122, N30123, N30124 } : 1'b0;
  assign N413 = N30242;
  assign { N30490, N30489, N30488, N30487 } = (N414)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30486)? { N30125, N30126, N30127, N30128 } : 1'b0;
  assign N414 = N30243;
  assign { N30495, N30494, N30493, N30492 } = (N415)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30491)? { N30129, N30130, N30131, N30132 } : 1'b0;
  assign N415 = N30244;
  assign { N30500, N30499, N30498, N30497 } = (N416)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30496)? { N30133, N30134, N30135, N30136 } : 1'b0;
  assign N416 = N30245;
  assign { N30505, N30504, N30503, N30502 } = (N417)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30501)? { N30137, N30138, N30139, N30140 } : 1'b0;
  assign N417 = N30246;
  assign { N30510, N30509, N30508, N30507 } = (N418)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30506)? { N30141, N30142, N30143, N30144 } : 1'b0;
  assign N418 = N30247;
  assign { N30515, N30514, N30513, N30512 } = (N419)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30511)? { N30145, N30146, N30147, N30148 } : 1'b0;
  assign N419 = N30248;
  assign { N30520, N30519, N30518, N30517 } = (N420)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30516)? { N30149, N30150, N30151, N30152 } : 1'b0;
  assign N420 = N30249;
  assign { N30525, N30524, N30523, N30522 } = (N421)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30521)? { N30153, N30154, N30155, N30156 } : 1'b0;
  assign N421 = N30250;
  assign { N30530, N30529, N30528, N30527 } = (N422)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30526)? { N30157, N30158, N30159, N30160 } : 1'b0;
  assign N422 = N30251;
  assign { N30535, N30534, N30533, N30532 } = (N423)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30531)? { N30161, N30162, N30163, N30164 } : 1'b0;
  assign N423 = N30252;
  assign { N30540, N30539, N30538, N30537 } = (N424)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30536)? { N30165, N30166, N30167, N30168 } : 1'b0;
  assign N424 = N30253;
  assign { N30545, N30544, N30543, N30542 } = (N425)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30541)? { N30169, N30170, N30171, N30172 } : 1'b0;
  assign N425 = N30254;
  assign { N30550, N30549, N30548, N30547 } = (N426)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30546)? { N30173, N30174, N30175, N30176 } : 1'b0;
  assign N426 = N30255;
  assign { N30555, N30554, N30553, N30552 } = (N427)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30551)? { N30177, N30178, N30179, N30180 } : 1'b0;
  assign N427 = N30256;
  assign { N30560, N30559, N30558, N30557 } = (N428)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30556)? { N30181, N30182, N30183, N30184 } : 1'b0;
  assign N428 = N30257;
  assign { N30565, N30564, N30563, N30562 } = (N429)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30561)? { N30185, N30186, N30187, N30188 } : 1'b0;
  assign N429 = N30258;
  assign { N30570, N30569, N30568, N30567 } = (N430)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30566)? { N30189, N30190, N30191, N30192 } : 1'b0;
  assign N430 = N30259;
  assign { N30575, N30574, N30573, N30572 } = (N431)? { mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020] } : 
                                              (N30571)? { N30193, N30194, N30195, N30196 } : 1'b0;
  assign N431 = N30260;
  assign { N30827, N30826, N30825, N30824, N30823, N30822, N30821, N30820, N30819, N30818, N30817, N30816, N30815, N30814, N30813, N30812, N30811, N30810, N30809, N30808, N30807, N30806, N30805, N30804, N30803, N30802, N30801, N30800, N30799, N30798, N30797, N30796, N30795, N30794, N30793, N30792, N30791, N30790, N30789, N30788, N30787, N30786, N30785, N30784, N30783, N30782, N30781, N30780, N30779, N30778, N30777, N30776, N30775, N30774, N30773, N30772, N30771, N30770, N30769, N30768, N30767, N30766, N30765, N30764, N30763, N30762, N30761, N30760, N30759, N30758, N30757, N30756, N30755, N30754, N30753, N30752, N30751, N30750, N30749, N30748, N30747, N30746, N30745, N30744, N30743, N30742, N30741, N30740, N30739, N30738, N30737, N30736, N30735, N30734, N30733, N30732, N30731, N30730, N30729, N30728, N30727, N30726, N30725, N30724, N30723, N30722, N30721, N30720, N30719, N30718, N30717, N30716, N30715, N30714, N30713, N30712, N30711, N30710, N30709, N30708, N30707, N30706, N30705, N30704, N30703, N30702, N30701, N30700, N30699, N30698, N30697, N30696, N30695, N30694, N30693, N30692, N30691, N30690, N30689, N30688, N30687, N30686, N30685, N30684, N30683, N30682, N30681, N30680, N30679, N30678, N30677, N30676, N30675, N30674, N30673, N30672, N30671, N30670, N30669, N30668, N30667, N30666, N30665, N30664, N30663, N30662, N30661, N30660, N30659, N30658, N30657, N30656, N30655, N30654, N30653, N30652, N30651, N30650, N30649, N30648, N30647, N30646, N30645, N30644, N30643, N30642, N30641, N30640, N30639, N30638, N30637, N30636, N30635, N30634, N30633, N30632, N30631, N30630, N30629, N30628, N30627, N30626, N30625, N30624, N30623, N30622, N30621, N30620, N30619, N30618, N30617, N30616, N30615, N30614, N30613, N30612, N30611, N30610, N30609, N30608, N30607, N30606, N30605, N30604, N30603, N30602, N30601, N30600, N30599, N30598, N30597, N30596, N30595, N30594, N30593, N30592, N30591, N30590, N30589, N30588, N30587, N30586, N30585, N30584, N30583, N30582, N30581, N30580, N30579, N30578, N30577, N30576 } = (N432)? { N30572, N30573, N30574, N30575, N30567, N30568, N30569, N30570, N30562, N30563, N30564, N30565, N30557, N30558, N30559, N30560, N30552, N30553, N30554, N30555, N30547, N30548, N30549, N30550, N30542, N30543, N30544, N30545, N30537, N30538, N30539, N30540, N30532, N30533, N30534, N30535, N30527, N30528, N30529, N30530, N30522, N30523, N30524, N30525, N30517, N30518, N30519, N30520, N30512, N30513, N30514, N30515, N30507, N30508, N30509, N30510, N30502, N30503, N30504, N30505, N30497, N30498, N30499, N30500, N30492, N30493, N30494, N30495, N30487, N30488, N30489, N30490, N30482, N30483, N30484, N30485, N30477, N30478, N30479, N30480, N30472, N30473, N30474, N30475, N30467, N30468, N30469, N30470, N30462, N30463, N30464, N30465, N30457, N30458, N30459, N30460, N30452, N30453, N30454, N30455, N30447, N30448, N30449, N30450, N30442, N30443, N30444, N30445, N30437, N30438, N30439, N30440, N30432, N30433, N30434, N30435, N30427, N30428, N30429, N30430, N30422, N30423, N30424, N30425, N30417, N30418, N30419, N30420, N30412, N30413, N30414, N30415, N30407, N30408, N30409, N30410, N30402, N30403, N30404, N30405, N30397, N30398, N30399, N30400, N30392, N30393, N30394, N30395, N30387, N30388, N30389, N30390, N30382, N30383, N30384, N30385, N30377, N30378, N30379, N30380, N30372, N30373, N30374, N30375, N30367, N30368, N30369, N30370, N30362, N30363, N30364, N30365, N30357, N30358, N30359, N30360, N30352, N30353, N30354, N30355, N30347, N30348, N30349, N30350, N30342, N30343, N30344, N30345, N30337, N30338, N30339, N30340, N30332, N30333, N30334, N30335, N30327, N30328, N30329, N30330, N30322, N30323, N30324, N30325, N30317, N30318, N30319, N30320, N30312, N30313, N30314, N30315, N30307, N30308, N30309, N30310, N30302, N30303, N30304, N30305, N30297, N30298, N30299, N30300, N30292, N30293, N30294, N30295, N30287, N30288, N30289, N30290, N30282, N30283, N30284, N30285, N30277, N30278, N30279, N30280, N30272, N30273, N30274, N30275, N30267, N30268, N30269, N30270, N30262, N30263, N30264, N30265 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N30197)? { N30196, N30195, N30194, N30193, N30192, N30191, N30190, N30189, N30188, N30187, N30186, N30185, N30184, N30183, N30182, N30181, N30180, N30179, N30178, N30177, N30176, N30175, N30174, N30173, N30172, N30171, N30170, N30169, N30168, N30167, N30166, N30165, N30164, N30163, N30162, N30161, N30160, N30159, N30158, N30157, N30156, N30155, N30154, N30153, N30152, N30151, N30150, N30149, N30148, N30147, N30146, N30145, N30144, N30143, N30142, N30141, N30140, N30139, N30138, N30137, N30136, N30135, N30134, N30133, N30132, N30131, N30130, N30129, N30128, N30127, N30126, N30125, N30124, N30123, N30122, N30121, N30120, N30119, N30118, N30117, N30116, N30115, N30114, N30113, N30112, N30111, N30110, N30109, N30108, N30107, N30106, N30105, N30104, N30103, N30102, N30101, N30100, N30099, N30098, N30097, N30096, N30095, N30094, N30093, N30092, N30091, N30090, N30089, N30088, N30087, N30086, N30085, N30084, N30083, N30082, N30081, N30080, N30079, N30078, N30077, N30076, N30075, N30074, N30073, N30072, N30071, N30070, N30069, N30068, N30067, N30066, N30065, N30064, N30063, N30062, N30061, N30060, N30059, N30058, N30057, N30056, N30055, N30054, N30053, N30052, N30051, N30050, N30049, N30048, N30047, N30046, N30045, N30044, N30043, N30042, N30041, N30040, N30039, N30038, N30037, N30036, N30035, N30034, N30033, N30032, N30031, N30030, N30029, N30028, N30027, N30026, N30025, N30024, N30023, N30022, N30021, N30020, N30019, N30018, N30017, N30016, N30015, N30014, N30013, N30012, N30011, N30010, N30009, N30008, N30007, N30006, N30005, N30004, N30003, N30002, N30001, N30000, N29999, N29998, N29997, N29996, N29995, N29994, N29993, N29992, N29991, N29990, N29989, N29988, N29987, N29986, N29985, N29984, N29983, N29982, N29981, N29980, N29979, N29978, N29977, N29976, N29975, N29974, N29973, N29972, N29971, N29970, N29969, N29968, N29967, N29966, N29965, N29964, N29963, N29962, N29961, N29960, N29959, N29958, N29957, N29956, N29955, N29954, N29953, N29952, N29951, N29950, N29949, N29948, N29947, N29946, N29945 } : 1'b0;
  assign N432 = mem_q[1088];
  assign { N30896, N30895, N30894, N30893 } = (N433)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30892)? { N30576, N30577, N30578, N30579 } : 1'b0;
  assign N433 = N30829;
  assign { N30901, N30900, N30899, N30898 } = (N434)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30897)? { N30580, N30581, N30582, N30583 } : 1'b0;
  assign N434 = N30830;
  assign { N30906, N30905, N30904, N30903 } = (N435)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30902)? { N30584, N30585, N30586, N30587 } : 1'b0;
  assign N435 = N30831;
  assign { N30911, N30910, N30909, N30908 } = (N436)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30907)? { N30588, N30589, N30590, N30591 } : 1'b0;
  assign N436 = N30832;
  assign { N30916, N30915, N30914, N30913 } = (N437)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30912)? { N30592, N30593, N30594, N30595 } : 1'b0;
  assign N437 = N30833;
  assign { N30921, N30920, N30919, N30918 } = (N438)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30917)? { N30596, N30597, N30598, N30599 } : 1'b0;
  assign N438 = N30834;
  assign { N30926, N30925, N30924, N30923 } = (N439)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30922)? { N30600, N30601, N30602, N30603 } : 1'b0;
  assign N439 = N30835;
  assign { N30931, N30930, N30929, N30928 } = (N440)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30927)? { N30604, N30605, N30606, N30607 } : 1'b0;
  assign N440 = N30836;
  assign { N30936, N30935, N30934, N30933 } = (N441)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30932)? { N30608, N30609, N30610, N30611 } : 1'b0;
  assign N441 = N30837;
  assign { N30941, N30940, N30939, N30938 } = (N442)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30937)? { N30612, N30613, N30614, N30615 } : 1'b0;
  assign N442 = N30838;
  assign { N30946, N30945, N30944, N30943 } = (N443)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30942)? { N30616, N30617, N30618, N30619 } : 1'b0;
  assign N443 = N30839;
  assign { N30951, N30950, N30949, N30948 } = (N444)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30947)? { N30620, N30621, N30622, N30623 } : 1'b0;
  assign N444 = N30840;
  assign { N30956, N30955, N30954, N30953 } = (N445)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30952)? { N30624, N30625, N30626, N30627 } : 1'b0;
  assign N445 = N30841;
  assign { N30961, N30960, N30959, N30958 } = (N446)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30957)? { N30628, N30629, N30630, N30631 } : 1'b0;
  assign N446 = N30842;
  assign { N30966, N30965, N30964, N30963 } = (N447)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30962)? { N30632, N30633, N30634, N30635 } : 1'b0;
  assign N447 = N30843;
  assign { N30971, N30970, N30969, N30968 } = (N448)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30967)? { N30636, N30637, N30638, N30639 } : 1'b0;
  assign N448 = N30844;
  assign { N30976, N30975, N30974, N30973 } = (N449)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30972)? { N30640, N30641, N30642, N30643 } : 1'b0;
  assign N449 = N30845;
  assign { N30981, N30980, N30979, N30978 } = (N450)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30977)? { N30644, N30645, N30646, N30647 } : 1'b0;
  assign N450 = N30846;
  assign { N30986, N30985, N30984, N30983 } = (N451)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30982)? { N30648, N30649, N30650, N30651 } : 1'b0;
  assign N451 = N30847;
  assign { N30991, N30990, N30989, N30988 } = (N452)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30987)? { N30652, N30653, N30654, N30655 } : 1'b0;
  assign N452 = N30848;
  assign { N30996, N30995, N30994, N30993 } = (N453)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30992)? { N30656, N30657, N30658, N30659 } : 1'b0;
  assign N453 = N30849;
  assign { N31001, N31000, N30999, N30998 } = (N454)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N30997)? { N30660, N30661, N30662, N30663 } : 1'b0;
  assign N454 = N30850;
  assign { N31006, N31005, N31004, N31003 } = (N455)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31002)? { N30664, N30665, N30666, N30667 } : 1'b0;
  assign N455 = N30851;
  assign { N31011, N31010, N31009, N31008 } = (N456)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31007)? { N30668, N30669, N30670, N30671 } : 1'b0;
  assign N456 = N30852;
  assign { N31016, N31015, N31014, N31013 } = (N457)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31012)? { N30672, N30673, N30674, N30675 } : 1'b0;
  assign N457 = N30853;
  assign { N31021, N31020, N31019, N31018 } = (N458)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31017)? { N30676, N30677, N30678, N30679 } : 1'b0;
  assign N458 = N30854;
  assign { N31026, N31025, N31024, N31023 } = (N459)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31022)? { N30680, N30681, N30682, N30683 } : 1'b0;
  assign N459 = N30855;
  assign { N31031, N31030, N31029, N31028 } = (N460)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31027)? { N30684, N30685, N30686, N30687 } : 1'b0;
  assign N460 = N30856;
  assign { N31036, N31035, N31034, N31033 } = (N461)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31032)? { N30688, N30689, N30690, N30691 } : 1'b0;
  assign N461 = N30857;
  assign { N31041, N31040, N31039, N31038 } = (N462)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31037)? { N30692, N30693, N30694, N30695 } : 1'b0;
  assign N462 = N30858;
  assign { N31046, N31045, N31044, N31043 } = (N463)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31042)? { N30696, N30697, N30698, N30699 } : 1'b0;
  assign N463 = N30859;
  assign { N31051, N31050, N31049, N31048 } = (N464)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31047)? { N30700, N30701, N30702, N30703 } : 1'b0;
  assign N464 = N30860;
  assign { N31056, N31055, N31054, N31053 } = (N465)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31052)? { N30704, N30705, N30706, N30707 } : 1'b0;
  assign N465 = N30861;
  assign { N31061, N31060, N31059, N31058 } = (N466)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31057)? { N30708, N30709, N30710, N30711 } : 1'b0;
  assign N466 = N30862;
  assign { N31066, N31065, N31064, N31063 } = (N467)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31062)? { N30712, N30713, N30714, N30715 } : 1'b0;
  assign N467 = N30863;
  assign { N31071, N31070, N31069, N31068 } = (N468)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31067)? { N30716, N30717, N30718, N30719 } : 1'b0;
  assign N468 = N30864;
  assign { N31076, N31075, N31074, N31073 } = (N469)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31072)? { N30720, N30721, N30722, N30723 } : 1'b0;
  assign N469 = N30865;
  assign { N31081, N31080, N31079, N31078 } = (N470)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31077)? { N30724, N30725, N30726, N30727 } : 1'b0;
  assign N470 = N30866;
  assign { N31086, N31085, N31084, N31083 } = (N471)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31082)? { N30728, N30729, N30730, N30731 } : 1'b0;
  assign N471 = N30867;
  assign { N31091, N31090, N31089, N31088 } = (N472)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31087)? { N30732, N30733, N30734, N30735 } : 1'b0;
  assign N472 = N30868;
  assign { N31096, N31095, N31094, N31093 } = (N473)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31092)? { N30736, N30737, N30738, N30739 } : 1'b0;
  assign N473 = N30869;
  assign { N31101, N31100, N31099, N31098 } = (N474)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31097)? { N30740, N30741, N30742, N30743 } : 1'b0;
  assign N474 = N30870;
  assign { N31106, N31105, N31104, N31103 } = (N475)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31102)? { N30744, N30745, N30746, N30747 } : 1'b0;
  assign N475 = N30871;
  assign { N31111, N31110, N31109, N31108 } = (N476)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31107)? { N30748, N30749, N30750, N30751 } : 1'b0;
  assign N476 = N30872;
  assign { N31116, N31115, N31114, N31113 } = (N477)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31112)? { N30752, N30753, N30754, N30755 } : 1'b0;
  assign N477 = N30873;
  assign { N31121, N31120, N31119, N31118 } = (N478)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31117)? { N30756, N30757, N30758, N30759 } : 1'b0;
  assign N478 = N30874;
  assign { N31126, N31125, N31124, N31123 } = (N479)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31122)? { N30760, N30761, N30762, N30763 } : 1'b0;
  assign N479 = N30875;
  assign { N31131, N31130, N31129, N31128 } = (N480)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31127)? { N30764, N30765, N30766, N30767 } : 1'b0;
  assign N480 = N30876;
  assign { N31136, N31135, N31134, N31133 } = (N481)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31132)? { N30768, N30769, N30770, N30771 } : 1'b0;
  assign N481 = N30877;
  assign { N31141, N31140, N31139, N31138 } = (N482)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31137)? { N30772, N30773, N30774, N30775 } : 1'b0;
  assign N482 = N30878;
  assign { N31146, N31145, N31144, N31143 } = (N483)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31142)? { N30776, N30777, N30778, N30779 } : 1'b0;
  assign N483 = N30879;
  assign { N31151, N31150, N31149, N31148 } = (N484)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31147)? { N30780, N30781, N30782, N30783 } : 1'b0;
  assign N484 = N30880;
  assign { N31156, N31155, N31154, N31153 } = (N485)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31152)? { N30784, N30785, N30786, N30787 } : 1'b0;
  assign N485 = N30881;
  assign { N31161, N31160, N31159, N31158 } = (N486)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31157)? { N30788, N30789, N30790, N30791 } : 1'b0;
  assign N486 = N30882;
  assign { N31166, N31165, N31164, N31163 } = (N487)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31162)? { N30792, N30793, N30794, N30795 } : 1'b0;
  assign N487 = N30883;
  assign { N31171, N31170, N31169, N31168 } = (N488)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31167)? { N30796, N30797, N30798, N30799 } : 1'b0;
  assign N488 = N30884;
  assign { N31176, N31175, N31174, N31173 } = (N489)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31172)? { N30800, N30801, N30802, N30803 } : 1'b0;
  assign N489 = N30885;
  assign { N31181, N31180, N31179, N31178 } = (N490)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31177)? { N30804, N30805, N30806, N30807 } : 1'b0;
  assign N490 = N30886;
  assign { N31186, N31185, N31184, N31183 } = (N491)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31182)? { N30808, N30809, N30810, N30811 } : 1'b0;
  assign N491 = N30887;
  assign { N31191, N31190, N31189, N31188 } = (N492)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31187)? { N30812, N30813, N30814, N30815 } : 1'b0;
  assign N492 = N30888;
  assign { N31196, N31195, N31194, N31193 } = (N493)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31192)? { N30816, N30817, N30818, N30819 } : 1'b0;
  assign N493 = N30889;
  assign { N31201, N31200, N31199, N31198 } = (N494)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31197)? { N30820, N30821, N30822, N30823 } : 1'b0;
  assign N494 = N30890;
  assign { N31206, N31205, N31204, N31203 } = (N495)? { mem_q[1380:1380], mem_q[1381:1381], mem_q[1382:1382], mem_q[1383:1383] } : 
                                              (N31202)? { N30824, N30825, N30826, N30827 } : 1'b0;
  assign N495 = N30891;
  assign { N31458, N31457, N31456, N31455, N31454, N31453, N31452, N31451, N31450, N31449, N31448, N31447, N31446, N31445, N31444, N31443, N31442, N31441, N31440, N31439, N31438, N31437, N31436, N31435, N31434, N31433, N31432, N31431, N31430, N31429, N31428, N31427, N31426, N31425, N31424, N31423, N31422, N31421, N31420, N31419, N31418, N31417, N31416, N31415, N31414, N31413, N31412, N31411, N31410, N31409, N31408, N31407, N31406, N31405, N31404, N31403, N31402, N31401, N31400, N31399, N31398, N31397, N31396, N31395, N31394, N31393, N31392, N31391, N31390, N31389, N31388, N31387, N31386, N31385, N31384, N31383, N31382, N31381, N31380, N31379, N31378, N31377, N31376, N31375, N31374, N31373, N31372, N31371, N31370, N31369, N31368, N31367, N31366, N31365, N31364, N31363, N31362, N31361, N31360, N31359, N31358, N31357, N31356, N31355, N31354, N31353, N31352, N31351, N31350, N31349, N31348, N31347, N31346, N31345, N31344, N31343, N31342, N31341, N31340, N31339, N31338, N31337, N31336, N31335, N31334, N31333, N31332, N31331, N31330, N31329, N31328, N31327, N31326, N31325, N31324, N31323, N31322, N31321, N31320, N31319, N31318, N31317, N31316, N31315, N31314, N31313, N31312, N31311, N31310, N31309, N31308, N31307, N31306, N31305, N31304, N31303, N31302, N31301, N31300, N31299, N31298, N31297, N31296, N31295, N31294, N31293, N31292, N31291, N31290, N31289, N31288, N31287, N31286, N31285, N31284, N31283, N31282, N31281, N31280, N31279, N31278, N31277, N31276, N31275, N31274, N31273, N31272, N31271, N31270, N31269, N31268, N31267, N31266, N31265, N31264, N31263, N31262, N31261, N31260, N31259, N31258, N31257, N31256, N31255, N31254, N31253, N31252, N31251, N31250, N31249, N31248, N31247, N31246, N31245, N31244, N31243, N31242, N31241, N31240, N31239, N31238, N31237, N31236, N31235, N31234, N31233, N31232, N31231, N31230, N31229, N31228, N31227, N31226, N31225, N31224, N31223, N31222, N31221, N31220, N31219, N31218, N31217, N31216, N31215, N31214, N31213, N31212, N31211, N31210, N31209, N31208, N31207 } = (N496)? { N31203, N31204, N31205, N31206, N31198, N31199, N31200, N31201, N31193, N31194, N31195, N31196, N31188, N31189, N31190, N31191, N31183, N31184, N31185, N31186, N31178, N31179, N31180, N31181, N31173, N31174, N31175, N31176, N31168, N31169, N31170, N31171, N31163, N31164, N31165, N31166, N31158, N31159, N31160, N31161, N31153, N31154, N31155, N31156, N31148, N31149, N31150, N31151, N31143, N31144, N31145, N31146, N31138, N31139, N31140, N31141, N31133, N31134, N31135, N31136, N31128, N31129, N31130, N31131, N31123, N31124, N31125, N31126, N31118, N31119, N31120, N31121, N31113, N31114, N31115, N31116, N31108, N31109, N31110, N31111, N31103, N31104, N31105, N31106, N31098, N31099, N31100, N31101, N31093, N31094, N31095, N31096, N31088, N31089, N31090, N31091, N31083, N31084, N31085, N31086, N31078, N31079, N31080, N31081, N31073, N31074, N31075, N31076, N31068, N31069, N31070, N31071, N31063, N31064, N31065, N31066, N31058, N31059, N31060, N31061, N31053, N31054, N31055, N31056, N31048, N31049, N31050, N31051, N31043, N31044, N31045, N31046, N31038, N31039, N31040, N31041, N31033, N31034, N31035, N31036, N31028, N31029, N31030, N31031, N31023, N31024, N31025, N31026, N31018, N31019, N31020, N31021, N31013, N31014, N31015, N31016, N31008, N31009, N31010, N31011, N31003, N31004, N31005, N31006, N30998, N30999, N31000, N31001, N30993, N30994, N30995, N30996, N30988, N30989, N30990, N30991, N30983, N30984, N30985, N30986, N30978, N30979, N30980, N30981, N30973, N30974, N30975, N30976, N30968, N30969, N30970, N30971, N30963, N30964, N30965, N30966, N30958, N30959, N30960, N30961, N30953, N30954, N30955, N30956, N30948, N30949, N30950, N30951, N30943, N30944, N30945, N30946, N30938, N30939, N30940, N30941, N30933, N30934, N30935, N30936, N30928, N30929, N30930, N30931, N30923, N30924, N30925, N30926, N30918, N30919, N30920, N30921, N30913, N30914, N30915, N30916, N30908, N30909, N30910, N30911, N30903, N30904, N30905, N30906, N30898, N30899, N30900, N30901, N30893, N30894, N30895, N30896 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N30828)? { N30827, N30826, N30825, N30824, N30823, N30822, N30821, N30820, N30819, N30818, N30817, N30816, N30815, N30814, N30813, N30812, N30811, N30810, N30809, N30808, N30807, N30806, N30805, N30804, N30803, N30802, N30801, N30800, N30799, N30798, N30797, N30796, N30795, N30794, N30793, N30792, N30791, N30790, N30789, N30788, N30787, N30786, N30785, N30784, N30783, N30782, N30781, N30780, N30779, N30778, N30777, N30776, N30775, N30774, N30773, N30772, N30771, N30770, N30769, N30768, N30767, N30766, N30765, N30764, N30763, N30762, N30761, N30760, N30759, N30758, N30757, N30756, N30755, N30754, N30753, N30752, N30751, N30750, N30749, N30748, N30747, N30746, N30745, N30744, N30743, N30742, N30741, N30740, N30739, N30738, N30737, N30736, N30735, N30734, N30733, N30732, N30731, N30730, N30729, N30728, N30727, N30726, N30725, N30724, N30723, N30722, N30721, N30720, N30719, N30718, N30717, N30716, N30715, N30714, N30713, N30712, N30711, N30710, N30709, N30708, N30707, N30706, N30705, N30704, N30703, N30702, N30701, N30700, N30699, N30698, N30697, N30696, N30695, N30694, N30693, N30692, N30691, N30690, N30689, N30688, N30687, N30686, N30685, N30684, N30683, N30682, N30681, N30680, N30679, N30678, N30677, N30676, N30675, N30674, N30673, N30672, N30671, N30670, N30669, N30668, N30667, N30666, N30665, N30664, N30663, N30662, N30661, N30660, N30659, N30658, N30657, N30656, N30655, N30654, N30653, N30652, N30651, N30650, N30649, N30648, N30647, N30646, N30645, N30644, N30643, N30642, N30641, N30640, N30639, N30638, N30637, N30636, N30635, N30634, N30633, N30632, N30631, N30630, N30629, N30628, N30627, N30626, N30625, N30624, N30623, N30622, N30621, N30620, N30619, N30618, N30617, N30616, N30615, N30614, N30613, N30612, N30611, N30610, N30609, N30608, N30607, N30606, N30605, N30604, N30603, N30602, N30601, N30600, N30599, N30598, N30597, N30596, N30595, N30594, N30593, N30592, N30591, N30590, N30589, N30588, N30587, N30586, N30585, N30584, N30583, N30582, N30581, N30580, N30579, N30578, N30577, N30576 } : 1'b0;
  assign N496 = mem_q[1451];
  assign { N31527, N31526, N31525, N31524 } = (N497)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31523)? { N31207, N31208, N31209, N31210 } : 1'b0;
  assign N497 = N31460;
  assign { N31532, N31531, N31530, N31529 } = (N498)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31528)? { N31211, N31212, N31213, N31214 } : 1'b0;
  assign N498 = N31461;
  assign { N31537, N31536, N31535, N31534 } = (N499)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31533)? { N31215, N31216, N31217, N31218 } : 1'b0;
  assign N499 = N31462;
  assign { N31542, N31541, N31540, N31539 } = (N500)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31538)? { N31219, N31220, N31221, N31222 } : 1'b0;
  assign N500 = N31463;
  assign { N31547, N31546, N31545, N31544 } = (N501)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31543)? { N31223, N31224, N31225, N31226 } : 1'b0;
  assign N501 = N31464;
  assign { N31552, N31551, N31550, N31549 } = (N502)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31548)? { N31227, N31228, N31229, N31230 } : 1'b0;
  assign N502 = N31465;
  assign { N31557, N31556, N31555, N31554 } = (N503)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31553)? { N31231, N31232, N31233, N31234 } : 1'b0;
  assign N503 = N31466;
  assign { N31562, N31561, N31560, N31559 } = (N504)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31558)? { N31235, N31236, N31237, N31238 } : 1'b0;
  assign N504 = N31467;
  assign { N31567, N31566, N31565, N31564 } = (N505)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31563)? { N31239, N31240, N31241, N31242 } : 1'b0;
  assign N505 = N31468;
  assign { N31572, N31571, N31570, N31569 } = (N506)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31568)? { N31243, N31244, N31245, N31246 } : 1'b0;
  assign N506 = N31469;
  assign { N31577, N31576, N31575, N31574 } = (N507)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31573)? { N31247, N31248, N31249, N31250 } : 1'b0;
  assign N507 = N31470;
  assign { N31582, N31581, N31580, N31579 } = (N508)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31578)? { N31251, N31252, N31253, N31254 } : 1'b0;
  assign N508 = N31471;
  assign { N31587, N31586, N31585, N31584 } = (N509)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31583)? { N31255, N31256, N31257, N31258 } : 1'b0;
  assign N509 = N31472;
  assign { N31592, N31591, N31590, N31589 } = (N510)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31588)? { N31259, N31260, N31261, N31262 } : 1'b0;
  assign N510 = N31473;
  assign { N31597, N31596, N31595, N31594 } = (N511)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31593)? { N31263, N31264, N31265, N31266 } : 1'b0;
  assign N511 = N31474;
  assign { N31602, N31601, N31600, N31599 } = (N512)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31598)? { N31267, N31268, N31269, N31270 } : 1'b0;
  assign N512 = N31475;
  assign { N31607, N31606, N31605, N31604 } = (N513)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31603)? { N31271, N31272, N31273, N31274 } : 1'b0;
  assign N513 = N31476;
  assign { N31612, N31611, N31610, N31609 } = (N514)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31608)? { N31275, N31276, N31277, N31278 } : 1'b0;
  assign N514 = N31477;
  assign { N31617, N31616, N31615, N31614 } = (N515)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31613)? { N31279, N31280, N31281, N31282 } : 1'b0;
  assign N515 = N31478;
  assign { N31622, N31621, N31620, N31619 } = (N516)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31618)? { N31283, N31284, N31285, N31286 } : 1'b0;
  assign N516 = N31479;
  assign { N31627, N31626, N31625, N31624 } = (N517)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31623)? { N31287, N31288, N31289, N31290 } : 1'b0;
  assign N517 = N31480;
  assign { N31632, N31631, N31630, N31629 } = (N518)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31628)? { N31291, N31292, N31293, N31294 } : 1'b0;
  assign N518 = N31481;
  assign { N31637, N31636, N31635, N31634 } = (N519)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31633)? { N31295, N31296, N31297, N31298 } : 1'b0;
  assign N519 = N31482;
  assign { N31642, N31641, N31640, N31639 } = (N520)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31638)? { N31299, N31300, N31301, N31302 } : 1'b0;
  assign N520 = N31483;
  assign { N31647, N31646, N31645, N31644 } = (N521)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31643)? { N31303, N31304, N31305, N31306 } : 1'b0;
  assign N521 = N31484;
  assign { N31652, N31651, N31650, N31649 } = (N522)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31648)? { N31307, N31308, N31309, N31310 } : 1'b0;
  assign N522 = N31485;
  assign { N31657, N31656, N31655, N31654 } = (N523)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31653)? { N31311, N31312, N31313, N31314 } : 1'b0;
  assign N523 = N31486;
  assign { N31662, N31661, N31660, N31659 } = (N524)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31658)? { N31315, N31316, N31317, N31318 } : 1'b0;
  assign N524 = N31487;
  assign { N31667, N31666, N31665, N31664 } = (N525)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31663)? { N31319, N31320, N31321, N31322 } : 1'b0;
  assign N525 = N31488;
  assign { N31672, N31671, N31670, N31669 } = (N526)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31668)? { N31323, N31324, N31325, N31326 } : 1'b0;
  assign N526 = N31489;
  assign { N31677, N31676, N31675, N31674 } = (N527)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31673)? { N31327, N31328, N31329, N31330 } : 1'b0;
  assign N527 = N31490;
  assign { N31682, N31681, N31680, N31679 } = (N528)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31678)? { N31331, N31332, N31333, N31334 } : 1'b0;
  assign N528 = N31491;
  assign { N31687, N31686, N31685, N31684 } = (N529)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31683)? { N31335, N31336, N31337, N31338 } : 1'b0;
  assign N529 = N31492;
  assign { N31692, N31691, N31690, N31689 } = (N530)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31688)? { N31339, N31340, N31341, N31342 } : 1'b0;
  assign N530 = N31493;
  assign { N31697, N31696, N31695, N31694 } = (N531)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31693)? { N31343, N31344, N31345, N31346 } : 1'b0;
  assign N531 = N31494;
  assign { N31702, N31701, N31700, N31699 } = (N532)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31698)? { N31347, N31348, N31349, N31350 } : 1'b0;
  assign N532 = N31495;
  assign { N31707, N31706, N31705, N31704 } = (N533)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31703)? { N31351, N31352, N31353, N31354 } : 1'b0;
  assign N533 = N31496;
  assign { N31712, N31711, N31710, N31709 } = (N534)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31708)? { N31355, N31356, N31357, N31358 } : 1'b0;
  assign N534 = N31497;
  assign { N31717, N31716, N31715, N31714 } = (N535)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31713)? { N31359, N31360, N31361, N31362 } : 1'b0;
  assign N535 = N31498;
  assign { N31722, N31721, N31720, N31719 } = (N536)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31718)? { N31363, N31364, N31365, N31366 } : 1'b0;
  assign N536 = N31499;
  assign { N31727, N31726, N31725, N31724 } = (N537)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31723)? { N31367, N31368, N31369, N31370 } : 1'b0;
  assign N537 = N31500;
  assign { N31732, N31731, N31730, N31729 } = (N538)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31728)? { N31371, N31372, N31373, N31374 } : 1'b0;
  assign N538 = N31501;
  assign { N31737, N31736, N31735, N31734 } = (N539)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31733)? { N31375, N31376, N31377, N31378 } : 1'b0;
  assign N539 = N31502;
  assign { N31742, N31741, N31740, N31739 } = (N540)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31738)? { N31379, N31380, N31381, N31382 } : 1'b0;
  assign N540 = N31503;
  assign { N31747, N31746, N31745, N31744 } = (N541)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31743)? { N31383, N31384, N31385, N31386 } : 1'b0;
  assign N541 = N31504;
  assign { N31752, N31751, N31750, N31749 } = (N542)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31748)? { N31387, N31388, N31389, N31390 } : 1'b0;
  assign N542 = N31505;
  assign { N31757, N31756, N31755, N31754 } = (N543)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31753)? { N31391, N31392, N31393, N31394 } : 1'b0;
  assign N543 = N31506;
  assign { N31762, N31761, N31760, N31759 } = (N544)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31758)? { N31395, N31396, N31397, N31398 } : 1'b0;
  assign N544 = N31507;
  assign { N31767, N31766, N31765, N31764 } = (N545)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31763)? { N31399, N31400, N31401, N31402 } : 1'b0;
  assign N545 = N31508;
  assign { N31772, N31771, N31770, N31769 } = (N546)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31768)? { N31403, N31404, N31405, N31406 } : 1'b0;
  assign N546 = N31509;
  assign { N31777, N31776, N31775, N31774 } = (N547)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31773)? { N31407, N31408, N31409, N31410 } : 1'b0;
  assign N547 = N31510;
  assign { N31782, N31781, N31780, N31779 } = (N548)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31778)? { N31411, N31412, N31413, N31414 } : 1'b0;
  assign N548 = N31511;
  assign { N31787, N31786, N31785, N31784 } = (N549)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31783)? { N31415, N31416, N31417, N31418 } : 1'b0;
  assign N549 = N31512;
  assign { N31792, N31791, N31790, N31789 } = (N550)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31788)? { N31419, N31420, N31421, N31422 } : 1'b0;
  assign N550 = N31513;
  assign { N31797, N31796, N31795, N31794 } = (N551)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31793)? { N31423, N31424, N31425, N31426 } : 1'b0;
  assign N551 = N31514;
  assign { N31802, N31801, N31800, N31799 } = (N552)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31798)? { N31427, N31428, N31429, N31430 } : 1'b0;
  assign N552 = N31515;
  assign { N31807, N31806, N31805, N31804 } = (N553)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31803)? { N31431, N31432, N31433, N31434 } : 1'b0;
  assign N553 = N31516;
  assign { N31812, N31811, N31810, N31809 } = (N554)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31808)? { N31435, N31436, N31437, N31438 } : 1'b0;
  assign N554 = N31517;
  assign { N31817, N31816, N31815, N31814 } = (N555)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31813)? { N31439, N31440, N31441, N31442 } : 1'b0;
  assign N555 = N31518;
  assign { N31822, N31821, N31820, N31819 } = (N556)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31818)? { N31443, N31444, N31445, N31446 } : 1'b0;
  assign N556 = N31519;
  assign { N31827, N31826, N31825, N31824 } = (N557)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31823)? { N31447, N31448, N31449, N31450 } : 1'b0;
  assign N557 = N31520;
  assign { N31832, N31831, N31830, N31829 } = (N558)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31828)? { N31451, N31452, N31453, N31454 } : 1'b0;
  assign N558 = N31521;
  assign { N31837, N31836, N31835, N31834 } = (N559)? { mem_q[1743:1743], mem_q[1744:1744], mem_q[1745:1745], mem_q[1746:1746] } : 
                                              (N31833)? { N31455, N31456, N31457, N31458 } : 1'b0;
  assign N559 = N31522;
  assign { N32089, N32088, N32087, N32086, N32085, N32084, N32083, N32082, N32081, N32080, N32079, N32078, N32077, N32076, N32075, N32074, N32073, N32072, N32071, N32070, N32069, N32068, N32067, N32066, N32065, N32064, N32063, N32062, N32061, N32060, N32059, N32058, N32057, N32056, N32055, N32054, N32053, N32052, N32051, N32050, N32049, N32048, N32047, N32046, N32045, N32044, N32043, N32042, N32041, N32040, N32039, N32038, N32037, N32036, N32035, N32034, N32033, N32032, N32031, N32030, N32029, N32028, N32027, N32026, N32025, N32024, N32023, N32022, N32021, N32020, N32019, N32018, N32017, N32016, N32015, N32014, N32013, N32012, N32011, N32010, N32009, N32008, N32007, N32006, N32005, N32004, N32003, N32002, N32001, N32000, N31999, N31998, N31997, N31996, N31995, N31994, N31993, N31992, N31991, N31990, N31989, N31988, N31987, N31986, N31985, N31984, N31983, N31982, N31981, N31980, N31979, N31978, N31977, N31976, N31975, N31974, N31973, N31972, N31971, N31970, N31969, N31968, N31967, N31966, N31965, N31964, N31963, N31962, N31961, N31960, N31959, N31958, N31957, N31956, N31955, N31954, N31953, N31952, N31951, N31950, N31949, N31948, N31947, N31946, N31945, N31944, N31943, N31942, N31941, N31940, N31939, N31938, N31937, N31936, N31935, N31934, N31933, N31932, N31931, N31930, N31929, N31928, N31927, N31926, N31925, N31924, N31923, N31922, N31921, N31920, N31919, N31918, N31917, N31916, N31915, N31914, N31913, N31912, N31911, N31910, N31909, N31908, N31907, N31906, N31905, N31904, N31903, N31902, N31901, N31900, N31899, N31898, N31897, N31896, N31895, N31894, N31893, N31892, N31891, N31890, N31889, N31888, N31887, N31886, N31885, N31884, N31883, N31882, N31881, N31880, N31879, N31878, N31877, N31876, N31875, N31874, N31873, N31872, N31871, N31870, N31869, N31868, N31867, N31866, N31865, N31864, N31863, N31862, N31861, N31860, N31859, N31858, N31857, N31856, N31855, N31854, N31853, N31852, N31851, N31850, N31849, N31848, N31847, N31846, N31845, N31844, N31843, N31842, N31841, N31840, N31839, N31838 } = (N560)? { N31834, N31835, N31836, N31837, N31829, N31830, N31831, N31832, N31824, N31825, N31826, N31827, N31819, N31820, N31821, N31822, N31814, N31815, N31816, N31817, N31809, N31810, N31811, N31812, N31804, N31805, N31806, N31807, N31799, N31800, N31801, N31802, N31794, N31795, N31796, N31797, N31789, N31790, N31791, N31792, N31784, N31785, N31786, N31787, N31779, N31780, N31781, N31782, N31774, N31775, N31776, N31777, N31769, N31770, N31771, N31772, N31764, N31765, N31766, N31767, N31759, N31760, N31761, N31762, N31754, N31755, N31756, N31757, N31749, N31750, N31751, N31752, N31744, N31745, N31746, N31747, N31739, N31740, N31741, N31742, N31734, N31735, N31736, N31737, N31729, N31730, N31731, N31732, N31724, N31725, N31726, N31727, N31719, N31720, N31721, N31722, N31714, N31715, N31716, N31717, N31709, N31710, N31711, N31712, N31704, N31705, N31706, N31707, N31699, N31700, N31701, N31702, N31694, N31695, N31696, N31697, N31689, N31690, N31691, N31692, N31684, N31685, N31686, N31687, N31679, N31680, N31681, N31682, N31674, N31675, N31676, N31677, N31669, N31670, N31671, N31672, N31664, N31665, N31666, N31667, N31659, N31660, N31661, N31662, N31654, N31655, N31656, N31657, N31649, N31650, N31651, N31652, N31644, N31645, N31646, N31647, N31639, N31640, N31641, N31642, N31634, N31635, N31636, N31637, N31629, N31630, N31631, N31632, N31624, N31625, N31626, N31627, N31619, N31620, N31621, N31622, N31614, N31615, N31616, N31617, N31609, N31610, N31611, N31612, N31604, N31605, N31606, N31607, N31599, N31600, N31601, N31602, N31594, N31595, N31596, N31597, N31589, N31590, N31591, N31592, N31584, N31585, N31586, N31587, N31579, N31580, N31581, N31582, N31574, N31575, N31576, N31577, N31569, N31570, N31571, N31572, N31564, N31565, N31566, N31567, N31559, N31560, N31561, N31562, N31554, N31555, N31556, N31557, N31549, N31550, N31551, N31552, N31544, N31545, N31546, N31547, N31539, N31540, N31541, N31542, N31534, N31535, N31536, N31537, N31529, N31530, N31531, N31532, N31524, N31525, N31526, N31527 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N31459)? { N31458, N31457, N31456, N31455, N31454, N31453, N31452, N31451, N31450, N31449, N31448, N31447, N31446, N31445, N31444, N31443, N31442, N31441, N31440, N31439, N31438, N31437, N31436, N31435, N31434, N31433, N31432, N31431, N31430, N31429, N31428, N31427, N31426, N31425, N31424, N31423, N31422, N31421, N31420, N31419, N31418, N31417, N31416, N31415, N31414, N31413, N31412, N31411, N31410, N31409, N31408, N31407, N31406, N31405, N31404, N31403, N31402, N31401, N31400, N31399, N31398, N31397, N31396, N31395, N31394, N31393, N31392, N31391, N31390, N31389, N31388, N31387, N31386, N31385, N31384, N31383, N31382, N31381, N31380, N31379, N31378, N31377, N31376, N31375, N31374, N31373, N31372, N31371, N31370, N31369, N31368, N31367, N31366, N31365, N31364, N31363, N31362, N31361, N31360, N31359, N31358, N31357, N31356, N31355, N31354, N31353, N31352, N31351, N31350, N31349, N31348, N31347, N31346, N31345, N31344, N31343, N31342, N31341, N31340, N31339, N31338, N31337, N31336, N31335, N31334, N31333, N31332, N31331, N31330, N31329, N31328, N31327, N31326, N31325, N31324, N31323, N31322, N31321, N31320, N31319, N31318, N31317, N31316, N31315, N31314, N31313, N31312, N31311, N31310, N31309, N31308, N31307, N31306, N31305, N31304, N31303, N31302, N31301, N31300, N31299, N31298, N31297, N31296, N31295, N31294, N31293, N31292, N31291, N31290, N31289, N31288, N31287, N31286, N31285, N31284, N31283, N31282, N31281, N31280, N31279, N31278, N31277, N31276, N31275, N31274, N31273, N31272, N31271, N31270, N31269, N31268, N31267, N31266, N31265, N31264, N31263, N31262, N31261, N31260, N31259, N31258, N31257, N31256, N31255, N31254, N31253, N31252, N31251, N31250, N31249, N31248, N31247, N31246, N31245, N31244, N31243, N31242, N31241, N31240, N31239, N31238, N31237, N31236, N31235, N31234, N31233, N31232, N31231, N31230, N31229, N31228, N31227, N31226, N31225, N31224, N31223, N31222, N31221, N31220, N31219, N31218, N31217, N31216, N31215, N31214, N31213, N31212, N31211, N31210, N31209, N31208, N31207 } : 1'b0;
  assign N560 = mem_q[1814];
  assign { N32158, N32157, N32156, N32155 } = (N561)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32154)? { N31838, N31839, N31840, N31841 } : 1'b0;
  assign N561 = N32091;
  assign { N32163, N32162, N32161, N32160 } = (N562)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32159)? { N31842, N31843, N31844, N31845 } : 1'b0;
  assign N562 = N32092;
  assign { N32168, N32167, N32166, N32165 } = (N563)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32164)? { N31846, N31847, N31848, N31849 } : 1'b0;
  assign N563 = N32093;
  assign { N32173, N32172, N32171, N32170 } = (N564)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32169)? { N31850, N31851, N31852, N31853 } : 1'b0;
  assign N564 = N32094;
  assign { N32178, N32177, N32176, N32175 } = (N565)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32174)? { N31854, N31855, N31856, N31857 } : 1'b0;
  assign N565 = N32095;
  assign { N32183, N32182, N32181, N32180 } = (N566)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32179)? { N31858, N31859, N31860, N31861 } : 1'b0;
  assign N566 = N32096;
  assign { N32188, N32187, N32186, N32185 } = (N567)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32184)? { N31862, N31863, N31864, N31865 } : 1'b0;
  assign N567 = N32097;
  assign { N32193, N32192, N32191, N32190 } = (N568)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32189)? { N31866, N31867, N31868, N31869 } : 1'b0;
  assign N568 = N32098;
  assign { N32198, N32197, N32196, N32195 } = (N569)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32194)? { N31870, N31871, N31872, N31873 } : 1'b0;
  assign N569 = N32099;
  assign { N32203, N32202, N32201, N32200 } = (N570)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32199)? { N31874, N31875, N31876, N31877 } : 1'b0;
  assign N570 = N32100;
  assign { N32208, N32207, N32206, N32205 } = (N571)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32204)? { N31878, N31879, N31880, N31881 } : 1'b0;
  assign N571 = N32101;
  assign { N32213, N32212, N32211, N32210 } = (N572)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32209)? { N31882, N31883, N31884, N31885 } : 1'b0;
  assign N572 = N32102;
  assign { N32218, N32217, N32216, N32215 } = (N573)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32214)? { N31886, N31887, N31888, N31889 } : 1'b0;
  assign N573 = N32103;
  assign { N32223, N32222, N32221, N32220 } = (N574)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32219)? { N31890, N31891, N31892, N31893 } : 1'b0;
  assign N574 = N32104;
  assign { N32228, N32227, N32226, N32225 } = (N575)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32224)? { N31894, N31895, N31896, N31897 } : 1'b0;
  assign N575 = N32105;
  assign { N32233, N32232, N32231, N32230 } = (N576)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32229)? { N31898, N31899, N31900, N31901 } : 1'b0;
  assign N576 = N32106;
  assign { N32238, N32237, N32236, N32235 } = (N577)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32234)? { N31902, N31903, N31904, N31905 } : 1'b0;
  assign N577 = N32107;
  assign { N32243, N32242, N32241, N32240 } = (N578)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32239)? { N31906, N31907, N31908, N31909 } : 1'b0;
  assign N578 = N32108;
  assign { N32248, N32247, N32246, N32245 } = (N579)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32244)? { N31910, N31911, N31912, N31913 } : 1'b0;
  assign N579 = N32109;
  assign { N32253, N32252, N32251, N32250 } = (N580)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32249)? { N31914, N31915, N31916, N31917 } : 1'b0;
  assign N580 = N32110;
  assign { N32258, N32257, N32256, N32255 } = (N581)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32254)? { N31918, N31919, N31920, N31921 } : 1'b0;
  assign N581 = N32111;
  assign { N32263, N32262, N32261, N32260 } = (N582)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32259)? { N31922, N31923, N31924, N31925 } : 1'b0;
  assign N582 = N32112;
  assign { N32268, N32267, N32266, N32265 } = (N583)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32264)? { N31926, N31927, N31928, N31929 } : 1'b0;
  assign N583 = N32113;
  assign { N32273, N32272, N32271, N32270 } = (N584)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32269)? { N31930, N31931, N31932, N31933 } : 1'b0;
  assign N584 = N32114;
  assign { N32278, N32277, N32276, N32275 } = (N585)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32274)? { N31934, N31935, N31936, N31937 } : 1'b0;
  assign N585 = N32115;
  assign { N32283, N32282, N32281, N32280 } = (N586)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32279)? { N31938, N31939, N31940, N31941 } : 1'b0;
  assign N586 = N32116;
  assign { N32288, N32287, N32286, N32285 } = (N587)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32284)? { N31942, N31943, N31944, N31945 } : 1'b0;
  assign N587 = N32117;
  assign { N32293, N32292, N32291, N32290 } = (N588)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32289)? { N31946, N31947, N31948, N31949 } : 1'b0;
  assign N588 = N32118;
  assign { N32298, N32297, N32296, N32295 } = (N589)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32294)? { N31950, N31951, N31952, N31953 } : 1'b0;
  assign N589 = N32119;
  assign { N32303, N32302, N32301, N32300 } = (N590)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32299)? { N31954, N31955, N31956, N31957 } : 1'b0;
  assign N590 = N32120;
  assign { N32308, N32307, N32306, N32305 } = (N591)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32304)? { N31958, N31959, N31960, N31961 } : 1'b0;
  assign N591 = N32121;
  assign { N32313, N32312, N32311, N32310 } = (N592)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32309)? { N31962, N31963, N31964, N31965 } : 1'b0;
  assign N592 = N32122;
  assign { N32318, N32317, N32316, N32315 } = (N593)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32314)? { N31966, N31967, N31968, N31969 } : 1'b0;
  assign N593 = N32123;
  assign { N32323, N32322, N32321, N32320 } = (N594)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32319)? { N31970, N31971, N31972, N31973 } : 1'b0;
  assign N594 = N32124;
  assign { N32328, N32327, N32326, N32325 } = (N595)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32324)? { N31974, N31975, N31976, N31977 } : 1'b0;
  assign N595 = N32125;
  assign { N32333, N32332, N32331, N32330 } = (N596)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32329)? { N31978, N31979, N31980, N31981 } : 1'b0;
  assign N596 = N32126;
  assign { N32338, N32337, N32336, N32335 } = (N597)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32334)? { N31982, N31983, N31984, N31985 } : 1'b0;
  assign N597 = N32127;
  assign { N32343, N32342, N32341, N32340 } = (N598)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32339)? { N31986, N31987, N31988, N31989 } : 1'b0;
  assign N598 = N32128;
  assign { N32348, N32347, N32346, N32345 } = (N599)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32344)? { N31990, N31991, N31992, N31993 } : 1'b0;
  assign N599 = N32129;
  assign { N32353, N32352, N32351, N32350 } = (N600)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32349)? { N31994, N31995, N31996, N31997 } : 1'b0;
  assign N600 = N32130;
  assign { N32358, N32357, N32356, N32355 } = (N601)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32354)? { N31998, N31999, N32000, N32001 } : 1'b0;
  assign N601 = N32131;
  assign { N32363, N32362, N32361, N32360 } = (N602)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32359)? { N32002, N32003, N32004, N32005 } : 1'b0;
  assign N602 = N32132;
  assign { N32368, N32367, N32366, N32365 } = (N603)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32364)? { N32006, N32007, N32008, N32009 } : 1'b0;
  assign N603 = N32133;
  assign { N32373, N32372, N32371, N32370 } = (N604)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32369)? { N32010, N32011, N32012, N32013 } : 1'b0;
  assign N604 = N32134;
  assign { N32378, N32377, N32376, N32375 } = (N605)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32374)? { N32014, N32015, N32016, N32017 } : 1'b0;
  assign N605 = N32135;
  assign { N32383, N32382, N32381, N32380 } = (N606)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32379)? { N32018, N32019, N32020, N32021 } : 1'b0;
  assign N606 = N32136;
  assign { N32388, N32387, N32386, N32385 } = (N607)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32384)? { N32022, N32023, N32024, N32025 } : 1'b0;
  assign N607 = N32137;
  assign { N32393, N32392, N32391, N32390 } = (N608)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32389)? { N32026, N32027, N32028, N32029 } : 1'b0;
  assign N608 = N32138;
  assign { N32398, N32397, N32396, N32395 } = (N609)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32394)? { N32030, N32031, N32032, N32033 } : 1'b0;
  assign N609 = N32139;
  assign { N32403, N32402, N32401, N32400 } = (N610)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32399)? { N32034, N32035, N32036, N32037 } : 1'b0;
  assign N610 = N32140;
  assign { N32408, N32407, N32406, N32405 } = (N611)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32404)? { N32038, N32039, N32040, N32041 } : 1'b0;
  assign N611 = N32141;
  assign { N32413, N32412, N32411, N32410 } = (N612)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32409)? { N32042, N32043, N32044, N32045 } : 1'b0;
  assign N612 = N32142;
  assign { N32418, N32417, N32416, N32415 } = (N613)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32414)? { N32046, N32047, N32048, N32049 } : 1'b0;
  assign N613 = N32143;
  assign { N32423, N32422, N32421, N32420 } = (N614)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32419)? { N32050, N32051, N32052, N32053 } : 1'b0;
  assign N614 = N32144;
  assign { N32428, N32427, N32426, N32425 } = (N615)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32424)? { N32054, N32055, N32056, N32057 } : 1'b0;
  assign N615 = N32145;
  assign { N32433, N32432, N32431, N32430 } = (N616)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32429)? { N32058, N32059, N32060, N32061 } : 1'b0;
  assign N616 = N32146;
  assign { N32438, N32437, N32436, N32435 } = (N617)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32434)? { N32062, N32063, N32064, N32065 } : 1'b0;
  assign N617 = N32147;
  assign { N32443, N32442, N32441, N32440 } = (N618)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32439)? { N32066, N32067, N32068, N32069 } : 1'b0;
  assign N618 = N32148;
  assign { N32448, N32447, N32446, N32445 } = (N619)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32444)? { N32070, N32071, N32072, N32073 } : 1'b0;
  assign N619 = N32149;
  assign { N32453, N32452, N32451, N32450 } = (N620)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32449)? { N32074, N32075, N32076, N32077 } : 1'b0;
  assign N620 = N32150;
  assign { N32458, N32457, N32456, N32455 } = (N621)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32454)? { N32078, N32079, N32080, N32081 } : 1'b0;
  assign N621 = N32151;
  assign { N32463, N32462, N32461, N32460 } = (N622)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32459)? { N32082, N32083, N32084, N32085 } : 1'b0;
  assign N622 = N32152;
  assign { N32468, N32467, N32466, N32465 } = (N623)? { mem_q[2106:2106], mem_q[2107:2107], mem_q[2108:2108], mem_q[2109:2109] } : 
                                              (N32464)? { N32086, N32087, N32088, N32089 } : 1'b0;
  assign N623 = N32153;
  assign { N32720, N32719, N32718, N32717, N32716, N32715, N32714, N32713, N32712, N32711, N32710, N32709, N32708, N32707, N32706, N32705, N32704, N32703, N32702, N32701, N32700, N32699, N32698, N32697, N32696, N32695, N32694, N32693, N32692, N32691, N32690, N32689, N32688, N32687, N32686, N32685, N32684, N32683, N32682, N32681, N32680, N32679, N32678, N32677, N32676, N32675, N32674, N32673, N32672, N32671, N32670, N32669, N32668, N32667, N32666, N32665, N32664, N32663, N32662, N32661, N32660, N32659, N32658, N32657, N32656, N32655, N32654, N32653, N32652, N32651, N32650, N32649, N32648, N32647, N32646, N32645, N32644, N32643, N32642, N32641, N32640, N32639, N32638, N32637, N32636, N32635, N32634, N32633, N32632, N32631, N32630, N32629, N32628, N32627, N32626, N32625, N32624, N32623, N32622, N32621, N32620, N32619, N32618, N32617, N32616, N32615, N32614, N32613, N32612, N32611, N32610, N32609, N32608, N32607, N32606, N32605, N32604, N32603, N32602, N32601, N32600, N32599, N32598, N32597, N32596, N32595, N32594, N32593, N32592, N32591, N32590, N32589, N32588, N32587, N32586, N32585, N32584, N32583, N32582, N32581, N32580, N32579, N32578, N32577, N32576, N32575, N32574, N32573, N32572, N32571, N32570, N32569, N32568, N32567, N32566, N32565, N32564, N32563, N32562, N32561, N32560, N32559, N32558, N32557, N32556, N32555, N32554, N32553, N32552, N32551, N32550, N32549, N32548, N32547, N32546, N32545, N32544, N32543, N32542, N32541, N32540, N32539, N32538, N32537, N32536, N32535, N32534, N32533, N32532, N32531, N32530, N32529, N32528, N32527, N32526, N32525, N32524, N32523, N32522, N32521, N32520, N32519, N32518, N32517, N32516, N32515, N32514, N32513, N32512, N32511, N32510, N32509, N32508, N32507, N32506, N32505, N32504, N32503, N32502, N32501, N32500, N32499, N32498, N32497, N32496, N32495, N32494, N32493, N32492, N32491, N32490, N32489, N32488, N32487, N32486, N32485, N32484, N32483, N32482, N32481, N32480, N32479, N32478, N32477, N32476, N32475, N32474, N32473, N32472, N32471, N32470, N32469 } = (N624)? { N32465, N32466, N32467, N32468, N32460, N32461, N32462, N32463, N32455, N32456, N32457, N32458, N32450, N32451, N32452, N32453, N32445, N32446, N32447, N32448, N32440, N32441, N32442, N32443, N32435, N32436, N32437, N32438, N32430, N32431, N32432, N32433, N32425, N32426, N32427, N32428, N32420, N32421, N32422, N32423, N32415, N32416, N32417, N32418, N32410, N32411, N32412, N32413, N32405, N32406, N32407, N32408, N32400, N32401, N32402, N32403, N32395, N32396, N32397, N32398, N32390, N32391, N32392, N32393, N32385, N32386, N32387, N32388, N32380, N32381, N32382, N32383, N32375, N32376, N32377, N32378, N32370, N32371, N32372, N32373, N32365, N32366, N32367, N32368, N32360, N32361, N32362, N32363, N32355, N32356, N32357, N32358, N32350, N32351, N32352, N32353, N32345, N32346, N32347, N32348, N32340, N32341, N32342, N32343, N32335, N32336, N32337, N32338, N32330, N32331, N32332, N32333, N32325, N32326, N32327, N32328, N32320, N32321, N32322, N32323, N32315, N32316, N32317, N32318, N32310, N32311, N32312, N32313, N32305, N32306, N32307, N32308, N32300, N32301, N32302, N32303, N32295, N32296, N32297, N32298, N32290, N32291, N32292, N32293, N32285, N32286, N32287, N32288, N32280, N32281, N32282, N32283, N32275, N32276, N32277, N32278, N32270, N32271, N32272, N32273, N32265, N32266, N32267, N32268, N32260, N32261, N32262, N32263, N32255, N32256, N32257, N32258, N32250, N32251, N32252, N32253, N32245, N32246, N32247, N32248, N32240, N32241, N32242, N32243, N32235, N32236, N32237, N32238, N32230, N32231, N32232, N32233, N32225, N32226, N32227, N32228, N32220, N32221, N32222, N32223, N32215, N32216, N32217, N32218, N32210, N32211, N32212, N32213, N32205, N32206, N32207, N32208, N32200, N32201, N32202, N32203, N32195, N32196, N32197, N32198, N32190, N32191, N32192, N32193, N32185, N32186, N32187, N32188, N32180, N32181, N32182, N32183, N32175, N32176, N32177, N32178, N32170, N32171, N32172, N32173, N32165, N32166, N32167, N32168, N32160, N32161, N32162, N32163, N32155, N32156, N32157, N32158 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N32090)? { N32089, N32088, N32087, N32086, N32085, N32084, N32083, N32082, N32081, N32080, N32079, N32078, N32077, N32076, N32075, N32074, N32073, N32072, N32071, N32070, N32069, N32068, N32067, N32066, N32065, N32064, N32063, N32062, N32061, N32060, N32059, N32058, N32057, N32056, N32055, N32054, N32053, N32052, N32051, N32050, N32049, N32048, N32047, N32046, N32045, N32044, N32043, N32042, N32041, N32040, N32039, N32038, N32037, N32036, N32035, N32034, N32033, N32032, N32031, N32030, N32029, N32028, N32027, N32026, N32025, N32024, N32023, N32022, N32021, N32020, N32019, N32018, N32017, N32016, N32015, N32014, N32013, N32012, N32011, N32010, N32009, N32008, N32007, N32006, N32005, N32004, N32003, N32002, N32001, N32000, N31999, N31998, N31997, N31996, N31995, N31994, N31993, N31992, N31991, N31990, N31989, N31988, N31987, N31986, N31985, N31984, N31983, N31982, N31981, N31980, N31979, N31978, N31977, N31976, N31975, N31974, N31973, N31972, N31971, N31970, N31969, N31968, N31967, N31966, N31965, N31964, N31963, N31962, N31961, N31960, N31959, N31958, N31957, N31956, N31955, N31954, N31953, N31952, N31951, N31950, N31949, N31948, N31947, N31946, N31945, N31944, N31943, N31942, N31941, N31940, N31939, N31938, N31937, N31936, N31935, N31934, N31933, N31932, N31931, N31930, N31929, N31928, N31927, N31926, N31925, N31924, N31923, N31922, N31921, N31920, N31919, N31918, N31917, N31916, N31915, N31914, N31913, N31912, N31911, N31910, N31909, N31908, N31907, N31906, N31905, N31904, N31903, N31902, N31901, N31900, N31899, N31898, N31897, N31896, N31895, N31894, N31893, N31892, N31891, N31890, N31889, N31888, N31887, N31886, N31885, N31884, N31883, N31882, N31881, N31880, N31879, N31878, N31877, N31876, N31875, N31874, N31873, N31872, N31871, N31870, N31869, N31868, N31867, N31866, N31865, N31864, N31863, N31862, N31861, N31860, N31859, N31858, N31857, N31856, N31855, N31854, N31853, N31852, N31851, N31850, N31849, N31848, N31847, N31846, N31845, N31844, N31843, N31842, N31841, N31840, N31839, N31838 } : 1'b0;
  assign N624 = mem_q[2177];
  assign { N32789, N32788, N32787, N32786 } = (N625)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32785)? { N32469, N32470, N32471, N32472 } : 1'b0;
  assign N625 = N32722;
  assign { N32794, N32793, N32792, N32791 } = (N626)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32790)? { N32473, N32474, N32475, N32476 } : 1'b0;
  assign N626 = N32723;
  assign { N32799, N32798, N32797, N32796 } = (N627)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32795)? { N32477, N32478, N32479, N32480 } : 1'b0;
  assign N627 = N32724;
  assign { N32804, N32803, N32802, N32801 } = (N628)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32800)? { N32481, N32482, N32483, N32484 } : 1'b0;
  assign N628 = N32725;
  assign { N32809, N32808, N32807, N32806 } = (N629)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32805)? { N32485, N32486, N32487, N32488 } : 1'b0;
  assign N629 = N32726;
  assign { N32814, N32813, N32812, N32811 } = (N630)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32810)? { N32489, N32490, N32491, N32492 } : 1'b0;
  assign N630 = N32727;
  assign { N32819, N32818, N32817, N32816 } = (N631)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32815)? { N32493, N32494, N32495, N32496 } : 1'b0;
  assign N631 = N32728;
  assign { N32824, N32823, N32822, N32821 } = (N632)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32820)? { N32497, N32498, N32499, N32500 } : 1'b0;
  assign N632 = N32729;
  assign { N32829, N32828, N32827, N32826 } = (N633)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32825)? { N32501, N32502, N32503, N32504 } : 1'b0;
  assign N633 = N32730;
  assign { N32834, N32833, N32832, N32831 } = (N634)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32830)? { N32505, N32506, N32507, N32508 } : 1'b0;
  assign N634 = N32731;
  assign { N32839, N32838, N32837, N32836 } = (N635)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32835)? { N32509, N32510, N32511, N32512 } : 1'b0;
  assign N635 = N32732;
  assign { N32844, N32843, N32842, N32841 } = (N636)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32840)? { N32513, N32514, N32515, N32516 } : 1'b0;
  assign N636 = N32733;
  assign { N32849, N32848, N32847, N32846 } = (N637)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32845)? { N32517, N32518, N32519, N32520 } : 1'b0;
  assign N637 = N32734;
  assign { N32854, N32853, N32852, N32851 } = (N638)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32850)? { N32521, N32522, N32523, N32524 } : 1'b0;
  assign N638 = N32735;
  assign { N32859, N32858, N32857, N32856 } = (N639)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32855)? { N32525, N32526, N32527, N32528 } : 1'b0;
  assign N639 = N32736;
  assign { N32864, N32863, N32862, N32861 } = (N640)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32860)? { N32529, N32530, N32531, N32532 } : 1'b0;
  assign N640 = N32737;
  assign { N32869, N32868, N32867, N32866 } = (N641)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32865)? { N32533, N32534, N32535, N32536 } : 1'b0;
  assign N641 = N32738;
  assign { N32874, N32873, N32872, N32871 } = (N642)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32870)? { N32537, N32538, N32539, N32540 } : 1'b0;
  assign N642 = N32739;
  assign { N32879, N32878, N32877, N32876 } = (N643)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32875)? { N32541, N32542, N32543, N32544 } : 1'b0;
  assign N643 = N32740;
  assign { N32884, N32883, N32882, N32881 } = (N644)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32880)? { N32545, N32546, N32547, N32548 } : 1'b0;
  assign N644 = N32741;
  assign { N32889, N32888, N32887, N32886 } = (N645)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32885)? { N32549, N32550, N32551, N32552 } : 1'b0;
  assign N645 = N32742;
  assign { N32894, N32893, N32892, N32891 } = (N646)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32890)? { N32553, N32554, N32555, N32556 } : 1'b0;
  assign N646 = N32743;
  assign { N32899, N32898, N32897, N32896 } = (N647)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32895)? { N32557, N32558, N32559, N32560 } : 1'b0;
  assign N647 = N32744;
  assign { N32904, N32903, N32902, N32901 } = (N648)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32900)? { N32561, N32562, N32563, N32564 } : 1'b0;
  assign N648 = N32745;
  assign { N32909, N32908, N32907, N32906 } = (N649)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32905)? { N32565, N32566, N32567, N32568 } : 1'b0;
  assign N649 = N32746;
  assign { N32914, N32913, N32912, N32911 } = (N650)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32910)? { N32569, N32570, N32571, N32572 } : 1'b0;
  assign N650 = N32747;
  assign { N32919, N32918, N32917, N32916 } = (N651)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32915)? { N32573, N32574, N32575, N32576 } : 1'b0;
  assign N651 = N32748;
  assign { N32924, N32923, N32922, N32921 } = (N652)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32920)? { N32577, N32578, N32579, N32580 } : 1'b0;
  assign N652 = N32749;
  assign { N32929, N32928, N32927, N32926 } = (N653)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32925)? { N32581, N32582, N32583, N32584 } : 1'b0;
  assign N653 = N32750;
  assign { N32934, N32933, N32932, N32931 } = (N654)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32930)? { N32585, N32586, N32587, N32588 } : 1'b0;
  assign N654 = N32751;
  assign { N32939, N32938, N32937, N32936 } = (N655)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32935)? { N32589, N32590, N32591, N32592 } : 1'b0;
  assign N655 = N32752;
  assign { N32944, N32943, N32942, N32941 } = (N656)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32940)? { N32593, N32594, N32595, N32596 } : 1'b0;
  assign N656 = N32753;
  assign { N32949, N32948, N32947, N32946 } = (N657)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32945)? { N32597, N32598, N32599, N32600 } : 1'b0;
  assign N657 = N32754;
  assign { N32954, N32953, N32952, N32951 } = (N658)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32950)? { N32601, N32602, N32603, N32604 } : 1'b0;
  assign N658 = N32755;
  assign { N32959, N32958, N32957, N32956 } = (N659)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32955)? { N32605, N32606, N32607, N32608 } : 1'b0;
  assign N659 = N32756;
  assign { N32964, N32963, N32962, N32961 } = (N660)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32960)? { N32609, N32610, N32611, N32612 } : 1'b0;
  assign N660 = N32757;
  assign { N32969, N32968, N32967, N32966 } = (N661)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32965)? { N32613, N32614, N32615, N32616 } : 1'b0;
  assign N661 = N32758;
  assign { N32974, N32973, N32972, N32971 } = (N662)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32970)? { N32617, N32618, N32619, N32620 } : 1'b0;
  assign N662 = N32759;
  assign { N32979, N32978, N32977, N32976 } = (N663)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32975)? { N32621, N32622, N32623, N32624 } : 1'b0;
  assign N663 = N32760;
  assign { N32984, N32983, N32982, N32981 } = (N664)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32980)? { N32625, N32626, N32627, N32628 } : 1'b0;
  assign N664 = N32761;
  assign { N32989, N32988, N32987, N32986 } = (N665)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32985)? { N32629, N32630, N32631, N32632 } : 1'b0;
  assign N665 = N32762;
  assign { N32994, N32993, N32992, N32991 } = (N666)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32990)? { N32633, N32634, N32635, N32636 } : 1'b0;
  assign N666 = N32763;
  assign { N32999, N32998, N32997, N32996 } = (N667)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N32995)? { N32637, N32638, N32639, N32640 } : 1'b0;
  assign N667 = N32764;
  assign { N33004, N33003, N33002, N33001 } = (N668)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33000)? { N32641, N32642, N32643, N32644 } : 1'b0;
  assign N668 = N32765;
  assign { N33009, N33008, N33007, N33006 } = (N669)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33005)? { N32645, N32646, N32647, N32648 } : 1'b0;
  assign N669 = N32766;
  assign { N33014, N33013, N33012, N33011 } = (N670)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33010)? { N32649, N32650, N32651, N32652 } : 1'b0;
  assign N670 = N32767;
  assign { N33019, N33018, N33017, N33016 } = (N671)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33015)? { N32653, N32654, N32655, N32656 } : 1'b0;
  assign N671 = N32768;
  assign { N33024, N33023, N33022, N33021 } = (N672)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33020)? { N32657, N32658, N32659, N32660 } : 1'b0;
  assign N672 = N32769;
  assign { N33029, N33028, N33027, N33026 } = (N673)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33025)? { N32661, N32662, N32663, N32664 } : 1'b0;
  assign N673 = N32770;
  assign { N33034, N33033, N33032, N33031 } = (N674)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33030)? { N32665, N32666, N32667, N32668 } : 1'b0;
  assign N674 = N32771;
  assign { N33039, N33038, N33037, N33036 } = (N675)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33035)? { N32669, N32670, N32671, N32672 } : 1'b0;
  assign N675 = N32772;
  assign { N33044, N33043, N33042, N33041 } = (N676)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33040)? { N32673, N32674, N32675, N32676 } : 1'b0;
  assign N676 = N32773;
  assign { N33049, N33048, N33047, N33046 } = (N677)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33045)? { N32677, N32678, N32679, N32680 } : 1'b0;
  assign N677 = N32774;
  assign { N33054, N33053, N33052, N33051 } = (N678)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33050)? { N32681, N32682, N32683, N32684 } : 1'b0;
  assign N678 = N32775;
  assign { N33059, N33058, N33057, N33056 } = (N679)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33055)? { N32685, N32686, N32687, N32688 } : 1'b0;
  assign N679 = N32776;
  assign { N33064, N33063, N33062, N33061 } = (N680)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33060)? { N32689, N32690, N32691, N32692 } : 1'b0;
  assign N680 = N32777;
  assign { N33069, N33068, N33067, N33066 } = (N681)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33065)? { N32693, N32694, N32695, N32696 } : 1'b0;
  assign N681 = N32778;
  assign { N33074, N33073, N33072, N33071 } = (N682)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33070)? { N32697, N32698, N32699, N32700 } : 1'b0;
  assign N682 = N32779;
  assign { N33079, N33078, N33077, N33076 } = (N683)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33075)? { N32701, N32702, N32703, N32704 } : 1'b0;
  assign N683 = N32780;
  assign { N33084, N33083, N33082, N33081 } = (N684)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33080)? { N32705, N32706, N32707, N32708 } : 1'b0;
  assign N684 = N32781;
  assign { N33089, N33088, N33087, N33086 } = (N685)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33085)? { N32709, N32710, N32711, N32712 } : 1'b0;
  assign N685 = N32782;
  assign { N33094, N33093, N33092, N33091 } = (N686)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33090)? { N32713, N32714, N32715, N32716 } : 1'b0;
  assign N686 = N32783;
  assign { N33099, N33098, N33097, N33096 } = (N687)? { mem_q[2469:2469], mem_q[2470:2470], mem_q[2471:2471], mem_q[2472:2472] } : 
                                              (N33095)? { N32717, N32718, N32719, N32720 } : 1'b0;
  assign N687 = N32784;
  assign { N33351, N33350, N33349, N33348, N33347, N33346, N33345, N33344, N33343, N33342, N33341, N33340, N33339, N33338, N33337, N33336, N33335, N33334, N33333, N33332, N33331, N33330, N33329, N33328, N33327, N33326, N33325, N33324, N33323, N33322, N33321, N33320, N33319, N33318, N33317, N33316, N33315, N33314, N33313, N33312, N33311, N33310, N33309, N33308, N33307, N33306, N33305, N33304, N33303, N33302, N33301, N33300, N33299, N33298, N33297, N33296, N33295, N33294, N33293, N33292, N33291, N33290, N33289, N33288, N33287, N33286, N33285, N33284, N33283, N33282, N33281, N33280, N33279, N33278, N33277, N33276, N33275, N33274, N33273, N33272, N33271, N33270, N33269, N33268, N33267, N33266, N33265, N33264, N33263, N33262, N33261, N33260, N33259, N33258, N33257, N33256, N33255, N33254, N33253, N33252, N33251, N33250, N33249, N33248, N33247, N33246, N33245, N33244, N33243, N33242, N33241, N33240, N33239, N33238, N33237, N33236, N33235, N33234, N33233, N33232, N33231, N33230, N33229, N33228, N33227, N33226, N33225, N33224, N33223, N33222, N33221, N33220, N33219, N33218, N33217, N33216, N33215, N33214, N33213, N33212, N33211, N33210, N33209, N33208, N33207, N33206, N33205, N33204, N33203, N33202, N33201, N33200, N33199, N33198, N33197, N33196, N33195, N33194, N33193, N33192, N33191, N33190, N33189, N33188, N33187, N33186, N33185, N33184, N33183, N33182, N33181, N33180, N33179, N33178, N33177, N33176, N33175, N33174, N33173, N33172, N33171, N33170, N33169, N33168, N33167, N33166, N33165, N33164, N33163, N33162, N33161, N33160, N33159, N33158, N33157, N33156, N33155, N33154, N33153, N33152, N33151, N33150, N33149, N33148, N33147, N33146, N33145, N33144, N33143, N33142, N33141, N33140, N33139, N33138, N33137, N33136, N33135, N33134, N33133, N33132, N33131, N33130, N33129, N33128, N33127, N33126, N33125, N33124, N33123, N33122, N33121, N33120, N33119, N33118, N33117, N33116, N33115, N33114, N33113, N33112, N33111, N33110, N33109, N33108, N33107, N33106, N33105, N33104, N33103, N33102, N33101, N33100 } = (N688)? { N33096, N33097, N33098, N33099, N33091, N33092, N33093, N33094, N33086, N33087, N33088, N33089, N33081, N33082, N33083, N33084, N33076, N33077, N33078, N33079, N33071, N33072, N33073, N33074, N33066, N33067, N33068, N33069, N33061, N33062, N33063, N33064, N33056, N33057, N33058, N33059, N33051, N33052, N33053, N33054, N33046, N33047, N33048, N33049, N33041, N33042, N33043, N33044, N33036, N33037, N33038, N33039, N33031, N33032, N33033, N33034, N33026, N33027, N33028, N33029, N33021, N33022, N33023, N33024, N33016, N33017, N33018, N33019, N33011, N33012, N33013, N33014, N33006, N33007, N33008, N33009, N33001, N33002, N33003, N33004, N32996, N32997, N32998, N32999, N32991, N32992, N32993, N32994, N32986, N32987, N32988, N32989, N32981, N32982, N32983, N32984, N32976, N32977, N32978, N32979, N32971, N32972, N32973, N32974, N32966, N32967, N32968, N32969, N32961, N32962, N32963, N32964, N32956, N32957, N32958, N32959, N32951, N32952, N32953, N32954, N32946, N32947, N32948, N32949, N32941, N32942, N32943, N32944, N32936, N32937, N32938, N32939, N32931, N32932, N32933, N32934, N32926, N32927, N32928, N32929, N32921, N32922, N32923, N32924, N32916, N32917, N32918, N32919, N32911, N32912, N32913, N32914, N32906, N32907, N32908, N32909, N32901, N32902, N32903, N32904, N32896, N32897, N32898, N32899, N32891, N32892, N32893, N32894, N32886, N32887, N32888, N32889, N32881, N32882, N32883, N32884, N32876, N32877, N32878, N32879, N32871, N32872, N32873, N32874, N32866, N32867, N32868, N32869, N32861, N32862, N32863, N32864, N32856, N32857, N32858, N32859, N32851, N32852, N32853, N32854, N32846, N32847, N32848, N32849, N32841, N32842, N32843, N32844, N32836, N32837, N32838, N32839, N32831, N32832, N32833, N32834, N32826, N32827, N32828, N32829, N32821, N32822, N32823, N32824, N32816, N32817, N32818, N32819, N32811, N32812, N32813, N32814, N32806, N32807, N32808, N32809, N32801, N32802, N32803, N32804, N32796, N32797, N32798, N32799, N32791, N32792, N32793, N32794, N32786, N32787, N32788, N32789 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N32721)? { N32720, N32719, N32718, N32717, N32716, N32715, N32714, N32713, N32712, N32711, N32710, N32709, N32708, N32707, N32706, N32705, N32704, N32703, N32702, N32701, N32700, N32699, N32698, N32697, N32696, N32695, N32694, N32693, N32692, N32691, N32690, N32689, N32688, N32687, N32686, N32685, N32684, N32683, N32682, N32681, N32680, N32679, N32678, N32677, N32676, N32675, N32674, N32673, N32672, N32671, N32670, N32669, N32668, N32667, N32666, N32665, N32664, N32663, N32662, N32661, N32660, N32659, N32658, N32657, N32656, N32655, N32654, N32653, N32652, N32651, N32650, N32649, N32648, N32647, N32646, N32645, N32644, N32643, N32642, N32641, N32640, N32639, N32638, N32637, N32636, N32635, N32634, N32633, N32632, N32631, N32630, N32629, N32628, N32627, N32626, N32625, N32624, N32623, N32622, N32621, N32620, N32619, N32618, N32617, N32616, N32615, N32614, N32613, N32612, N32611, N32610, N32609, N32608, N32607, N32606, N32605, N32604, N32603, N32602, N32601, N32600, N32599, N32598, N32597, N32596, N32595, N32594, N32593, N32592, N32591, N32590, N32589, N32588, N32587, N32586, N32585, N32584, N32583, N32582, N32581, N32580, N32579, N32578, N32577, N32576, N32575, N32574, N32573, N32572, N32571, N32570, N32569, N32568, N32567, N32566, N32565, N32564, N32563, N32562, N32561, N32560, N32559, N32558, N32557, N32556, N32555, N32554, N32553, N32552, N32551, N32550, N32549, N32548, N32547, N32546, N32545, N32544, N32543, N32542, N32541, N32540, N32539, N32538, N32537, N32536, N32535, N32534, N32533, N32532, N32531, N32530, N32529, N32528, N32527, N32526, N32525, N32524, N32523, N32522, N32521, N32520, N32519, N32518, N32517, N32516, N32515, N32514, N32513, N32512, N32511, N32510, N32509, N32508, N32507, N32506, N32505, N32504, N32503, N32502, N32501, N32500, N32499, N32498, N32497, N32496, N32495, N32494, N32493, N32492, N32491, N32490, N32489, N32488, N32487, N32486, N32485, N32484, N32483, N32482, N32481, N32480, N32479, N32478, N32477, N32476, N32475, N32474, N32473, N32472, N32471, N32470, N32469 } : 1'b0;
  assign N688 = mem_q[2540];
  assign { N33420, N33419, N33418, N33417 } = (N689)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33416)? { N33100, N33101, N33102, N33103 } : 1'b0;
  assign N689 = N33353;
  assign { N33425, N33424, N33423, N33422 } = (N690)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33421)? { N33104, N33105, N33106, N33107 } : 1'b0;
  assign N690 = N33354;
  assign { N33430, N33429, N33428, N33427 } = (N691)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33426)? { N33108, N33109, N33110, N33111 } : 1'b0;
  assign N691 = N33355;
  assign { N33435, N33434, N33433, N33432 } = (N692)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33431)? { N33112, N33113, N33114, N33115 } : 1'b0;
  assign N692 = N33356;
  assign { N33440, N33439, N33438, N33437 } = (N693)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33436)? { N33116, N33117, N33118, N33119 } : 1'b0;
  assign N693 = N33357;
  assign { N33445, N33444, N33443, N33442 } = (N694)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33441)? { N33120, N33121, N33122, N33123 } : 1'b0;
  assign N694 = N33358;
  assign { N33450, N33449, N33448, N33447 } = (N695)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33446)? { N33124, N33125, N33126, N33127 } : 1'b0;
  assign N695 = N33359;
  assign { N33455, N33454, N33453, N33452 } = (N696)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33451)? { N33128, N33129, N33130, N33131 } : 1'b0;
  assign N696 = N33360;
  assign { N33460, N33459, N33458, N33457 } = (N697)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33456)? { N33132, N33133, N33134, N33135 } : 1'b0;
  assign N697 = N33361;
  assign { N33465, N33464, N33463, N33462 } = (N698)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33461)? { N33136, N33137, N33138, N33139 } : 1'b0;
  assign N698 = N33362;
  assign { N33470, N33469, N33468, N33467 } = (N699)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33466)? { N33140, N33141, N33142, N33143 } : 1'b0;
  assign N699 = N33363;
  assign { N33475, N33474, N33473, N33472 } = (N700)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33471)? { N33144, N33145, N33146, N33147 } : 1'b0;
  assign N700 = N33364;
  assign { N33480, N33479, N33478, N33477 } = (N701)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33476)? { N33148, N33149, N33150, N33151 } : 1'b0;
  assign N701 = N33365;
  assign { N33485, N33484, N33483, N33482 } = (N702)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33481)? { N33152, N33153, N33154, N33155 } : 1'b0;
  assign N702 = N33366;
  assign { N33490, N33489, N33488, N33487 } = (N703)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33486)? { N33156, N33157, N33158, N33159 } : 1'b0;
  assign N703 = N33367;
  assign { N33495, N33494, N33493, N33492 } = (N704)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33491)? { N33160, N33161, N33162, N33163 } : 1'b0;
  assign N704 = N33368;
  assign { N33500, N33499, N33498, N33497 } = (N705)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33496)? { N33164, N33165, N33166, N33167 } : 1'b0;
  assign N705 = N33369;
  assign { N33505, N33504, N33503, N33502 } = (N706)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33501)? { N33168, N33169, N33170, N33171 } : 1'b0;
  assign N706 = N33370;
  assign { N33510, N33509, N33508, N33507 } = (N707)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33506)? { N33172, N33173, N33174, N33175 } : 1'b0;
  assign N707 = N33371;
  assign { N33515, N33514, N33513, N33512 } = (N708)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33511)? { N33176, N33177, N33178, N33179 } : 1'b0;
  assign N708 = N33372;
  assign { N33520, N33519, N33518, N33517 } = (N709)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33516)? { N33180, N33181, N33182, N33183 } : 1'b0;
  assign N709 = N33373;
  assign { N33525, N33524, N33523, N33522 } = (N710)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33521)? { N33184, N33185, N33186, N33187 } : 1'b0;
  assign N710 = N33374;
  assign { N33530, N33529, N33528, N33527 } = (N711)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33526)? { N33188, N33189, N33190, N33191 } : 1'b0;
  assign N711 = N33375;
  assign { N33535, N33534, N33533, N33532 } = (N712)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33531)? { N33192, N33193, N33194, N33195 } : 1'b0;
  assign N712 = N33376;
  assign { N33540, N33539, N33538, N33537 } = (N713)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33536)? { N33196, N33197, N33198, N33199 } : 1'b0;
  assign N713 = N33377;
  assign { N33545, N33544, N33543, N33542 } = (N714)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33541)? { N33200, N33201, N33202, N33203 } : 1'b0;
  assign N714 = N33378;
  assign { N33550, N33549, N33548, N33547 } = (N715)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33546)? { N33204, N33205, N33206, N33207 } : 1'b0;
  assign N715 = N33379;
  assign { N33555, N33554, N33553, N33552 } = (N716)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33551)? { N33208, N33209, N33210, N33211 } : 1'b0;
  assign N716 = N33380;
  assign { N33560, N33559, N33558, N33557 } = (N717)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33556)? { N33212, N33213, N33214, N33215 } : 1'b0;
  assign N717 = N33381;
  assign { N33565, N33564, N33563, N33562 } = (N718)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33561)? { N33216, N33217, N33218, N33219 } : 1'b0;
  assign N718 = N33382;
  assign { N33570, N33569, N33568, N33567 } = (N719)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33566)? { N33220, N33221, N33222, N33223 } : 1'b0;
  assign N719 = N33383;
  assign { N33575, N33574, N33573, N33572 } = (N720)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33571)? { N33224, N33225, N33226, N33227 } : 1'b0;
  assign N720 = N33384;
  assign { N33580, N33579, N33578, N33577 } = (N721)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33576)? { N33228, N33229, N33230, N33231 } : 1'b0;
  assign N721 = N33385;
  assign { N33585, N33584, N33583, N33582 } = (N722)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33581)? { N33232, N33233, N33234, N33235 } : 1'b0;
  assign N722 = N33386;
  assign { N33590, N33589, N33588, N33587 } = (N723)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33586)? { N33236, N33237, N33238, N33239 } : 1'b0;
  assign N723 = N33387;
  assign { N33595, N33594, N33593, N33592 } = (N724)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33591)? { N33240, N33241, N33242, N33243 } : 1'b0;
  assign N724 = N33388;
  assign { N33600, N33599, N33598, N33597 } = (N725)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33596)? { N33244, N33245, N33246, N33247 } : 1'b0;
  assign N725 = N33389;
  assign { N33605, N33604, N33603, N33602 } = (N726)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33601)? { N33248, N33249, N33250, N33251 } : 1'b0;
  assign N726 = N33390;
  assign { N33610, N33609, N33608, N33607 } = (N727)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33606)? { N33252, N33253, N33254, N33255 } : 1'b0;
  assign N727 = N33391;
  assign { N33615, N33614, N33613, N33612 } = (N728)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33611)? { N33256, N33257, N33258, N33259 } : 1'b0;
  assign N728 = N33392;
  assign { N33620, N33619, N33618, N33617 } = (N729)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33616)? { N33260, N33261, N33262, N33263 } : 1'b0;
  assign N729 = N33393;
  assign { N33625, N33624, N33623, N33622 } = (N730)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33621)? { N33264, N33265, N33266, N33267 } : 1'b0;
  assign N730 = N33394;
  assign { N33630, N33629, N33628, N33627 } = (N731)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33626)? { N33268, N33269, N33270, N33271 } : 1'b0;
  assign N731 = N33395;
  assign { N33635, N33634, N33633, N33632 } = (N732)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33631)? { N33272, N33273, N33274, N33275 } : 1'b0;
  assign N732 = N33396;
  assign { N33640, N33639, N33638, N33637 } = (N733)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33636)? { N33276, N33277, N33278, N33279 } : 1'b0;
  assign N733 = N33397;
  assign { N33645, N33644, N33643, N33642 } = (N734)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33641)? { N33280, N33281, N33282, N33283 } : 1'b0;
  assign N734 = N33398;
  assign { N33650, N33649, N33648, N33647 } = (N735)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33646)? { N33284, N33285, N33286, N33287 } : 1'b0;
  assign N735 = N33399;
  assign { N33655, N33654, N33653, N33652 } = (N736)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33651)? { N33288, N33289, N33290, N33291 } : 1'b0;
  assign N736 = N33400;
  assign { N33660, N33659, N33658, N33657 } = (N737)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33656)? { N33292, N33293, N33294, N33295 } : 1'b0;
  assign N737 = N33401;
  assign { N33665, N33664, N33663, N33662 } = (N738)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33661)? { N33296, N33297, N33298, N33299 } : 1'b0;
  assign N738 = N33402;
  assign { N33670, N33669, N33668, N33667 } = (N739)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33666)? { N33300, N33301, N33302, N33303 } : 1'b0;
  assign N739 = N33403;
  assign { N33675, N33674, N33673, N33672 } = (N740)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33671)? { N33304, N33305, N33306, N33307 } : 1'b0;
  assign N740 = N33404;
  assign { N33680, N33679, N33678, N33677 } = (N741)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33676)? { N33308, N33309, N33310, N33311 } : 1'b0;
  assign N741 = N33405;
  assign { N33685, N33684, N33683, N33682 } = (N742)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33681)? { N33312, N33313, N33314, N33315 } : 1'b0;
  assign N742 = N33406;
  assign { N33690, N33689, N33688, N33687 } = (N743)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33686)? { N33316, N33317, N33318, N33319 } : 1'b0;
  assign N743 = N33407;
  assign { N33695, N33694, N33693, N33692 } = (N744)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33691)? { N33320, N33321, N33322, N33323 } : 1'b0;
  assign N744 = N33408;
  assign { N33700, N33699, N33698, N33697 } = (N745)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33696)? { N33324, N33325, N33326, N33327 } : 1'b0;
  assign N745 = N33409;
  assign { N33705, N33704, N33703, N33702 } = (N746)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33701)? { N33328, N33329, N33330, N33331 } : 1'b0;
  assign N746 = N33410;
  assign { N33710, N33709, N33708, N33707 } = (N747)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33706)? { N33332, N33333, N33334, N33335 } : 1'b0;
  assign N747 = N33411;
  assign { N33715, N33714, N33713, N33712 } = (N748)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33711)? { N33336, N33337, N33338, N33339 } : 1'b0;
  assign N748 = N33412;
  assign { N33720, N33719, N33718, N33717 } = (N749)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33716)? { N33340, N33341, N33342, N33343 } : 1'b0;
  assign N749 = N33413;
  assign { N33725, N33724, N33723, N33722 } = (N750)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33721)? { N33344, N33345, N33346, N33347 } : 1'b0;
  assign N750 = N33414;
  assign { N33730, N33729, N33728, N33727 } = (N751)? { mem_q[2832:2832], mem_q[2833:2833], mem_q[2834:2834], mem_q[2835:2835] } : 
                                              (N33726)? { N33348, N33349, N33350, N33351 } : 1'b0;
  assign N751 = N33415;
  assign rd_clobber_gpr_o[255:4] = (N752)? { N33727, N33728, N33729, N33730, N33722, N33723, N33724, N33725, N33717, N33718, N33719, N33720, N33712, N33713, N33714, N33715, N33707, N33708, N33709, N33710, N33702, N33703, N33704, N33705, N33697, N33698, N33699, N33700, N33692, N33693, N33694, N33695, N33687, N33688, N33689, N33690, N33682, N33683, N33684, N33685, N33677, N33678, N33679, N33680, N33672, N33673, N33674, N33675, N33667, N33668, N33669, N33670, N33662, N33663, N33664, N33665, N33657, N33658, N33659, N33660, N33652, N33653, N33654, N33655, N33647, N33648, N33649, N33650, N33642, N33643, N33644, N33645, N33637, N33638, N33639, N33640, N33632, N33633, N33634, N33635, N33627, N33628, N33629, N33630, N33622, N33623, N33624, N33625, N33617, N33618, N33619, N33620, N33612, N33613, N33614, N33615, N33607, N33608, N33609, N33610, N33602, N33603, N33604, N33605, N33597, N33598, N33599, N33600, N33592, N33593, N33594, N33595, N33587, N33588, N33589, N33590, N33582, N33583, N33584, N33585, N33577, N33578, N33579, N33580, N33572, N33573, N33574, N33575, N33567, N33568, N33569, N33570, N33562, N33563, N33564, N33565, N33557, N33558, N33559, N33560, N33552, N33553, N33554, N33555, N33547, N33548, N33549, N33550, N33542, N33543, N33544, N33545, N33537, N33538, N33539, N33540, N33532, N33533, N33534, N33535, N33527, N33528, N33529, N33530, N33522, N33523, N33524, N33525, N33517, N33518, N33519, N33520, N33512, N33513, N33514, N33515, N33507, N33508, N33509, N33510, N33502, N33503, N33504, N33505, N33497, N33498, N33499, N33500, N33492, N33493, N33494, N33495, N33487, N33488, N33489, N33490, N33482, N33483, N33484, N33485, N33477, N33478, N33479, N33480, N33472, N33473, N33474, N33475, N33467, N33468, N33469, N33470, N33462, N33463, N33464, N33465, N33457, N33458, N33459, N33460, N33452, N33453, N33454, N33455, N33447, N33448, N33449, N33450, N33442, N33443, N33444, N33445, N33437, N33438, N33439, N33440, N33432, N33433, N33434, N33435, N33427, N33428, N33429, N33430, N33422, N33423, N33424, N33425, N33417, N33418, N33419, N33420 } : 
                                   (N33352)? { N33351, N33350, N33349, N33348, N33347, N33346, N33345, N33344, N33343, N33342, N33341, N33340, N33339, N33338, N33337, N33336, N33335, N33334, N33333, N33332, N33331, N33330, N33329, N33328, N33327, N33326, N33325, N33324, N33323, N33322, N33321, N33320, N33319, N33318, N33317, N33316, N33315, N33314, N33313, N33312, N33311, N33310, N33309, N33308, N33307, N33306, N33305, N33304, N33303, N33302, N33301, N33300, N33299, N33298, N33297, N33296, N33295, N33294, N33293, N33292, N33291, N33290, N33289, N33288, N33287, N33286, N33285, N33284, N33283, N33282, N33281, N33280, N33279, N33278, N33277, N33276, N33275, N33274, N33273, N33272, N33271, N33270, N33269, N33268, N33267, N33266, N33265, N33264, N33263, N33262, N33261, N33260, N33259, N33258, N33257, N33256, N33255, N33254, N33253, N33252, N33251, N33250, N33249, N33248, N33247, N33246, N33245, N33244, N33243, N33242, N33241, N33240, N33239, N33238, N33237, N33236, N33235, N33234, N33233, N33232, N33231, N33230, N33229, N33228, N33227, N33226, N33225, N33224, N33223, N33222, N33221, N33220, N33219, N33218, N33217, N33216, N33215, N33214, N33213, N33212, N33211, N33210, N33209, N33208, N33207, N33206, N33205, N33204, N33203, N33202, N33201, N33200, N33199, N33198, N33197, N33196, N33195, N33194, N33193, N33192, N33191, N33190, N33189, N33188, N33187, N33186, N33185, N33184, N33183, N33182, N33181, N33180, N33179, N33178, N33177, N33176, N33175, N33174, N33173, N33172, N33171, N33170, N33169, N33168, N33167, N33166, N33165, N33164, N33163, N33162, N33161, N33160, N33159, N33158, N33157, N33156, N33155, N33154, N33153, N33152, N33151, N33150, N33149, N33148, N33147, N33146, N33145, N33144, N33143, N33142, N33141, N33140, N33139, N33138, N33137, N33136, N33135, N33134, N33133, N33132, N33131, N33130, N33129, N33128, N33127, N33126, N33125, N33124, N33123, N33122, N33121, N33120, N33119, N33118, N33117, N33116, N33115, N33114, N33113, N33112, N33111, N33110, N33109, N33108, N33107, N33106, N33105, N33104, N33103, N33102, N33101, N33100 } : 1'b0;
  assign N752 = mem_q[2903];
  assign { N33740, N33739 } = (N753)? mem_q[203:202] : 
                              (N754)? { 1'b0, 1'b0 } : 1'b0;
  assign N753 = N33737;
  assign N754 = N33738;
  assign N33741 = (N753)? mem_q[201] : 
                  (N754)? 1'b0 : 1'b0;
  assign { N33805, N33804, N33803, N33802, N33801, N33800, N33799, N33798, N33797, N33796, N33795, N33794, N33793, N33792, N33791, N33790, N33789, N33788, N33787, N33786, N33785, N33784, N33783, N33782, N33781, N33780, N33779, N33778, N33777, N33776, N33775, N33774, N33773, N33772, N33771, N33770, N33769, N33768, N33767, N33766, N33765, N33764, N33763, N33762, N33761, N33760, N33759, N33758, N33757, N33756, N33755, N33754, N33753, N33752, N33751, N33750, N33749, N33748, N33747, N33746, N33745, N33744, N33743, N33742 } = (N755)? mem_q[265:202] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N756)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N755 = N33735;
  assign N756 = N33736;
  assign N33806 = (N755)? mem_q[201] : 
                  (N756)? 1'b0 : 1'b0;
  assign { N33808, N33807 } = (N755)? { 1'b0, 1'b0 } : 
                              (N756)? { N33740, N33739 } : 1'b0;
  assign N33809 = (N755)? 1'b0 : 
                  (N756)? N33741 : 1'b0;
  assign { N33873, N33872, N33871, N33870, N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, N33861, N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, N33852, N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, N33843, N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, N33834, N33833, N33832, N33831, N33830, N33829, N33828, N33827, N33826, N33825, N33824, N33823, N33822, N33821, N33820, N33819, N33818, N33817, N33816, N33815, N33814, N33813, N33812, N33811, N33810 } = (N757)? mem_q[265:202] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N758)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N757 = N33732;
  assign N758 = N33733;
  assign N33874 = (N757)? mem_q[201] : 
                  (N758)? 1'b0 : 1'b0;
  assign { N33876, N33875 } = (N757)? { 1'b0, 1'b0 } : 
                              (N758)? { N33808, N33807 } : 1'b0;
  assign N33877 = (N757)? 1'b0 : 
                  (N758)? N33809 : 1'b0;
  assign { N33941, N33940, N33939, N33938, N33937, N33936, N33935, N33934, N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, N33925, N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, N33916, N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, N33907, N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, N33898, N33897, N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, N33888, N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, N33879, N33878 } = (N757)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N758)? { N33805, N33804, N33803, N33802, N33801, N33800, N33799, N33798, N33797, N33796, N33795, N33794, N33793, N33792, N33791, N33790, N33789, N33788, N33787, N33786, N33785, N33784, N33783, N33782, N33781, N33780, N33779, N33778, N33777, N33776, N33775, N33774, N33773, N33772, N33771, N33770, N33769, N33768, N33767, N33766, N33765, N33764, N33763, N33762, N33761, N33760, N33759, N33758, N33757, N33756, N33755, N33754, N33753, N33752, N33751, N33750, N33749, N33748, N33747, N33746, N33745, N33744, N33743, N33742 } : 1'b0;
  assign N33942 = (N757)? 1'b0 : 
                  (N758)? N33806 : 1'b0;
  assign { N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962, N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, N33943 } = (N304)? { N33941, N33940, N33939, N33938, N33937, N33936, N33935, N33934, N33933, N33932, N33931, N33930, N33929, N33928, N33927, N33926, N33925, N33924, N33923, N33922, N33921, N33920, N33919, N33918, N33917, N33916, N33915, N33914, N33913, N33912, N33911, N33910, N33909, N33908, N33907, N33906, N33905, N33904, N33903, N33902, N33901, N33900, N33899, N33898, N33897, N33896, N33895, N33894, N33893, N33892, N33891, N33890, N33889, N33888, N33887, N33886, N33885, N33884, N33883, N33882, N33881, N33880, N33879, N33878 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N28935)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34007 = (N304)? N33942 : 
                  (N28935)? 1'b0 : 1'b0;
  assign { N34071, N34070, N34069, N34068, N34067, N34066, N34065, N34064, N34063, N34062, N34061, N34060, N34059, N34058, N34057, N34056, N34055, N34054, N34053, N34052, N34051, N34050, N34049, N34048, N34047, N34046, N34045, N34044, N34043, N34042, N34041, N34040, N34039, N34038, N34037, N34036, N34035, N34034, N34033, N34032, N34031, N34030, N34029, N34028, N34027, N34026, N34025, N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008 } = (N304)? { N33873, N33872, N33871, N33870, N33869, N33868, N33867, N33866, N33865, N33864, N33863, N33862, N33861, N33860, N33859, N33858, N33857, N33856, N33855, N33854, N33853, N33852, N33851, N33850, N33849, N33848, N33847, N33846, N33845, N33844, N33843, N33842, N33841, N33840, N33839, N33838, N33837, N33836, N33835, N33834, N33833, N33832, N33831, N33830, N33829, N33828, N33827, N33826, N33825, N33824, N33823, N33822, N33821, N33820, N33819, N33818, N33817, N33816, N33815, N33814, N33813, N33812, N33811, N33810 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N28935)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34072 = (N304)? N33874 : 
                  (N28935)? 1'b0 : 1'b0;
  assign { N34074, N34073 } = (N304)? { N33876, N33875 } : 
                              (N28935)? { 1'b0, 1'b0 } : 1'b0;
  assign N34075 = (N304)? N33877 : 
                  (N28935)? 1'b0 : 1'b0;
  assign { N34085, N34084 } = (N759)? mem_q[566:565] : 
                              (N760)? { N34074, N34073 } : 1'b0;
  assign N759 = N34082;
  assign N760 = N34083;
  assign N34086 = (N759)? mem_q[564] : 
                  (N760)? N34075 : 1'b0;
  assign { N34150, N34149, N34148, N34147, N34146, N34145, N34144, N34143, N34142, N34141, N34140, N34139, N34138, N34137, N34136, N34135, N34134, N34133, N34132, N34131, N34130, N34129, N34128, N34127, N34126, N34125, N34124, N34123, N34122, N34121, N34120, N34119, N34118, N34117, N34116, N34115, N34114, N34113, N34112, N34111, N34110, N34109, N34108, N34107, N34106, N34105, N34104, N34103, N34102, N34101, N34100, N34099, N34098, N34097, N34096, N34095, N34094, N34093, N34092, N34091, N34090, N34089, N34088, N34087 } = (N761)? mem_q[628:565] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N762)? { N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962, N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, N33943 } : 1'b0;
  assign N761 = N34080;
  assign N762 = N34081;
  assign N34151 = (N761)? mem_q[564] : 
                  (N762)? N34007 : 1'b0;
  assign { N34153, N34152 } = (N761)? { N34074, N34073 } : 
                              (N762)? { N34085, N34084 } : 1'b0;
  assign N34154 = (N761)? N34075 : 
                  (N762)? N34086 : 1'b0;
  assign { N34218, N34217, N34216, N34215, N34214, N34213, N34212, N34211, N34210, N34209, N34208, N34207, N34206, N34205, N34204, N34203, N34202, N34201, N34200, N34199, N34198, N34197, N34196, N34195, N34194, N34193, N34192, N34191, N34190, N34189, N34188, N34187, N34186, N34185, N34184, N34183, N34182, N34181, N34180, N34179, N34178, N34177, N34176, N34175, N34174, N34173, N34172, N34171, N34170, N34169, N34168, N34167, N34166, N34165, N34164, N34163, N34162, N34161, N34160, N34159, N34158, N34157, N34156, N34155 } = (N763)? mem_q[628:565] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N764)? { N34071, N34070, N34069, N34068, N34067, N34066, N34065, N34064, N34063, N34062, N34061, N34060, N34059, N34058, N34057, N34056, N34055, N34054, N34053, N34052, N34051, N34050, N34049, N34048, N34047, N34046, N34045, N34044, N34043, N34042, N34041, N34040, N34039, N34038, N34037, N34036, N34035, N34034, N34033, N34032, N34031, N34030, N34029, N34028, N34027, N34026, N34025, N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008 } : 1'b0;
  assign N763 = N34077;
  assign N764 = N34078;
  assign N34219 = (N763)? mem_q[564] : 
                  (N764)? N34072 : 1'b0;
  assign { N34221, N34220 } = (N763)? { N34074, N34073 } : 
                              (N764)? { N34153, N34152 } : 1'b0;
  assign N34222 = (N763)? N34075 : 
                  (N764)? N34154 : 1'b0;
  assign { N34286, N34285, N34284, N34283, N34282, N34281, N34280, N34279, N34278, N34277, N34276, N34275, N34274, N34273, N34272, N34271, N34270, N34269, N34268, N34267, N34266, N34265, N34264, N34263, N34262, N34261, N34260, N34259, N34258, N34257, N34256, N34255, N34254, N34253, N34252, N34251, N34250, N34249, N34248, N34247, N34246, N34245, N34244, N34243, N34242, N34241, N34240, N34239, N34238, N34237, N34236, N34235, N34234, N34233, N34232, N34231, N34230, N34229, N34228, N34227, N34226, N34225, N34224, N34223 } = (N763)? { N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962, N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, N33943 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N764)? { N34150, N34149, N34148, N34147, N34146, N34145, N34144, N34143, N34142, N34141, N34140, N34139, N34138, N34137, N34136, N34135, N34134, N34133, N34132, N34131, N34130, N34129, N34128, N34127, N34126, N34125, N34124, N34123, N34122, N34121, N34120, N34119, N34118, N34117, N34116, N34115, N34114, N34113, N34112, N34111, N34110, N34109, N34108, N34107, N34106, N34105, N34104, N34103, N34102, N34101, N34100, N34099, N34098, N34097, N34096, N34095, N34094, N34093, N34092, N34091, N34090, N34089, N34088, N34087 } : 1'b0;
  assign N34287 = (N763)? N34007 : 
                  (N764)? N34151 : 1'b0;
  assign { N34351, N34350, N34349, N34348, N34347, N34346, N34345, N34344, N34343, N34342, N34341, N34340, N34339, N34338, N34337, N34336, N34335, N34334, N34333, N34332, N34331, N34330, N34329, N34328, N34327, N34326, N34325, N34324, N34323, N34322, N34321, N34320, N34319, N34318, N34317, N34316, N34315, N34314, N34313, N34312, N34311, N34310, N34309, N34308, N34307, N34306, N34305, N34304, N34303, N34302, N34301, N34300, N34299, N34298, N34297, N34296, N34295, N34294, N34293, N34292, N34291, N34290, N34289, N34288 } = (N368)? { N34286, N34285, N34284, N34283, N34282, N34281, N34280, N34279, N34278, N34277, N34276, N34275, N34274, N34273, N34272, N34271, N34270, N34269, N34268, N34267, N34266, N34265, N34264, N34263, N34262, N34261, N34260, N34259, N34258, N34257, N34256, N34255, N34254, N34253, N34252, N34251, N34250, N34249, N34248, N34247, N34246, N34245, N34244, N34243, N34242, N34241, N34240, N34239, N34238, N34237, N34236, N34235, N34234, N34233, N34232, N34231, N34230, N34229, N34228, N34227, N34226, N34225, N34224, N34223 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N29566)? { N34006, N34005, N34004, N34003, N34002, N34001, N34000, N33999, N33998, N33997, N33996, N33995, N33994, N33993, N33992, N33991, N33990, N33989, N33988, N33987, N33986, N33985, N33984, N33983, N33982, N33981, N33980, N33979, N33978, N33977, N33976, N33975, N33974, N33973, N33972, N33971, N33970, N33969, N33968, N33967, N33966, N33965, N33964, N33963, N33962, N33961, N33960, N33959, N33958, N33957, N33956, N33955, N33954, N33953, N33952, N33951, N33950, N33949, N33948, N33947, N33946, N33945, N33944, N33943 } : 1'b0;
  assign N34352 = (N368)? N34287 : 
                  (N29566)? N34007 : 1'b0;
  assign { N34416, N34415, N34414, N34413, N34412, N34411, N34410, N34409, N34408, N34407, N34406, N34405, N34404, N34403, N34402, N34401, N34400, N34399, N34398, N34397, N34396, N34395, N34394, N34393, N34392, N34391, N34390, N34389, N34388, N34387, N34386, N34385, N34384, N34383, N34382, N34381, N34380, N34379, N34378, N34377, N34376, N34375, N34374, N34373, N34372, N34371, N34370, N34369, N34368, N34367, N34366, N34365, N34364, N34363, N34362, N34361, N34360, N34359, N34358, N34357, N34356, N34355, N34354, N34353 } = (N368)? { N34218, N34217, N34216, N34215, N34214, N34213, N34212, N34211, N34210, N34209, N34208, N34207, N34206, N34205, N34204, N34203, N34202, N34201, N34200, N34199, N34198, N34197, N34196, N34195, N34194, N34193, N34192, N34191, N34190, N34189, N34188, N34187, N34186, N34185, N34184, N34183, N34182, N34181, N34180, N34179, N34178, N34177, N34176, N34175, N34174, N34173, N34172, N34171, N34170, N34169, N34168, N34167, N34166, N34165, N34164, N34163, N34162, N34161, N34160, N34159, N34158, N34157, N34156, N34155 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N29566)? { N34071, N34070, N34069, N34068, N34067, N34066, N34065, N34064, N34063, N34062, N34061, N34060, N34059, N34058, N34057, N34056, N34055, N34054, N34053, N34052, N34051, N34050, N34049, N34048, N34047, N34046, N34045, N34044, N34043, N34042, N34041, N34040, N34039, N34038, N34037, N34036, N34035, N34034, N34033, N34032, N34031, N34030, N34029, N34028, N34027, N34026, N34025, N34024, N34023, N34022, N34021, N34020, N34019, N34018, N34017, N34016, N34015, N34014, N34013, N34012, N34011, N34010, N34009, N34008 } : 1'b0;
  assign N34417 = (N368)? N34219 : 
                  (N29566)? N34072 : 1'b0;
  assign { N34419, N34418 } = (N368)? { N34221, N34220 } : 
                              (N29566)? { N34074, N34073 } : 1'b0;
  assign N34420 = (N368)? N34222 : 
                  (N29566)? N34075 : 1'b0;
  assign { N34430, N34429 } = (N765)? mem_q[929:928] : 
                              (N766)? { N34419, N34418 } : 1'b0;
  assign N765 = N34427;
  assign N766 = N34428;
  assign N34431 = (N765)? mem_q[927] : 
                  (N766)? N34420 : 1'b0;
  assign { N34495, N34494, N34493, N34492, N34491, N34490, N34489, N34488, N34487, N34486, N34485, N34484, N34483, N34482, N34481, N34480, N34479, N34478, N34477, N34476, N34475, N34474, N34473, N34472, N34471, N34470, N34469, N34468, N34467, N34466, N34465, N34464, N34463, N34462, N34461, N34460, N34459, N34458, N34457, N34456, N34455, N34454, N34453, N34452, N34451, N34450, N34449, N34448, N34447, N34446, N34445, N34444, N34443, N34442, N34441, N34440, N34439, N34438, N34437, N34436, N34435, N34434, N34433, N34432 } = (N767)? mem_q[991:928] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N768)? { N34351, N34350, N34349, N34348, N34347, N34346, N34345, N34344, N34343, N34342, N34341, N34340, N34339, N34338, N34337, N34336, N34335, N34334, N34333, N34332, N34331, N34330, N34329, N34328, N34327, N34326, N34325, N34324, N34323, N34322, N34321, N34320, N34319, N34318, N34317, N34316, N34315, N34314, N34313, N34312, N34311, N34310, N34309, N34308, N34307, N34306, N34305, N34304, N34303, N34302, N34301, N34300, N34299, N34298, N34297, N34296, N34295, N34294, N34293, N34292, N34291, N34290, N34289, N34288 } : 1'b0;
  assign N767 = N34425;
  assign N768 = N34426;
  assign N34496 = (N767)? mem_q[927] : 
                  (N768)? N34352 : 1'b0;
  assign { N34498, N34497 } = (N767)? { N34419, N34418 } : 
                              (N768)? { N34430, N34429 } : 1'b0;
  assign N34499 = (N767)? N34420 : 
                  (N768)? N34431 : 1'b0;
  assign { N34563, N34562, N34561, N34560, N34559, N34558, N34557, N34556, N34555, N34554, N34553, N34552, N34551, N34550, N34549, N34548, N34547, N34546, N34545, N34544, N34543, N34542, N34541, N34540, N34539, N34538, N34537, N34536, N34535, N34534, N34533, N34532, N34531, N34530, N34529, N34528, N34527, N34526, N34525, N34524, N34523, N34522, N34521, N34520, N34519, N34518, N34517, N34516, N34515, N34514, N34513, N34512, N34511, N34510, N34509, N34508, N34507, N34506, N34505, N34504, N34503, N34502, N34501, N34500 } = (N769)? mem_q[991:928] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N770)? { N34416, N34415, N34414, N34413, N34412, N34411, N34410, N34409, N34408, N34407, N34406, N34405, N34404, N34403, N34402, N34401, N34400, N34399, N34398, N34397, N34396, N34395, N34394, N34393, N34392, N34391, N34390, N34389, N34388, N34387, N34386, N34385, N34384, N34383, N34382, N34381, N34380, N34379, N34378, N34377, N34376, N34375, N34374, N34373, N34372, N34371, N34370, N34369, N34368, N34367, N34366, N34365, N34364, N34363, N34362, N34361, N34360, N34359, N34358, N34357, N34356, N34355, N34354, N34353 } : 1'b0;
  assign N769 = N34422;
  assign N770 = N34423;
  assign N34564 = (N769)? mem_q[927] : 
                  (N770)? N34417 : 1'b0;
  assign { N34566, N34565 } = (N769)? { N34419, N34418 } : 
                              (N770)? { N34498, N34497 } : 1'b0;
  assign N34567 = (N769)? N34420 : 
                  (N770)? N34499 : 1'b0;
  assign { N34631, N34630, N34629, N34628, N34627, N34626, N34625, N34624, N34623, N34622, N34621, N34620, N34619, N34618, N34617, N34616, N34615, N34614, N34613, N34612, N34611, N34610, N34609, N34608, N34607, N34606, N34605, N34604, N34603, N34602, N34601, N34600, N34599, N34598, N34597, N34596, N34595, N34594, N34593, N34592, N34591, N34590, N34589, N34588, N34587, N34586, N34585, N34584, N34583, N34582, N34581, N34580, N34579, N34578, N34577, N34576, N34575, N34574, N34573, N34572, N34571, N34570, N34569, N34568 } = (N769)? { N34351, N34350, N34349, N34348, N34347, N34346, N34345, N34344, N34343, N34342, N34341, N34340, N34339, N34338, N34337, N34336, N34335, N34334, N34333, N34332, N34331, N34330, N34329, N34328, N34327, N34326, N34325, N34324, N34323, N34322, N34321, N34320, N34319, N34318, N34317, N34316, N34315, N34314, N34313, N34312, N34311, N34310, N34309, N34308, N34307, N34306, N34305, N34304, N34303, N34302, N34301, N34300, N34299, N34298, N34297, N34296, N34295, N34294, N34293, N34292, N34291, N34290, N34289, N34288 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N770)? { N34495, N34494, N34493, N34492, N34491, N34490, N34489, N34488, N34487, N34486, N34485, N34484, N34483, N34482, N34481, N34480, N34479, N34478, N34477, N34476, N34475, N34474, N34473, N34472, N34471, N34470, N34469, N34468, N34467, N34466, N34465, N34464, N34463, N34462, N34461, N34460, N34459, N34458, N34457, N34456, N34455, N34454, N34453, N34452, N34451, N34450, N34449, N34448, N34447, N34446, N34445, N34444, N34443, N34442, N34441, N34440, N34439, N34438, N34437, N34436, N34435, N34434, N34433, N34432 } : 1'b0;
  assign N34632 = (N769)? N34352 : 
                  (N770)? N34496 : 1'b0;
  assign { N34696, N34695, N34694, N34693, N34692, N34691, N34690, N34689, N34688, N34687, N34686, N34685, N34684, N34683, N34682, N34681, N34680, N34679, N34678, N34677, N34676, N34675, N34674, N34673, N34672, N34671, N34670, N34669, N34668, N34667, N34666, N34665, N34664, N34663, N34662, N34661, N34660, N34659, N34658, N34657, N34656, N34655, N34654, N34653, N34652, N34651, N34650, N34649, N34648, N34647, N34646, N34645, N34644, N34643, N34642, N34641, N34640, N34639, N34638, N34637, N34636, N34635, N34634, N34633 } = (N432)? { N34631, N34630, N34629, N34628, N34627, N34626, N34625, N34624, N34623, N34622, N34621, N34620, N34619, N34618, N34617, N34616, N34615, N34614, N34613, N34612, N34611, N34610, N34609, N34608, N34607, N34606, N34605, N34604, N34603, N34602, N34601, N34600, N34599, N34598, N34597, N34596, N34595, N34594, N34593, N34592, N34591, N34590, N34589, N34588, N34587, N34586, N34585, N34584, N34583, N34582, N34581, N34580, N34579, N34578, N34577, N34576, N34575, N34574, N34573, N34572, N34571, N34570, N34569, N34568 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N30197)? { N34351, N34350, N34349, N34348, N34347, N34346, N34345, N34344, N34343, N34342, N34341, N34340, N34339, N34338, N34337, N34336, N34335, N34334, N34333, N34332, N34331, N34330, N34329, N34328, N34327, N34326, N34325, N34324, N34323, N34322, N34321, N34320, N34319, N34318, N34317, N34316, N34315, N34314, N34313, N34312, N34311, N34310, N34309, N34308, N34307, N34306, N34305, N34304, N34303, N34302, N34301, N34300, N34299, N34298, N34297, N34296, N34295, N34294, N34293, N34292, N34291, N34290, N34289, N34288 } : 1'b0;
  assign N34697 = (N432)? N34632 : 
                  (N30197)? N34352 : 1'b0;
  assign { N34761, N34760, N34759, N34758, N34757, N34756, N34755, N34754, N34753, N34752, N34751, N34750, N34749, N34748, N34747, N34746, N34745, N34744, N34743, N34742, N34741, N34740, N34739, N34738, N34737, N34736, N34735, N34734, N34733, N34732, N34731, N34730, N34729, N34728, N34727, N34726, N34725, N34724, N34723, N34722, N34721, N34720, N34719, N34718, N34717, N34716, N34715, N34714, N34713, N34712, N34711, N34710, N34709, N34708, N34707, N34706, N34705, N34704, N34703, N34702, N34701, N34700, N34699, N34698 } = (N432)? { N34563, N34562, N34561, N34560, N34559, N34558, N34557, N34556, N34555, N34554, N34553, N34552, N34551, N34550, N34549, N34548, N34547, N34546, N34545, N34544, N34543, N34542, N34541, N34540, N34539, N34538, N34537, N34536, N34535, N34534, N34533, N34532, N34531, N34530, N34529, N34528, N34527, N34526, N34525, N34524, N34523, N34522, N34521, N34520, N34519, N34518, N34517, N34516, N34515, N34514, N34513, N34512, N34511, N34510, N34509, N34508, N34507, N34506, N34505, N34504, N34503, N34502, N34501, N34500 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N30197)? { N34416, N34415, N34414, N34413, N34412, N34411, N34410, N34409, N34408, N34407, N34406, N34405, N34404, N34403, N34402, N34401, N34400, N34399, N34398, N34397, N34396, N34395, N34394, N34393, N34392, N34391, N34390, N34389, N34388, N34387, N34386, N34385, N34384, N34383, N34382, N34381, N34380, N34379, N34378, N34377, N34376, N34375, N34374, N34373, N34372, N34371, N34370, N34369, N34368, N34367, N34366, N34365, N34364, N34363, N34362, N34361, N34360, N34359, N34358, N34357, N34356, N34355, N34354, N34353 } : 1'b0;
  assign N34762 = (N432)? N34564 : 
                  (N30197)? N34417 : 1'b0;
  assign { N34764, N34763 } = (N432)? { N34566, N34565 } : 
                              (N30197)? { N34419, N34418 } : 1'b0;
  assign N34765 = (N432)? N34567 : 
                  (N30197)? N34420 : 1'b0;
  assign { N34775, N34774 } = (N771)? mem_q[1292:1291] : 
                              (N772)? { N34764, N34763 } : 1'b0;
  assign N771 = N34772;
  assign N772 = N34773;
  assign N34776 = (N771)? mem_q[1290] : 
                  (N772)? N34765 : 1'b0;
  assign { N34840, N34839, N34838, N34837, N34836, N34835, N34834, N34833, N34832, N34831, N34830, N34829, N34828, N34827, N34826, N34825, N34824, N34823, N34822, N34821, N34820, N34819, N34818, N34817, N34816, N34815, N34814, N34813, N34812, N34811, N34810, N34809, N34808, N34807, N34806, N34805, N34804, N34803, N34802, N34801, N34800, N34799, N34798, N34797, N34796, N34795, N34794, N34793, N34792, N34791, N34790, N34789, N34788, N34787, N34786, N34785, N34784, N34783, N34782, N34781, N34780, N34779, N34778, N34777 } = (N773)? mem_q[1354:1291] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N774)? { N34696, N34695, N34694, N34693, N34692, N34691, N34690, N34689, N34688, N34687, N34686, N34685, N34684, N34683, N34682, N34681, N34680, N34679, N34678, N34677, N34676, N34675, N34674, N34673, N34672, N34671, N34670, N34669, N34668, N34667, N34666, N34665, N34664, N34663, N34662, N34661, N34660, N34659, N34658, N34657, N34656, N34655, N34654, N34653, N34652, N34651, N34650, N34649, N34648, N34647, N34646, N34645, N34644, N34643, N34642, N34641, N34640, N34639, N34638, N34637, N34636, N34635, N34634, N34633 } : 1'b0;
  assign N773 = N34770;
  assign N774 = N34771;
  assign N34841 = (N773)? mem_q[1290] : 
                  (N774)? N34697 : 1'b0;
  assign { N34843, N34842 } = (N773)? { N34764, N34763 } : 
                              (N774)? { N34775, N34774 } : 1'b0;
  assign N34844 = (N773)? N34765 : 
                  (N774)? N34776 : 1'b0;
  assign { N34908, N34907, N34906, N34905, N34904, N34903, N34902, N34901, N34900, N34899, N34898, N34897, N34896, N34895, N34894, N34893, N34892, N34891, N34890, N34889, N34888, N34887, N34886, N34885, N34884, N34883, N34882, N34881, N34880, N34879, N34878, N34877, N34876, N34875, N34874, N34873, N34872, N34871, N34870, N34869, N34868, N34867, N34866, N34865, N34864, N34863, N34862, N34861, N34860, N34859, N34858, N34857, N34856, N34855, N34854, N34853, N34852, N34851, N34850, N34849, N34848, N34847, N34846, N34845 } = (N775)? mem_q[1354:1291] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N776)? { N34761, N34760, N34759, N34758, N34757, N34756, N34755, N34754, N34753, N34752, N34751, N34750, N34749, N34748, N34747, N34746, N34745, N34744, N34743, N34742, N34741, N34740, N34739, N34738, N34737, N34736, N34735, N34734, N34733, N34732, N34731, N34730, N34729, N34728, N34727, N34726, N34725, N34724, N34723, N34722, N34721, N34720, N34719, N34718, N34717, N34716, N34715, N34714, N34713, N34712, N34711, N34710, N34709, N34708, N34707, N34706, N34705, N34704, N34703, N34702, N34701, N34700, N34699, N34698 } : 1'b0;
  assign N775 = N34767;
  assign N776 = N34768;
  assign N34909 = (N775)? mem_q[1290] : 
                  (N776)? N34762 : 1'b0;
  assign { N34911, N34910 } = (N775)? { N34764, N34763 } : 
                              (N776)? { N34843, N34842 } : 1'b0;
  assign N34912 = (N775)? N34765 : 
                  (N776)? N34844 : 1'b0;
  assign { N34976, N34975, N34974, N34973, N34972, N34971, N34970, N34969, N34968, N34967, N34966, N34965, N34964, N34963, N34962, N34961, N34960, N34959, N34958, N34957, N34956, N34955, N34954, N34953, N34952, N34951, N34950, N34949, N34948, N34947, N34946, N34945, N34944, N34943, N34942, N34941, N34940, N34939, N34938, N34937, N34936, N34935, N34934, N34933, N34932, N34931, N34930, N34929, N34928, N34927, N34926, N34925, N34924, N34923, N34922, N34921, N34920, N34919, N34918, N34917, N34916, N34915, N34914, N34913 } = (N775)? { N34696, N34695, N34694, N34693, N34692, N34691, N34690, N34689, N34688, N34687, N34686, N34685, N34684, N34683, N34682, N34681, N34680, N34679, N34678, N34677, N34676, N34675, N34674, N34673, N34672, N34671, N34670, N34669, N34668, N34667, N34666, N34665, N34664, N34663, N34662, N34661, N34660, N34659, N34658, N34657, N34656, N34655, N34654, N34653, N34652, N34651, N34650, N34649, N34648, N34647, N34646, N34645, N34644, N34643, N34642, N34641, N34640, N34639, N34638, N34637, N34636, N34635, N34634, N34633 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N776)? { N34840, N34839, N34838, N34837, N34836, N34835, N34834, N34833, N34832, N34831, N34830, N34829, N34828, N34827, N34826, N34825, N34824, N34823, N34822, N34821, N34820, N34819, N34818, N34817, N34816, N34815, N34814, N34813, N34812, N34811, N34810, N34809, N34808, N34807, N34806, N34805, N34804, N34803, N34802, N34801, N34800, N34799, N34798, N34797, N34796, N34795, N34794, N34793, N34792, N34791, N34790, N34789, N34788, N34787, N34786, N34785, N34784, N34783, N34782, N34781, N34780, N34779, N34778, N34777 } : 1'b0;
  assign N34977 = (N775)? N34697 : 
                  (N776)? N34841 : 1'b0;
  assign { N35041, N35040, N35039, N35038, N35037, N35036, N35035, N35034, N35033, N35032, N35031, N35030, N35029, N35028, N35027, N35026, N35025, N35024, N35023, N35022, N35021, N35020, N35019, N35018, N35017, N35016, N35015, N35014, N35013, N35012, N35011, N35010, N35009, N35008, N35007, N35006, N35005, N35004, N35003, N35002, N35001, N35000, N34999, N34998, N34997, N34996, N34995, N34994, N34993, N34992, N34991, N34990, N34989, N34988, N34987, N34986, N34985, N34984, N34983, N34982, N34981, N34980, N34979, N34978 } = (N496)? { N34976, N34975, N34974, N34973, N34972, N34971, N34970, N34969, N34968, N34967, N34966, N34965, N34964, N34963, N34962, N34961, N34960, N34959, N34958, N34957, N34956, N34955, N34954, N34953, N34952, N34951, N34950, N34949, N34948, N34947, N34946, N34945, N34944, N34943, N34942, N34941, N34940, N34939, N34938, N34937, N34936, N34935, N34934, N34933, N34932, N34931, N34930, N34929, N34928, N34927, N34926, N34925, N34924, N34923, N34922, N34921, N34920, N34919, N34918, N34917, N34916, N34915, N34914, N34913 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N30828)? { N34696, N34695, N34694, N34693, N34692, N34691, N34690, N34689, N34688, N34687, N34686, N34685, N34684, N34683, N34682, N34681, N34680, N34679, N34678, N34677, N34676, N34675, N34674, N34673, N34672, N34671, N34670, N34669, N34668, N34667, N34666, N34665, N34664, N34663, N34662, N34661, N34660, N34659, N34658, N34657, N34656, N34655, N34654, N34653, N34652, N34651, N34650, N34649, N34648, N34647, N34646, N34645, N34644, N34643, N34642, N34641, N34640, N34639, N34638, N34637, N34636, N34635, N34634, N34633 } : 1'b0;
  assign N35042 = (N496)? N34977 : 
                  (N30828)? N34697 : 1'b0;
  assign { N35106, N35105, N35104, N35103, N35102, N35101, N35100, N35099, N35098, N35097, N35096, N35095, N35094, N35093, N35092, N35091, N35090, N35089, N35088, N35087, N35086, N35085, N35084, N35083, N35082, N35081, N35080, N35079, N35078, N35077, N35076, N35075, N35074, N35073, N35072, N35071, N35070, N35069, N35068, N35067, N35066, N35065, N35064, N35063, N35062, N35061, N35060, N35059, N35058, N35057, N35056, N35055, N35054, N35053, N35052, N35051, N35050, N35049, N35048, N35047, N35046, N35045, N35044, N35043 } = (N496)? { N34908, N34907, N34906, N34905, N34904, N34903, N34902, N34901, N34900, N34899, N34898, N34897, N34896, N34895, N34894, N34893, N34892, N34891, N34890, N34889, N34888, N34887, N34886, N34885, N34884, N34883, N34882, N34881, N34880, N34879, N34878, N34877, N34876, N34875, N34874, N34873, N34872, N34871, N34870, N34869, N34868, N34867, N34866, N34865, N34864, N34863, N34862, N34861, N34860, N34859, N34858, N34857, N34856, N34855, N34854, N34853, N34852, N34851, N34850, N34849, N34848, N34847, N34846, N34845 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N30828)? { N34761, N34760, N34759, N34758, N34757, N34756, N34755, N34754, N34753, N34752, N34751, N34750, N34749, N34748, N34747, N34746, N34745, N34744, N34743, N34742, N34741, N34740, N34739, N34738, N34737, N34736, N34735, N34734, N34733, N34732, N34731, N34730, N34729, N34728, N34727, N34726, N34725, N34724, N34723, N34722, N34721, N34720, N34719, N34718, N34717, N34716, N34715, N34714, N34713, N34712, N34711, N34710, N34709, N34708, N34707, N34706, N34705, N34704, N34703, N34702, N34701, N34700, N34699, N34698 } : 1'b0;
  assign N35107 = (N496)? N34909 : 
                  (N30828)? N34762 : 1'b0;
  assign { N35109, N35108 } = (N496)? { N34911, N34910 } : 
                              (N30828)? { N34764, N34763 } : 1'b0;
  assign N35110 = (N496)? N34912 : 
                  (N30828)? N34765 : 1'b0;
  assign { N35120, N35119 } = (N777)? mem_q[1655:1654] : 
                              (N778)? { N35109, N35108 } : 1'b0;
  assign N777 = N35117;
  assign N778 = N35118;
  assign N35121 = (N777)? mem_q[1653] : 
                  (N778)? N35110 : 1'b0;
  assign { N35185, N35184, N35183, N35182, N35181, N35180, N35179, N35178, N35177, N35176, N35175, N35174, N35173, N35172, N35171, N35170, N35169, N35168, N35167, N35166, N35165, N35164, N35163, N35162, N35161, N35160, N35159, N35158, N35157, N35156, N35155, N35154, N35153, N35152, N35151, N35150, N35149, N35148, N35147, N35146, N35145, N35144, N35143, N35142, N35141, N35140, N35139, N35138, N35137, N35136, N35135, N35134, N35133, N35132, N35131, N35130, N35129, N35128, N35127, N35126, N35125, N35124, N35123, N35122 } = (N779)? mem_q[1717:1654] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N780)? { N35041, N35040, N35039, N35038, N35037, N35036, N35035, N35034, N35033, N35032, N35031, N35030, N35029, N35028, N35027, N35026, N35025, N35024, N35023, N35022, N35021, N35020, N35019, N35018, N35017, N35016, N35015, N35014, N35013, N35012, N35011, N35010, N35009, N35008, N35007, N35006, N35005, N35004, N35003, N35002, N35001, N35000, N34999, N34998, N34997, N34996, N34995, N34994, N34993, N34992, N34991, N34990, N34989, N34988, N34987, N34986, N34985, N34984, N34983, N34982, N34981, N34980, N34979, N34978 } : 1'b0;
  assign N779 = N35115;
  assign N780 = N35116;
  assign N35186 = (N779)? mem_q[1653] : 
                  (N780)? N35042 : 1'b0;
  assign { N35188, N35187 } = (N779)? { N35109, N35108 } : 
                              (N780)? { N35120, N35119 } : 1'b0;
  assign N35189 = (N779)? N35110 : 
                  (N780)? N35121 : 1'b0;
  assign { N35253, N35252, N35251, N35250, N35249, N35248, N35247, N35246, N35245, N35244, N35243, N35242, N35241, N35240, N35239, N35238, N35237, N35236, N35235, N35234, N35233, N35232, N35231, N35230, N35229, N35228, N35227, N35226, N35225, N35224, N35223, N35222, N35221, N35220, N35219, N35218, N35217, N35216, N35215, N35214, N35213, N35212, N35211, N35210, N35209, N35208, N35207, N35206, N35205, N35204, N35203, N35202, N35201, N35200, N35199, N35198, N35197, N35196, N35195, N35194, N35193, N35192, N35191, N35190 } = (N781)? mem_q[1717:1654] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N782)? { N35106, N35105, N35104, N35103, N35102, N35101, N35100, N35099, N35098, N35097, N35096, N35095, N35094, N35093, N35092, N35091, N35090, N35089, N35088, N35087, N35086, N35085, N35084, N35083, N35082, N35081, N35080, N35079, N35078, N35077, N35076, N35075, N35074, N35073, N35072, N35071, N35070, N35069, N35068, N35067, N35066, N35065, N35064, N35063, N35062, N35061, N35060, N35059, N35058, N35057, N35056, N35055, N35054, N35053, N35052, N35051, N35050, N35049, N35048, N35047, N35046, N35045, N35044, N35043 } : 1'b0;
  assign N781 = N35112;
  assign N782 = N35113;
  assign N35254 = (N781)? mem_q[1653] : 
                  (N782)? N35107 : 1'b0;
  assign { N35256, N35255 } = (N781)? { N35109, N35108 } : 
                              (N782)? { N35188, N35187 } : 1'b0;
  assign N35257 = (N781)? N35110 : 
                  (N782)? N35189 : 1'b0;
  assign { N35321, N35320, N35319, N35318, N35317, N35316, N35315, N35314, N35313, N35312, N35311, N35310, N35309, N35308, N35307, N35306, N35305, N35304, N35303, N35302, N35301, N35300, N35299, N35298, N35297, N35296, N35295, N35294, N35293, N35292, N35291, N35290, N35289, N35288, N35287, N35286, N35285, N35284, N35283, N35282, N35281, N35280, N35279, N35278, N35277, N35276, N35275, N35274, N35273, N35272, N35271, N35270, N35269, N35268, N35267, N35266, N35265, N35264, N35263, N35262, N35261, N35260, N35259, N35258 } = (N781)? { N35041, N35040, N35039, N35038, N35037, N35036, N35035, N35034, N35033, N35032, N35031, N35030, N35029, N35028, N35027, N35026, N35025, N35024, N35023, N35022, N35021, N35020, N35019, N35018, N35017, N35016, N35015, N35014, N35013, N35012, N35011, N35010, N35009, N35008, N35007, N35006, N35005, N35004, N35003, N35002, N35001, N35000, N34999, N34998, N34997, N34996, N34995, N34994, N34993, N34992, N34991, N34990, N34989, N34988, N34987, N34986, N34985, N34984, N34983, N34982, N34981, N34980, N34979, N34978 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N782)? { N35185, N35184, N35183, N35182, N35181, N35180, N35179, N35178, N35177, N35176, N35175, N35174, N35173, N35172, N35171, N35170, N35169, N35168, N35167, N35166, N35165, N35164, N35163, N35162, N35161, N35160, N35159, N35158, N35157, N35156, N35155, N35154, N35153, N35152, N35151, N35150, N35149, N35148, N35147, N35146, N35145, N35144, N35143, N35142, N35141, N35140, N35139, N35138, N35137, N35136, N35135, N35134, N35133, N35132, N35131, N35130, N35129, N35128, N35127, N35126, N35125, N35124, N35123, N35122 } : 1'b0;
  assign N35322 = (N781)? N35042 : 
                  (N782)? N35186 : 1'b0;
  assign { N35386, N35385, N35384, N35383, N35382, N35381, N35380, N35379, N35378, N35377, N35376, N35375, N35374, N35373, N35372, N35371, N35370, N35369, N35368, N35367, N35366, N35365, N35364, N35363, N35362, N35361, N35360, N35359, N35358, N35357, N35356, N35355, N35354, N35353, N35352, N35351, N35350, N35349, N35348, N35347, N35346, N35345, N35344, N35343, N35342, N35341, N35340, N35339, N35338, N35337, N35336, N35335, N35334, N35333, N35332, N35331, N35330, N35329, N35328, N35327, N35326, N35325, N35324, N35323 } = (N560)? { N35321, N35320, N35319, N35318, N35317, N35316, N35315, N35314, N35313, N35312, N35311, N35310, N35309, N35308, N35307, N35306, N35305, N35304, N35303, N35302, N35301, N35300, N35299, N35298, N35297, N35296, N35295, N35294, N35293, N35292, N35291, N35290, N35289, N35288, N35287, N35286, N35285, N35284, N35283, N35282, N35281, N35280, N35279, N35278, N35277, N35276, N35275, N35274, N35273, N35272, N35271, N35270, N35269, N35268, N35267, N35266, N35265, N35264, N35263, N35262, N35261, N35260, N35259, N35258 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N31459)? { N35041, N35040, N35039, N35038, N35037, N35036, N35035, N35034, N35033, N35032, N35031, N35030, N35029, N35028, N35027, N35026, N35025, N35024, N35023, N35022, N35021, N35020, N35019, N35018, N35017, N35016, N35015, N35014, N35013, N35012, N35011, N35010, N35009, N35008, N35007, N35006, N35005, N35004, N35003, N35002, N35001, N35000, N34999, N34998, N34997, N34996, N34995, N34994, N34993, N34992, N34991, N34990, N34989, N34988, N34987, N34986, N34985, N34984, N34983, N34982, N34981, N34980, N34979, N34978 } : 1'b0;
  assign N35387 = (N560)? N35322 : 
                  (N31459)? N35042 : 1'b0;
  assign { N35451, N35450, N35449, N35448, N35447, N35446, N35445, N35444, N35443, N35442, N35441, N35440, N35439, N35438, N35437, N35436, N35435, N35434, N35433, N35432, N35431, N35430, N35429, N35428, N35427, N35426, N35425, N35424, N35423, N35422, N35421, N35420, N35419, N35418, N35417, N35416, N35415, N35414, N35413, N35412, N35411, N35410, N35409, N35408, N35407, N35406, N35405, N35404, N35403, N35402, N35401, N35400, N35399, N35398, N35397, N35396, N35395, N35394, N35393, N35392, N35391, N35390, N35389, N35388 } = (N560)? { N35253, N35252, N35251, N35250, N35249, N35248, N35247, N35246, N35245, N35244, N35243, N35242, N35241, N35240, N35239, N35238, N35237, N35236, N35235, N35234, N35233, N35232, N35231, N35230, N35229, N35228, N35227, N35226, N35225, N35224, N35223, N35222, N35221, N35220, N35219, N35218, N35217, N35216, N35215, N35214, N35213, N35212, N35211, N35210, N35209, N35208, N35207, N35206, N35205, N35204, N35203, N35202, N35201, N35200, N35199, N35198, N35197, N35196, N35195, N35194, N35193, N35192, N35191, N35190 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N31459)? { N35106, N35105, N35104, N35103, N35102, N35101, N35100, N35099, N35098, N35097, N35096, N35095, N35094, N35093, N35092, N35091, N35090, N35089, N35088, N35087, N35086, N35085, N35084, N35083, N35082, N35081, N35080, N35079, N35078, N35077, N35076, N35075, N35074, N35073, N35072, N35071, N35070, N35069, N35068, N35067, N35066, N35065, N35064, N35063, N35062, N35061, N35060, N35059, N35058, N35057, N35056, N35055, N35054, N35053, N35052, N35051, N35050, N35049, N35048, N35047, N35046, N35045, N35044, N35043 } : 1'b0;
  assign N35452 = (N560)? N35254 : 
                  (N31459)? N35107 : 1'b0;
  assign { N35454, N35453 } = (N560)? { N35256, N35255 } : 
                              (N31459)? { N35109, N35108 } : 1'b0;
  assign N35455 = (N560)? N35257 : 
                  (N31459)? N35110 : 1'b0;
  assign { N35465, N35464 } = (N783)? mem_q[2018:2017] : 
                              (N784)? { N35454, N35453 } : 1'b0;
  assign N783 = N35462;
  assign N784 = N35463;
  assign N35466 = (N783)? mem_q[2016] : 
                  (N784)? N35455 : 1'b0;
  assign { N35530, N35529, N35528, N35527, N35526, N35525, N35524, N35523, N35522, N35521, N35520, N35519, N35518, N35517, N35516, N35515, N35514, N35513, N35512, N35511, N35510, N35509, N35508, N35507, N35506, N35505, N35504, N35503, N35502, N35501, N35500, N35499, N35498, N35497, N35496, N35495, N35494, N35493, N35492, N35491, N35490, N35489, N35488, N35487, N35486, N35485, N35484, N35483, N35482, N35481, N35480, N35479, N35478, N35477, N35476, N35475, N35474, N35473, N35472, N35471, N35470, N35469, N35468, N35467 } = (N785)? mem_q[2080:2017] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N786)? { N35386, N35385, N35384, N35383, N35382, N35381, N35380, N35379, N35378, N35377, N35376, N35375, N35374, N35373, N35372, N35371, N35370, N35369, N35368, N35367, N35366, N35365, N35364, N35363, N35362, N35361, N35360, N35359, N35358, N35357, N35356, N35355, N35354, N35353, N35352, N35351, N35350, N35349, N35348, N35347, N35346, N35345, N35344, N35343, N35342, N35341, N35340, N35339, N35338, N35337, N35336, N35335, N35334, N35333, N35332, N35331, N35330, N35329, N35328, N35327, N35326, N35325, N35324, N35323 } : 1'b0;
  assign N785 = N35460;
  assign N786 = N35461;
  assign N35531 = (N785)? mem_q[2016] : 
                  (N786)? N35387 : 1'b0;
  assign { N35533, N35532 } = (N785)? { N35454, N35453 } : 
                              (N786)? { N35465, N35464 } : 1'b0;
  assign N35534 = (N785)? N35455 : 
                  (N786)? N35466 : 1'b0;
  assign { N35598, N35597, N35596, N35595, N35594, N35593, N35592, N35591, N35590, N35589, N35588, N35587, N35586, N35585, N35584, N35583, N35582, N35581, N35580, N35579, N35578, N35577, N35576, N35575, N35574, N35573, N35572, N35571, N35570, N35569, N35568, N35567, N35566, N35565, N35564, N35563, N35562, N35561, N35560, N35559, N35558, N35557, N35556, N35555, N35554, N35553, N35552, N35551, N35550, N35549, N35548, N35547, N35546, N35545, N35544, N35543, N35542, N35541, N35540, N35539, N35538, N35537, N35536, N35535 } = (N787)? mem_q[2080:2017] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N788)? { N35451, N35450, N35449, N35448, N35447, N35446, N35445, N35444, N35443, N35442, N35441, N35440, N35439, N35438, N35437, N35436, N35435, N35434, N35433, N35432, N35431, N35430, N35429, N35428, N35427, N35426, N35425, N35424, N35423, N35422, N35421, N35420, N35419, N35418, N35417, N35416, N35415, N35414, N35413, N35412, N35411, N35410, N35409, N35408, N35407, N35406, N35405, N35404, N35403, N35402, N35401, N35400, N35399, N35398, N35397, N35396, N35395, N35394, N35393, N35392, N35391, N35390, N35389, N35388 } : 1'b0;
  assign N787 = N35457;
  assign N788 = N35458;
  assign N35599 = (N787)? mem_q[2016] : 
                  (N788)? N35452 : 1'b0;
  assign { N35601, N35600 } = (N787)? { N35454, N35453 } : 
                              (N788)? { N35533, N35532 } : 1'b0;
  assign N35602 = (N787)? N35455 : 
                  (N788)? N35534 : 1'b0;
  assign { N35666, N35665, N35664, N35663, N35662, N35661, N35660, N35659, N35658, N35657, N35656, N35655, N35654, N35653, N35652, N35651, N35650, N35649, N35648, N35647, N35646, N35645, N35644, N35643, N35642, N35641, N35640, N35639, N35638, N35637, N35636, N35635, N35634, N35633, N35632, N35631, N35630, N35629, N35628, N35627, N35626, N35625, N35624, N35623, N35622, N35621, N35620, N35619, N35618, N35617, N35616, N35615, N35614, N35613, N35612, N35611, N35610, N35609, N35608, N35607, N35606, N35605, N35604, N35603 } = (N787)? { N35386, N35385, N35384, N35383, N35382, N35381, N35380, N35379, N35378, N35377, N35376, N35375, N35374, N35373, N35372, N35371, N35370, N35369, N35368, N35367, N35366, N35365, N35364, N35363, N35362, N35361, N35360, N35359, N35358, N35357, N35356, N35355, N35354, N35353, N35352, N35351, N35350, N35349, N35348, N35347, N35346, N35345, N35344, N35343, N35342, N35341, N35340, N35339, N35338, N35337, N35336, N35335, N35334, N35333, N35332, N35331, N35330, N35329, N35328, N35327, N35326, N35325, N35324, N35323 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N788)? { N35530, N35529, N35528, N35527, N35526, N35525, N35524, N35523, N35522, N35521, N35520, N35519, N35518, N35517, N35516, N35515, N35514, N35513, N35512, N35511, N35510, N35509, N35508, N35507, N35506, N35505, N35504, N35503, N35502, N35501, N35500, N35499, N35498, N35497, N35496, N35495, N35494, N35493, N35492, N35491, N35490, N35489, N35488, N35487, N35486, N35485, N35484, N35483, N35482, N35481, N35480, N35479, N35478, N35477, N35476, N35475, N35474, N35473, N35472, N35471, N35470, N35469, N35468, N35467 } : 1'b0;
  assign N35667 = (N787)? N35387 : 
                  (N788)? N35531 : 1'b0;
  assign { N35731, N35730, N35729, N35728, N35727, N35726, N35725, N35724, N35723, N35722, N35721, N35720, N35719, N35718, N35717, N35716, N35715, N35714, N35713, N35712, N35711, N35710, N35709, N35708, N35707, N35706, N35705, N35704, N35703, N35702, N35701, N35700, N35699, N35698, N35697, N35696, N35695, N35694, N35693, N35692, N35691, N35690, N35689, N35688, N35687, N35686, N35685, N35684, N35683, N35682, N35681, N35680, N35679, N35678, N35677, N35676, N35675, N35674, N35673, N35672, N35671, N35670, N35669, N35668 } = (N624)? { N35666, N35665, N35664, N35663, N35662, N35661, N35660, N35659, N35658, N35657, N35656, N35655, N35654, N35653, N35652, N35651, N35650, N35649, N35648, N35647, N35646, N35645, N35644, N35643, N35642, N35641, N35640, N35639, N35638, N35637, N35636, N35635, N35634, N35633, N35632, N35631, N35630, N35629, N35628, N35627, N35626, N35625, N35624, N35623, N35622, N35621, N35620, N35619, N35618, N35617, N35616, N35615, N35614, N35613, N35612, N35611, N35610, N35609, N35608, N35607, N35606, N35605, N35604, N35603 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N32090)? { N35386, N35385, N35384, N35383, N35382, N35381, N35380, N35379, N35378, N35377, N35376, N35375, N35374, N35373, N35372, N35371, N35370, N35369, N35368, N35367, N35366, N35365, N35364, N35363, N35362, N35361, N35360, N35359, N35358, N35357, N35356, N35355, N35354, N35353, N35352, N35351, N35350, N35349, N35348, N35347, N35346, N35345, N35344, N35343, N35342, N35341, N35340, N35339, N35338, N35337, N35336, N35335, N35334, N35333, N35332, N35331, N35330, N35329, N35328, N35327, N35326, N35325, N35324, N35323 } : 1'b0;
  assign N35732 = (N624)? N35667 : 
                  (N32090)? N35387 : 1'b0;
  assign { N35796, N35795, N35794, N35793, N35792, N35791, N35790, N35789, N35788, N35787, N35786, N35785, N35784, N35783, N35782, N35781, N35780, N35779, N35778, N35777, N35776, N35775, N35774, N35773, N35772, N35771, N35770, N35769, N35768, N35767, N35766, N35765, N35764, N35763, N35762, N35761, N35760, N35759, N35758, N35757, N35756, N35755, N35754, N35753, N35752, N35751, N35750, N35749, N35748, N35747, N35746, N35745, N35744, N35743, N35742, N35741, N35740, N35739, N35738, N35737, N35736, N35735, N35734, N35733 } = (N624)? { N35598, N35597, N35596, N35595, N35594, N35593, N35592, N35591, N35590, N35589, N35588, N35587, N35586, N35585, N35584, N35583, N35582, N35581, N35580, N35579, N35578, N35577, N35576, N35575, N35574, N35573, N35572, N35571, N35570, N35569, N35568, N35567, N35566, N35565, N35564, N35563, N35562, N35561, N35560, N35559, N35558, N35557, N35556, N35555, N35554, N35553, N35552, N35551, N35550, N35549, N35548, N35547, N35546, N35545, N35544, N35543, N35542, N35541, N35540, N35539, N35538, N35537, N35536, N35535 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N32090)? { N35451, N35450, N35449, N35448, N35447, N35446, N35445, N35444, N35443, N35442, N35441, N35440, N35439, N35438, N35437, N35436, N35435, N35434, N35433, N35432, N35431, N35430, N35429, N35428, N35427, N35426, N35425, N35424, N35423, N35422, N35421, N35420, N35419, N35418, N35417, N35416, N35415, N35414, N35413, N35412, N35411, N35410, N35409, N35408, N35407, N35406, N35405, N35404, N35403, N35402, N35401, N35400, N35399, N35398, N35397, N35396, N35395, N35394, N35393, N35392, N35391, N35390, N35389, N35388 } : 1'b0;
  assign N35797 = (N624)? N35599 : 
                  (N32090)? N35452 : 1'b0;
  assign { N35799, N35798 } = (N624)? { N35601, N35600 } : 
                              (N32090)? { N35454, N35453 } : 1'b0;
  assign N35800 = (N624)? N35602 : 
                  (N32090)? N35455 : 1'b0;
  assign { N35810, N35809 } = (N789)? mem_q[2381:2380] : 
                              (N790)? { N35799, N35798 } : 1'b0;
  assign N789 = N35807;
  assign N790 = N35808;
  assign N35811 = (N789)? mem_q[2379] : 
                  (N790)? N35800 : 1'b0;
  assign { N35875, N35874, N35873, N35872, N35871, N35870, N35869, N35868, N35867, N35866, N35865, N35864, N35863, N35862, N35861, N35860, N35859, N35858, N35857, N35856, N35855, N35854, N35853, N35852, N35851, N35850, N35849, N35848, N35847, N35846, N35845, N35844, N35843, N35842, N35841, N35840, N35839, N35838, N35837, N35836, N35835, N35834, N35833, N35832, N35831, N35830, N35829, N35828, N35827, N35826, N35825, N35824, N35823, N35822, N35821, N35820, N35819, N35818, N35817, N35816, N35815, N35814, N35813, N35812 } = (N791)? mem_q[2443:2380] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N792)? { N35731, N35730, N35729, N35728, N35727, N35726, N35725, N35724, N35723, N35722, N35721, N35720, N35719, N35718, N35717, N35716, N35715, N35714, N35713, N35712, N35711, N35710, N35709, N35708, N35707, N35706, N35705, N35704, N35703, N35702, N35701, N35700, N35699, N35698, N35697, N35696, N35695, N35694, N35693, N35692, N35691, N35690, N35689, N35688, N35687, N35686, N35685, N35684, N35683, N35682, N35681, N35680, N35679, N35678, N35677, N35676, N35675, N35674, N35673, N35672, N35671, N35670, N35669, N35668 } : 1'b0;
  assign N791 = N35805;
  assign N792 = N35806;
  assign N35876 = (N791)? mem_q[2379] : 
                  (N792)? N35732 : 1'b0;
  assign { N35878, N35877 } = (N791)? { N35799, N35798 } : 
                              (N792)? { N35810, N35809 } : 1'b0;
  assign N35879 = (N791)? N35800 : 
                  (N792)? N35811 : 1'b0;
  assign { N35943, N35942, N35941, N35940, N35939, N35938, N35937, N35936, N35935, N35934, N35933, N35932, N35931, N35930, N35929, N35928, N35927, N35926, N35925, N35924, N35923, N35922, N35921, N35920, N35919, N35918, N35917, N35916, N35915, N35914, N35913, N35912, N35911, N35910, N35909, N35908, N35907, N35906, N35905, N35904, N35903, N35902, N35901, N35900, N35899, N35898, N35897, N35896, N35895, N35894, N35893, N35892, N35891, N35890, N35889, N35888, N35887, N35886, N35885, N35884, N35883, N35882, N35881, N35880 } = (N793)? mem_q[2443:2380] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N794)? { N35796, N35795, N35794, N35793, N35792, N35791, N35790, N35789, N35788, N35787, N35786, N35785, N35784, N35783, N35782, N35781, N35780, N35779, N35778, N35777, N35776, N35775, N35774, N35773, N35772, N35771, N35770, N35769, N35768, N35767, N35766, N35765, N35764, N35763, N35762, N35761, N35760, N35759, N35758, N35757, N35756, N35755, N35754, N35753, N35752, N35751, N35750, N35749, N35748, N35747, N35746, N35745, N35744, N35743, N35742, N35741, N35740, N35739, N35738, N35737, N35736, N35735, N35734, N35733 } : 1'b0;
  assign N793 = N35802;
  assign N794 = N35803;
  assign N35944 = (N793)? mem_q[2379] : 
                  (N794)? N35797 : 1'b0;
  assign { N35946, N35945 } = (N793)? { N35799, N35798 } : 
                              (N794)? { N35878, N35877 } : 1'b0;
  assign N35947 = (N793)? N35800 : 
                  (N794)? N35879 : 1'b0;
  assign { N36011, N36010, N36009, N36008, N36007, N36006, N36005, N36004, N36003, N36002, N36001, N36000, N35999, N35998, N35997, N35996, N35995, N35994, N35993, N35992, N35991, N35990, N35989, N35988, N35987, N35986, N35985, N35984, N35983, N35982, N35981, N35980, N35979, N35978, N35977, N35976, N35975, N35974, N35973, N35972, N35971, N35970, N35969, N35968, N35967, N35966, N35965, N35964, N35963, N35962, N35961, N35960, N35959, N35958, N35957, N35956, N35955, N35954, N35953, N35952, N35951, N35950, N35949, N35948 } = (N793)? { N35731, N35730, N35729, N35728, N35727, N35726, N35725, N35724, N35723, N35722, N35721, N35720, N35719, N35718, N35717, N35716, N35715, N35714, N35713, N35712, N35711, N35710, N35709, N35708, N35707, N35706, N35705, N35704, N35703, N35702, N35701, N35700, N35699, N35698, N35697, N35696, N35695, N35694, N35693, N35692, N35691, N35690, N35689, N35688, N35687, N35686, N35685, N35684, N35683, N35682, N35681, N35680, N35679, N35678, N35677, N35676, N35675, N35674, N35673, N35672, N35671, N35670, N35669, N35668 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N794)? { N35875, N35874, N35873, N35872, N35871, N35870, N35869, N35868, N35867, N35866, N35865, N35864, N35863, N35862, N35861, N35860, N35859, N35858, N35857, N35856, N35855, N35854, N35853, N35852, N35851, N35850, N35849, N35848, N35847, N35846, N35845, N35844, N35843, N35842, N35841, N35840, N35839, N35838, N35837, N35836, N35835, N35834, N35833, N35832, N35831, N35830, N35829, N35828, N35827, N35826, N35825, N35824, N35823, N35822, N35821, N35820, N35819, N35818, N35817, N35816, N35815, N35814, N35813, N35812 } : 1'b0;
  assign N36012 = (N793)? N35732 : 
                  (N794)? N35876 : 1'b0;
  assign { N36076, N36075, N36074, N36073, N36072, N36071, N36070, N36069, N36068, N36067, N36066, N36065, N36064, N36063, N36062, N36061, N36060, N36059, N36058, N36057, N36056, N36055, N36054, N36053, N36052, N36051, N36050, N36049, N36048, N36047, N36046, N36045, N36044, N36043, N36042, N36041, N36040, N36039, N36038, N36037, N36036, N36035, N36034, N36033, N36032, N36031, N36030, N36029, N36028, N36027, N36026, N36025, N36024, N36023, N36022, N36021, N36020, N36019, N36018, N36017, N36016, N36015, N36014, N36013 } = (N688)? { N36011, N36010, N36009, N36008, N36007, N36006, N36005, N36004, N36003, N36002, N36001, N36000, N35999, N35998, N35997, N35996, N35995, N35994, N35993, N35992, N35991, N35990, N35989, N35988, N35987, N35986, N35985, N35984, N35983, N35982, N35981, N35980, N35979, N35978, N35977, N35976, N35975, N35974, N35973, N35972, N35971, N35970, N35969, N35968, N35967, N35966, N35965, N35964, N35963, N35962, N35961, N35960, N35959, N35958, N35957, N35956, N35955, N35954, N35953, N35952, N35951, N35950, N35949, N35948 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N32721)? { N35731, N35730, N35729, N35728, N35727, N35726, N35725, N35724, N35723, N35722, N35721, N35720, N35719, N35718, N35717, N35716, N35715, N35714, N35713, N35712, N35711, N35710, N35709, N35708, N35707, N35706, N35705, N35704, N35703, N35702, N35701, N35700, N35699, N35698, N35697, N35696, N35695, N35694, N35693, N35692, N35691, N35690, N35689, N35688, N35687, N35686, N35685, N35684, N35683, N35682, N35681, N35680, N35679, N35678, N35677, N35676, N35675, N35674, N35673, N35672, N35671, N35670, N35669, N35668 } : 1'b0;
  assign N36077 = (N688)? N36012 : 
                  (N32721)? N35732 : 1'b0;
  assign { N36141, N36140, N36139, N36138, N36137, N36136, N36135, N36134, N36133, N36132, N36131, N36130, N36129, N36128, N36127, N36126, N36125, N36124, N36123, N36122, N36121, N36120, N36119, N36118, N36117, N36116, N36115, N36114, N36113, N36112, N36111, N36110, N36109, N36108, N36107, N36106, N36105, N36104, N36103, N36102, N36101, N36100, N36099, N36098, N36097, N36096, N36095, N36094, N36093, N36092, N36091, N36090, N36089, N36088, N36087, N36086, N36085, N36084, N36083, N36082, N36081, N36080, N36079, N36078 } = (N688)? { N35943, N35942, N35941, N35940, N35939, N35938, N35937, N35936, N35935, N35934, N35933, N35932, N35931, N35930, N35929, N35928, N35927, N35926, N35925, N35924, N35923, N35922, N35921, N35920, N35919, N35918, N35917, N35916, N35915, N35914, N35913, N35912, N35911, N35910, N35909, N35908, N35907, N35906, N35905, N35904, N35903, N35902, N35901, N35900, N35899, N35898, N35897, N35896, N35895, N35894, N35893, N35892, N35891, N35890, N35889, N35888, N35887, N35886, N35885, N35884, N35883, N35882, N35881, N35880 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N32721)? { N35796, N35795, N35794, N35793, N35792, N35791, N35790, N35789, N35788, N35787, N35786, N35785, N35784, N35783, N35782, N35781, N35780, N35779, N35778, N35777, N35776, N35775, N35774, N35773, N35772, N35771, N35770, N35769, N35768, N35767, N35766, N35765, N35764, N35763, N35762, N35761, N35760, N35759, N35758, N35757, N35756, N35755, N35754, N35753, N35752, N35751, N35750, N35749, N35748, N35747, N35746, N35745, N35744, N35743, N35742, N35741, N35740, N35739, N35738, N35737, N35736, N35735, N35734, N35733 } : 1'b0;
  assign N36142 = (N688)? N35944 : 
                  (N32721)? N35797 : 1'b0;
  assign { N36144, N36143 } = (N688)? { N35946, N35945 } : 
                              (N32721)? { N35799, N35798 } : 1'b0;
  assign N36145 = (N688)? N35947 : 
                  (N32721)? N35800 : 1'b0;
  assign { N36155, N36154 } = (N795)? mem_q[2744:2743] : 
                              (N796)? { N36144, N36143 } : 1'b0;
  assign N795 = N36152;
  assign N796 = N36153;
  assign N36156 = (N795)? mem_q[2742] : 
                  (N796)? N36145 : 1'b0;
  assign { N36220, N36219, N36218, N36217, N36216, N36215, N36214, N36213, N36212, N36211, N36210, N36209, N36208, N36207, N36206, N36205, N36204, N36203, N36202, N36201, N36200, N36199, N36198, N36197, N36196, N36195, N36194, N36193, N36192, N36191, N36190, N36189, N36188, N36187, N36186, N36185, N36184, N36183, N36182, N36181, N36180, N36179, N36178, N36177, N36176, N36175, N36174, N36173, N36172, N36171, N36170, N36169, N36168, N36167, N36166, N36165, N36164, N36163, N36162, N36161, N36160, N36159, N36158, N36157 } = (N797)? mem_q[2806:2743] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N798)? { N36076, N36075, N36074, N36073, N36072, N36071, N36070, N36069, N36068, N36067, N36066, N36065, N36064, N36063, N36062, N36061, N36060, N36059, N36058, N36057, N36056, N36055, N36054, N36053, N36052, N36051, N36050, N36049, N36048, N36047, N36046, N36045, N36044, N36043, N36042, N36041, N36040, N36039, N36038, N36037, N36036, N36035, N36034, N36033, N36032, N36031, N36030, N36029, N36028, N36027, N36026, N36025, N36024, N36023, N36022, N36021, N36020, N36019, N36018, N36017, N36016, N36015, N36014, N36013 } : 1'b0;
  assign N797 = N36150;
  assign N798 = N36151;
  assign N36221 = (N797)? mem_q[2742] : 
                  (N798)? N36077 : 1'b0;
  assign { N36223, N36222 } = (N797)? { N36144, N36143 } : 
                              (N798)? { N36155, N36154 } : 1'b0;
  assign N36224 = (N797)? N36145 : 
                  (N798)? N36156 : 1'b0;
  assign { N36288, N36287, N36286, N36285, N36284, N36283, N36282, N36281, N36280, N36279, N36278, N36277, N36276, N36275, N36274, N36273, N36272, N36271, N36270, N36269, N36268, N36267, N36266, N36265, N36264, N36263, N36262, N36261, N36260, N36259, N36258, N36257, N36256, N36255, N36254, N36253, N36252, N36251, N36250, N36249, N36248, N36247, N36246, N36245, N36244, N36243, N36242, N36241, N36240, N36239, N36238, N36237, N36236, N36235, N36234, N36233, N36232, N36231, N36230, N36229, N36228, N36227, N36226, N36225 } = (N799)? mem_q[2806:2743] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N800)? { N36141, N36140, N36139, N36138, N36137, N36136, N36135, N36134, N36133, N36132, N36131, N36130, N36129, N36128, N36127, N36126, N36125, N36124, N36123, N36122, N36121, N36120, N36119, N36118, N36117, N36116, N36115, N36114, N36113, N36112, N36111, N36110, N36109, N36108, N36107, N36106, N36105, N36104, N36103, N36102, N36101, N36100, N36099, N36098, N36097, N36096, N36095, N36094, N36093, N36092, N36091, N36090, N36089, N36088, N36087, N36086, N36085, N36084, N36083, N36082, N36081, N36080, N36079, N36078 } : 1'b0;
  assign N799 = N36147;
  assign N800 = N36148;
  assign N36289 = (N799)? mem_q[2742] : 
                  (N800)? N36142 : 1'b0;
  assign { N36291, N36290 } = (N799)? { N36144, N36143 } : 
                              (N800)? { N36223, N36222 } : 1'b0;
  assign N36292 = (N799)? N36145 : 
                  (N800)? N36224 : 1'b0;
  assign { N36356, N36355, N36354, N36353, N36352, N36351, N36350, N36349, N36348, N36347, N36346, N36345, N36344, N36343, N36342, N36341, N36340, N36339, N36338, N36337, N36336, N36335, N36334, N36333, N36332, N36331, N36330, N36329, N36328, N36327, N36326, N36325, N36324, N36323, N36322, N36321, N36320, N36319, N36318, N36317, N36316, N36315, N36314, N36313, N36312, N36311, N36310, N36309, N36308, N36307, N36306, N36305, N36304, N36303, N36302, N36301, N36300, N36299, N36298, N36297, N36296, N36295, N36294, N36293 } = (N799)? { N36076, N36075, N36074, N36073, N36072, N36071, N36070, N36069, N36068, N36067, N36066, N36065, N36064, N36063, N36062, N36061, N36060, N36059, N36058, N36057, N36056, N36055, N36054, N36053, N36052, N36051, N36050, N36049, N36048, N36047, N36046, N36045, N36044, N36043, N36042, N36041, N36040, N36039, N36038, N36037, N36036, N36035, N36034, N36033, N36032, N36031, N36030, N36029, N36028, N36027, N36026, N36025, N36024, N36023, N36022, N36021, N36020, N36019, N36018, N36017, N36016, N36015, N36014, N36013 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N800)? { N36220, N36219, N36218, N36217, N36216, N36215, N36214, N36213, N36212, N36211, N36210, N36209, N36208, N36207, N36206, N36205, N36204, N36203, N36202, N36201, N36200, N36199, N36198, N36197, N36196, N36195, N36194, N36193, N36192, N36191, N36190, N36189, N36188, N36187, N36186, N36185, N36184, N36183, N36182, N36181, N36180, N36179, N36178, N36177, N36176, N36175, N36174, N36173, N36172, N36171, N36170, N36169, N36168, N36167, N36166, N36165, N36164, N36163, N36162, N36161, N36160, N36159, N36158, N36157 } : 1'b0;
  assign N36357 = (N799)? N36077 : 
                  (N800)? N36221 : 1'b0;
  assign { N36421, N36420, N36419, N36418, N36417, N36416, N36415, N36414, N36413, N36412, N36411, N36410, N36409, N36408, N36407, N36406, N36405, N36404, N36403, N36402, N36401, N36400, N36399, N36398, N36397, N36396, N36395, N36394, N36393, N36392, N36391, N36390, N36389, N36388, N36387, N36386, N36385, N36384, N36383, N36382, N36381, N36380, N36379, N36378, N36377, N36376, N36375, N36374, N36373, N36372, N36371, N36370, N36369, N36368, N36367, N36366, N36365, N36364, N36363, N36362, N36361, N36360, N36359, N36358 } = (N752)? { N36356, N36355, N36354, N36353, N36352, N36351, N36350, N36349, N36348, N36347, N36346, N36345, N36344, N36343, N36342, N36341, N36340, N36339, N36338, N36337, N36336, N36335, N36334, N36333, N36332, N36331, N36330, N36329, N36328, N36327, N36326, N36325, N36324, N36323, N36322, N36321, N36320, N36319, N36318, N36317, N36316, N36315, N36314, N36313, N36312, N36311, N36310, N36309, N36308, N36307, N36306, N36305, N36304, N36303, N36302, N36301, N36300, N36299, N36298, N36297, N36296, N36295, N36294, N36293 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N33352)? { N36076, N36075, N36074, N36073, N36072, N36071, N36070, N36069, N36068, N36067, N36066, N36065, N36064, N36063, N36062, N36061, N36060, N36059, N36058, N36057, N36056, N36055, N36054, N36053, N36052, N36051, N36050, N36049, N36048, N36047, N36046, N36045, N36044, N36043, N36042, N36041, N36040, N36039, N36038, N36037, N36036, N36035, N36034, N36033, N36032, N36031, N36030, N36029, N36028, N36027, N36026, N36025, N36024, N36023, N36022, N36021, N36020, N36019, N36018, N36017, N36016, N36015, N36014, N36013 } : 1'b0;
  assign N36422 = (N752)? N36357 : 
                  (N33352)? N36077 : 1'b0;
  assign { N36486, N36485, N36484, N36483, N36482, N36481, N36480, N36479, N36478, N36477, N36476, N36475, N36474, N36473, N36472, N36471, N36470, N36469, N36468, N36467, N36466, N36465, N36464, N36463, N36462, N36461, N36460, N36459, N36458, N36457, N36456, N36455, N36454, N36453, N36452, N36451, N36450, N36449, N36448, N36447, N36446, N36445, N36444, N36443, N36442, N36441, N36440, N36439, N36438, N36437, N36436, N36435, N36434, N36433, N36432, N36431, N36430, N36429, N36428, N36427, N36426, N36425, N36424, N36423 } = (N752)? { N36288, N36287, N36286, N36285, N36284, N36283, N36282, N36281, N36280, N36279, N36278, N36277, N36276, N36275, N36274, N36273, N36272, N36271, N36270, N36269, N36268, N36267, N36266, N36265, N36264, N36263, N36262, N36261, N36260, N36259, N36258, N36257, N36256, N36255, N36254, N36253, N36252, N36251, N36250, N36249, N36248, N36247, N36246, N36245, N36244, N36243, N36242, N36241, N36240, N36239, N36238, N36237, N36236, N36235, N36234, N36233, N36232, N36231, N36230, N36229, N36228, N36227, N36226, N36225 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N33352)? { N36141, N36140, N36139, N36138, N36137, N36136, N36135, N36134, N36133, N36132, N36131, N36130, N36129, N36128, N36127, N36126, N36125, N36124, N36123, N36122, N36121, N36120, N36119, N36118, N36117, N36116, N36115, N36114, N36113, N36112, N36111, N36110, N36109, N36108, N36107, N36106, N36105, N36104, N36103, N36102, N36101, N36100, N36099, N36098, N36097, N36096, N36095, N36094, N36093, N36092, N36091, N36090, N36089, N36088, N36087, N36086, N36085, N36084, N36083, N36082, N36081, N36080, N36079, N36078 } : 1'b0;
  assign N36487 = (N752)? N36289 : 
                  (N33352)? N36142 : 1'b0;
  assign { N36489, N36488 } = (N752)? { N36291, N36290 } : 
                              (N33352)? { N36144, N36143 } : 1'b0;
  assign N36490 = (N752)? N36292 : 
                  (N33352)? N36145 : 1'b0;
  assign { N36564, N36563, N36562, N36561, N36560, N36559, N36558, N36557, N36556, N36555, N36554, N36553, N36552, N36551, N36550, N36549, N36548, N36547, N36546, N36545, N36544, N36543, N36542, N36541, N36540, N36539, N36538, N36537, N36536, N36535, N36534, N36533, N36532, N36531, N36530, N36529, N36528, N36527, N36526, N36525, N36524, N36523, N36522, N36521, N36520, N36519, N36518, N36517, N36516, N36515, N36514, N36513, N36512, N36511, N36510, N36509, N36508, N36507, N36506, N36505, N36504, N36503, N36502, N36501 } = (N801)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N802)? { N36486, N36485, N36484, N36483, N36482, N36481, N36480, N36479, N36478, N36477, N36476, N36475, N36474, N36473, N36472, N36471, N36470, N36469, N36468, N36467, N36466, N36465, N36464, N36463, N36462, N36461, N36460, N36459, N36458, N36457, N36456, N36455, N36454, N36453, N36452, N36451, N36450, N36449, N36448, N36447, N36446, N36445, N36444, N36443, N36442, N36441, N36440, N36439, N36438, N36437, N36436, N36435, N36434, N36433, N36432, N36431, N36430, N36429, N36428, N36427, N36426, N36425, N36424, N36423 } : 1'b0;
  assign N801 = N36499;
  assign N802 = N36500;
  assign N36565 = (N801)? wb_valid_i[0] : 
                  (N802)? N36487 : 1'b0;
  assign { N36633, N36632, N36631, N36630, N36629, N36628, N36627, N36626, N36625, N36624, N36623, N36622, N36621, N36620, N36619, N36618, N36617, N36616, N36615, N36614, N36613, N36612, N36611, N36610, N36609, N36608, N36607, N36606, N36605, N36604, N36603, N36602, N36601, N36600, N36599, N36598, N36597, N36596, N36595, N36594, N36593, N36592, N36591, N36590, N36589, N36588, N36587, N36586, N36585, N36584, N36583, N36582, N36581, N36580, N36579, N36578, N36577, N36576, N36575, N36574, N36573, N36572, N36571, N36570 } = (N803)? wbdata_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N804)? { N36421, N36420, N36419, N36418, N36417, N36416, N36415, N36414, N36413, N36412, N36411, N36410, N36409, N36408, N36407, N36406, N36405, N36404, N36403, N36402, N36401, N36400, N36399, N36398, N36397, N36396, N36395, N36394, N36393, N36392, N36391, N36390, N36389, N36388, N36387, N36386, N36385, N36384, N36383, N36382, N36381, N36380, N36379, N36378, N36377, N36376, N36375, N36374, N36373, N36372, N36371, N36370, N36369, N36368, N36367, N36366, N36365, N36364, N36363, N36362, N36361, N36360, N36359, N36358 } : 1'b0;
  assign N803 = N36568;
  assign N804 = N36569;
  assign N36634 = (N803)? wb_valid_i[0] : 
                  (N804)? N36422 : 1'b0;
  assign N36635 = (N803)? 1'b0 : 
                  (N804)? N36500 : 1'b0;
  assign { N36642, N36641 } = (N805)? wbdata_i[1:0] : 
                              (N806)? { N36489, N36488 } : 1'b0;
  assign N805 = N36639;
  assign N806 = N36640;
  assign N36643 = (N805)? wb_valid_i[0] : 
                  (N806)? N36490 : 1'b0;
  assign N36644 = (N805)? 1'b0 : 
                  (N806)? N36635 : 1'b0;
  assign { N36721, N36720, N36719, N36718, N36717, N36716, N36715, N36714, N36713, N36712, N36711, N36710, N36709, N36708, N36707, N36706, N36705, N36704, N36703, N36702, N36701, N36700, N36699, N36698, N36697, N36696, N36695, N36694, N36693, N36692, N36691, N36690, N36689, N36688, N36687, N36686, N36685, N36684, N36683, N36682, N36681, N36680, N36679, N36678, N36677, N36676, N36675, N36674, N36673, N36672, N36671, N36670, N36669, N36668, N36667, N36666, N36665, N36664, N36663, N36662, N36661, N36660, N36659, N36658 } = (N807)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N808)? { N36564, N36563, N36562, N36561, N36560, N36559, N36558, N36557, N36556, N36555, N36554, N36553, N36552, N36551, N36550, N36549, N36548, N36547, N36546, N36545, N36544, N36543, N36542, N36541, N36540, N36539, N36538, N36537, N36536, N36535, N36534, N36533, N36532, N36531, N36530, N36529, N36528, N36527, N36526, N36525, N36524, N36523, N36522, N36521, N36520, N36519, N36518, N36517, N36516, N36515, N36514, N36513, N36512, N36511, N36510, N36509, N36508, N36507, N36506, N36505, N36504, N36503, N36502, N36501 } : 1'b0;
  assign N807 = N36656;
  assign N808 = N36657;
  assign N36722 = (N807)? wb_valid_i[1] : 
                  (N808)? N36565 : 1'b0;
  assign N36723 = (N807)? 1'b0 : 
                  (N808)? N36644 : 1'b0;
  assign { N36792, N36791, N36790, N36789, N36788, N36787, N36786, N36785, N36784, N36783, N36782, N36781, N36780, N36779, N36778, N36777, N36776, N36775, N36774, N36773, N36772, N36771, N36770, N36769, N36768, N36767, N36766, N36765, N36764, N36763, N36762, N36761, N36760, N36759, N36758, N36757, N36756, N36755, N36754, N36753, N36752, N36751, N36750, N36749, N36748, N36747, N36746, N36745, N36744, N36743, N36742, N36741, N36740, N36739, N36738, N36737, N36736, N36735, N36734, N36733, N36732, N36731, N36730, N36729 } = (N809)? wbdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N810)? { N36633, N36632, N36631, N36630, N36629, N36628, N36627, N36626, N36625, N36624, N36623, N36622, N36621, N36620, N36619, N36618, N36617, N36616, N36615, N36614, N36613, N36612, N36611, N36610, N36609, N36608, N36607, N36606, N36605, N36604, N36603, N36602, N36601, N36600, N36599, N36598, N36597, N36596, N36595, N36594, N36593, N36592, N36591, N36590, N36589, N36588, N36587, N36586, N36585, N36584, N36583, N36582, N36581, N36580, N36579, N36578, N36577, N36576, N36575, N36574, N36573, N36572, N36571, N36570 } : 1'b0;
  assign N809 = N36727;
  assign N810 = N36728;
  assign N36793 = (N809)? wb_valid_i[1] : 
                  (N810)? N36634 : 1'b0;
  assign N36794 = (N809)? 1'b0 : 
                  (N810)? N36723 : 1'b0;
  assign { N36801, N36800 } = (N811)? wbdata_i[65:64] : 
                              (N812)? { N36642, N36641 } : 1'b0;
  assign N811 = N36798;
  assign N812 = N36799;
  assign N36802 = (N811)? wb_valid_i[1] : 
                  (N812)? N36643 : 1'b0;
  assign N36803 = (N811)? 1'b0 : 
                  (N812)? N36794 : 1'b0;
  assign { N36880, N36879, N36878, N36877, N36876, N36875, N36874, N36873, N36872, N36871, N36870, N36869, N36868, N36867, N36866, N36865, N36864, N36863, N36862, N36861, N36860, N36859, N36858, N36857, N36856, N36855, N36854, N36853, N36852, N36851, N36850, N36849, N36848, N36847, N36846, N36845, N36844, N36843, N36842, N36841, N36840, N36839, N36838, N36837, N36836, N36835, N36834, N36833, N36832, N36831, N36830, N36829, N36828, N36827, N36826, N36825, N36824, N36823, N36822, N36821, N36820, N36819, N36818, N36817 } = (N813)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N814)? { N36721, N36720, N36719, N36718, N36717, N36716, N36715, N36714, N36713, N36712, N36711, N36710, N36709, N36708, N36707, N36706, N36705, N36704, N36703, N36702, N36701, N36700, N36699, N36698, N36697, N36696, N36695, N36694, N36693, N36692, N36691, N36690, N36689, N36688, N36687, N36686, N36685, N36684, N36683, N36682, N36681, N36680, N36679, N36678, N36677, N36676, N36675, N36674, N36673, N36672, N36671, N36670, N36669, N36668, N36667, N36666, N36665, N36664, N36663, N36662, N36661, N36660, N36659, N36658 } : 1'b0;
  assign N813 = N36815;
  assign N814 = N36816;
  assign N36881 = (N813)? wb_valid_i[2] : 
                  (N814)? N36722 : 1'b0;
  assign N36882 = (N813)? 1'b0 : 
                  (N814)? N36803 : 1'b0;
  assign { N36951, N36950, N36949, N36948, N36947, N36946, N36945, N36944, N36943, N36942, N36941, N36940, N36939, N36938, N36937, N36936, N36935, N36934, N36933, N36932, N36931, N36930, N36929, N36928, N36927, N36926, N36925, N36924, N36923, N36922, N36921, N36920, N36919, N36918, N36917, N36916, N36915, N36914, N36913, N36912, N36911, N36910, N36909, N36908, N36907, N36906, N36905, N36904, N36903, N36902, N36901, N36900, N36899, N36898, N36897, N36896, N36895, N36894, N36893, N36892, N36891, N36890, N36889, N36888 } = (N815)? wbdata_i[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N816)? { N36792, N36791, N36790, N36789, N36788, N36787, N36786, N36785, N36784, N36783, N36782, N36781, N36780, N36779, N36778, N36777, N36776, N36775, N36774, N36773, N36772, N36771, N36770, N36769, N36768, N36767, N36766, N36765, N36764, N36763, N36762, N36761, N36760, N36759, N36758, N36757, N36756, N36755, N36754, N36753, N36752, N36751, N36750, N36749, N36748, N36747, N36746, N36745, N36744, N36743, N36742, N36741, N36740, N36739, N36738, N36737, N36736, N36735, N36734, N36733, N36732, N36731, N36730, N36729 } : 1'b0;
  assign N815 = N36886;
  assign N816 = N36887;
  assign N36952 = (N815)? wb_valid_i[2] : 
                  (N816)? N36793 : 1'b0;
  assign N36953 = (N815)? 1'b0 : 
                  (N816)? N36882 : 1'b0;
  assign { N36960, N36959 } = (N817)? wbdata_i[129:128] : 
                              (N818)? { N36801, N36800 } : 1'b0;
  assign N817 = N36957;
  assign N818 = N36958;
  assign N36961 = (N817)? wb_valid_i[2] : 
                  (N818)? N36802 : 1'b0;
  assign N36962 = (N817)? 1'b0 : 
                  (N818)? N36953 : 1'b0;
  assign { N37039, N37038, N37037, N37036, N37035, N37034, N37033, N37032, N37031, N37030, N37029, N37028, N37027, N37026, N37025, N37024, N37023, N37022, N37021, N37020, N37019, N37018, N37017, N37016, N37015, N37014, N37013, N37012, N37011, N37010, N37009, N37008, N37007, N37006, N37005, N37004, N37003, N37002, N37001, N37000, N36999, N36998, N36997, N36996, N36995, N36994, N36993, N36992, N36991, N36990, N36989, N36988, N36987, N36986, N36985, N36984, N36983, N36982, N36981, N36980, N36979, N36978, N36977, N36976 } = (N819)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N820)? { N36880, N36879, N36878, N36877, N36876, N36875, N36874, N36873, N36872, N36871, N36870, N36869, N36868, N36867, N36866, N36865, N36864, N36863, N36862, N36861, N36860, N36859, N36858, N36857, N36856, N36855, N36854, N36853, N36852, N36851, N36850, N36849, N36848, N36847, N36846, N36845, N36844, N36843, N36842, N36841, N36840, N36839, N36838, N36837, N36836, N36835, N36834, N36833, N36832, N36831, N36830, N36829, N36828, N36827, N36826, N36825, N36824, N36823, N36822, N36821, N36820, N36819, N36818, N36817 } : 1'b0;
  assign N819 = N36974;
  assign N820 = N36975;
  assign N37040 = (N819)? wb_valid_i[3] : 
                  (N820)? N36881 : 1'b0;
  assign N37041 = (N819)? 1'b0 : 
                  (N820)? N36962 : 1'b0;
  assign { N37110, N37109, N37108, N37107, N37106, N37105, N37104, N37103, N37102, N37101, N37100, N37099, N37098, N37097, N37096, N37095, N37094, N37093, N37092, N37091, N37090, N37089, N37088, N37087, N37086, N37085, N37084, N37083, N37082, N37081, N37080, N37079, N37078, N37077, N37076, N37075, N37074, N37073, N37072, N37071, N37070, N37069, N37068, N37067, N37066, N37065, N37064, N37063, N37062, N37061, N37060, N37059, N37058, N37057, N37056, N37055, N37054, N37053, N37052, N37051, N37050, N37049, N37048, N37047 } = (N821)? wbdata_i[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N822)? { N36951, N36950, N36949, N36948, N36947, N36946, N36945, N36944, N36943, N36942, N36941, N36940, N36939, N36938, N36937, N36936, N36935, N36934, N36933, N36932, N36931, N36930, N36929, N36928, N36927, N36926, N36925, N36924, N36923, N36922, N36921, N36920, N36919, N36918, N36917, N36916, N36915, N36914, N36913, N36912, N36911, N36910, N36909, N36908, N36907, N36906, N36905, N36904, N36903, N36902, N36901, N36900, N36899, N36898, N36897, N36896, N36895, N36894, N36893, N36892, N36891, N36890, N36889, N36888 } : 1'b0;
  assign N821 = N37045;
  assign N822 = N37046;
  assign N37111 = (N821)? wb_valid_i[3] : 
                  (N822)? N36952 : 1'b0;
  assign N37112 = (N821)? 1'b0 : 
                  (N822)? N37041 : 1'b0;
  assign { N37118, N37117 } = (N823)? wbdata_i[193:192] : 
                              (N824)? { N36960, N36959 } : 1'b0;
  assign N823 = N37115;
  assign N824 = N37116;
  assign N37119 = (N823)? wb_valid_i[3] : 
                  (N824)? N36961 : 1'b0;
  assign { N37121, N37120 } = (N825)? { N37118, N37117 } : 
                              (N826)? { N36960, N36959 } : 1'b0;
  assign N825 = N37112;
  assign N826 = N37113;
  assign N37122 = (N825)? N37119 : 
                  (N826)? N36961 : 1'b0;
  assign { N37186, N37185, N37184, N37183, N37182, N37181, N37180, N37179, N37178, N37177, N37176, N37175, N37174, N37173, N37172, N37171, N37170, N37169, N37168, N37167, N37166, N37165, N37164, N37163, N37162, N37161, N37160, N37159, N37158, N37157, N37156, N37155, N37154, N37153, N37152, N37151, N37150, N37149, N37148, N37147, N37146, N37145, N37144, N37143, N37142, N37141, N37140, N37139, N37138, N37137, N37136, N37135, N37134, N37133, N37132, N37131, N37130, N37129, N37128, N37127, N37126, N37125, N37124, N37123 } = (N827)? { N37110, N37109, N37108, N37107, N37106, N37105, N37104, N37103, N37102, N37101, N37100, N37099, N37098, N37097, N37096, N37095, N37094, N37093, N37092, N37091, N37090, N37089, N37088, N37087, N37086, N37085, N37084, N37083, N37082, N37081, N37080, N37079, N37078, N37077, N37076, N37075, N37074, N37073, N37072, N37071, N37070, N37069, N37068, N37067, N37066, N37065, N37064, N37063, N37062, N37061, N37060, N37059, N37058, N37057, N37056, N37055, N37054, N37053, N37052, N37051, N37050, N37049, N37048, N37047 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N828)? { N36951, N36950, N36949, N36948, N36947, N36946, N36945, N36944, N36943, N36942, N36941, N36940, N36939, N36938, N36937, N36936, N36935, N36934, N36933, N36932, N36931, N36930, N36929, N36928, N36927, N36926, N36925, N36924, N36923, N36922, N36921, N36920, N36919, N36918, N36917, N36916, N36915, N36914, N36913, N36912, N36911, N36910, N36909, N36908, N36907, N36906, N36905, N36904, N36903, N36902, N36901, N36900, N36899, N36898, N36897, N36896, N36895, N36894, N36893, N36892, N36891, N36890, N36889, N36888 } : 1'b0;
  assign N827 = N37041;
  assign N828 = N37042;
  assign N37187 = (N827)? N37111 : 
                  (N828)? N36952 : 1'b0;
  assign { N37189, N37188 } = (N827)? { N37121, N37120 } : 
                              (N828)? { N36960, N36959 } : 1'b0;
  assign N37190 = (N827)? N37122 : 
                  (N828)? N36961 : 1'b0;
  assign { N37193, N37192 } = (N829)? { N37189, N37188 } : 
                              (N37191)? { N36960, N36959 } : 1'b0;
  assign N829 = N36962;
  assign N37194 = (N829)? N37190 : 
                  (N37191)? N36961 : 1'b0;
  assign N37195 = (N829)? N37187 : 
                  (N37191)? N36952 : 1'b0;
  assign { N37259, N37258, N37257, N37256, N37255, N37254, N37253, N37252, N37251, N37250, N37249, N37248, N37247, N37246, N37245, N37244, N37243, N37242, N37241, N37240, N37239, N37238, N37237, N37236, N37235, N37234, N37233, N37232, N37231, N37230, N37229, N37228, N37227, N37226, N37225, N37224, N37223, N37222, N37221, N37220, N37219, N37218, N37217, N37216, N37215, N37214, N37213, N37212, N37211, N37210, N37209, N37208, N37207, N37206, N37205, N37204, N37203, N37202, N37201, N37200, N37199, N37198, N37197, N37196 } = (N829)? { N37039, N37038, N37037, N37036, N37035, N37034, N37033, N37032, N37031, N37030, N37029, N37028, N37027, N37026, N37025, N37024, N37023, N37022, N37021, N37020, N37019, N37018, N37017, N37016, N37015, N37014, N37013, N37012, N37011, N37010, N37009, N37008, N37007, N37006, N37005, N37004, N37003, N37002, N37001, N37000, N36999, N36998, N36997, N36996, N36995, N36994, N36993, N36992, N36991, N36990, N36989, N36988, N36987, N36986, N36985, N36984, N36983, N36982, N36981, N36980, N36979, N36978, N36977, N36976 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N37191)? { N36880, N36879, N36878, N36877, N36876, N36875, N36874, N36873, N36872, N36871, N36870, N36869, N36868, N36867, N36866, N36865, N36864, N36863, N36862, N36861, N36860, N36859, N36858, N36857, N36856, N36855, N36854, N36853, N36852, N36851, N36850, N36849, N36848, N36847, N36846, N36845, N36844, N36843, N36842, N36841, N36840, N36839, N36838, N36837, N36836, N36835, N36834, N36833, N36832, N36831, N36830, N36829, N36828, N36827, N36826, N36825, N36824, N36823, N36822, N36821, N36820, N36819, N36818, N36817 } : 1'b0;
  assign N37260 = (N829)? N37040 : 
                  (N37191)? N36881 : 1'b0;
  assign { N37324, N37323, N37322, N37321, N37320, N37319, N37318, N37317, N37316, N37315, N37314, N37313, N37312, N37311, N37310, N37309, N37308, N37307, N37306, N37305, N37304, N37303, N37302, N37301, N37300, N37299, N37298, N37297, N37296, N37295, N37294, N37293, N37292, N37291, N37290, N37289, N37288, N37287, N37286, N37285, N37284, N37283, N37282, N37281, N37280, N37279, N37278, N37277, N37276, N37275, N37274, N37273, N37272, N37271, N37270, N37269, N37268, N37267, N37266, N37265, N37264, N37263, N37262, N37261 } = (N829)? { N37186, N37185, N37184, N37183, N37182, N37181, N37180, N37179, N37178, N37177, N37176, N37175, N37174, N37173, N37172, N37171, N37170, N37169, N37168, N37167, N37166, N37165, N37164, N37163, N37162, N37161, N37160, N37159, N37158, N37157, N37156, N37155, N37154, N37153, N37152, N37151, N37150, N37149, N37148, N37147, N37146, N37145, N37144, N37143, N37142, N37141, N37140, N37139, N37138, N37137, N37136, N37135, N37134, N37133, N37132, N37131, N37130, N37129, N37128, N37127, N37126, N37125, N37124, N37123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N37191)? { N36951, N36950, N36949, N36948, N36947, N36946, N36945, N36944, N36943, N36942, N36941, N36940, N36939, N36938, N36937, N36936, N36935, N36934, N36933, N36932, N36931, N36930, N36929, N36928, N36927, N36926, N36925, N36924, N36923, N36922, N36921, N36920, N36919, N36918, N36917, N36916, N36915, N36914, N36913, N36912, N36911, N36910, N36909, N36908, N36907, N36906, N36905, N36904, N36903, N36902, N36901, N36900, N36899, N36898, N36897, N36896, N36895, N36894, N36893, N36892, N36891, N36890, N36889, N36888 } : 1'b0;
  assign { N37326, N37325 } = (N829)? { N37193, N37192 } : 
                              (N830)? { N36960, N36959 } : 1'b0;
  assign N830 = N36963;
  assign N37327 = (N829)? N37194 : 
                  (N830)? N36961 : 1'b0;
  assign N37328 = (N829)? N37195 : 
                  (N830)? N36952 : 1'b0;
  assign { N37392, N37391, N37390, N37389, N37388, N37387, N37386, N37385, N37384, N37383, N37382, N37381, N37380, N37379, N37378, N37377, N37376, N37375, N37374, N37373, N37372, N37371, N37370, N37369, N37368, N37367, N37366, N37365, N37364, N37363, N37362, N37361, N37360, N37359, N37358, N37357, N37356, N37355, N37354, N37353, N37352, N37351, N37350, N37349, N37348, N37347, N37346, N37345, N37344, N37343, N37342, N37341, N37340, N37339, N37338, N37337, N37336, N37335, N37334, N37333, N37332, N37331, N37330, N37329 } = (N829)? { N37259, N37258, N37257, N37256, N37255, N37254, N37253, N37252, N37251, N37250, N37249, N37248, N37247, N37246, N37245, N37244, N37243, N37242, N37241, N37240, N37239, N37238, N37237, N37236, N37235, N37234, N37233, N37232, N37231, N37230, N37229, N37228, N37227, N37226, N37225, N37224, N37223, N37222, N37221, N37220, N37219, N37218, N37217, N37216, N37215, N37214, N37213, N37212, N37211, N37210, N37209, N37208, N37207, N37206, N37205, N37204, N37203, N37202, N37201, N37200, N37199, N37198, N37197, N37196 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N830)? { N36880, N36879, N36878, N36877, N36876, N36875, N36874, N36873, N36872, N36871, N36870, N36869, N36868, N36867, N36866, N36865, N36864, N36863, N36862, N36861, N36860, N36859, N36858, N36857, N36856, N36855, N36854, N36853, N36852, N36851, N36850, N36849, N36848, N36847, N36846, N36845, N36844, N36843, N36842, N36841, N36840, N36839, N36838, N36837, N36836, N36835, N36834, N36833, N36832, N36831, N36830, N36829, N36828, N36827, N36826, N36825, N36824, N36823, N36822, N36821, N36820, N36819, N36818, N36817 } : 1'b0;
  assign N37393 = (N829)? N37260 : 
                  (N830)? N36881 : 1'b0;
  assign { N37457, N37456, N37455, N37454, N37453, N37452, N37451, N37450, N37449, N37448, N37447, N37446, N37445, N37444, N37443, N37442, N37441, N37440, N37439, N37438, N37437, N37436, N37435, N37434, N37433, N37432, N37431, N37430, N37429, N37428, N37427, N37426, N37425, N37424, N37423, N37422, N37421, N37420, N37419, N37418, N37417, N37416, N37415, N37414, N37413, N37412, N37411, N37410, N37409, N37408, N37407, N37406, N37405, N37404, N37403, N37402, N37401, N37400, N37399, N37398, N37397, N37396, N37395, N37394 } = (N829)? { N37324, N37323, N37322, N37321, N37320, N37319, N37318, N37317, N37316, N37315, N37314, N37313, N37312, N37311, N37310, N37309, N37308, N37307, N37306, N37305, N37304, N37303, N37302, N37301, N37300, N37299, N37298, N37297, N37296, N37295, N37294, N37293, N37292, N37291, N37290, N37289, N37288, N37287, N37286, N37285, N37284, N37283, N37282, N37281, N37280, N37279, N37278, N37277, N37276, N37275, N37274, N37273, N37272, N37271, N37270, N37269, N37268, N37267, N37266, N37265, N37264, N37263, N37262, N37261 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N830)? { N36951, N36950, N36949, N36948, N36947, N36946, N36945, N36944, N36943, N36942, N36941, N36940, N36939, N36938, N36937, N36936, N36935, N36934, N36933, N36932, N36931, N36930, N36929, N36928, N36927, N36926, N36925, N36924, N36923, N36922, N36921, N36920, N36919, N36918, N36917, N36916, N36915, N36914, N36913, N36912, N36911, N36910, N36909, N36908, N36907, N36906, N36905, N36904, N36903, N36902, N36901, N36900, N36899, N36898, N36897, N36896, N36895, N36894, N36893, N36892, N36891, N36890, N36889, N36888 } : 1'b0;
  assign N37458 = (N831)? N37393 : 
                  (N832)? N36881 : 1'b0;
  assign N831 = N36953;
  assign N832 = N36954;
  assign { N37460, N37459 } = (N831)? { N37326, N37325 } : 
                              (N832)? { N36801, N36800 } : 1'b0;
  assign N37461 = (N831)? N37327 : 
                  (N832)? N36802 : 1'b0;
  assign { N37525, N37524, N37523, N37522, N37521, N37520, N37519, N37518, N37517, N37516, N37515, N37514, N37513, N37512, N37511, N37510, N37509, N37508, N37507, N37506, N37505, N37504, N37503, N37502, N37501, N37500, N37499, N37498, N37497, N37496, N37495, N37494, N37493, N37492, N37491, N37490, N37489, N37488, N37487, N37486, N37485, N37484, N37483, N37482, N37481, N37480, N37479, N37478, N37477, N37476, N37475, N37474, N37473, N37472, N37471, N37470, N37469, N37468, N37467, N37466, N37465, N37464, N37463, N37462 } = (N831)? { N37457, N37456, N37455, N37454, N37453, N37452, N37451, N37450, N37449, N37448, N37447, N37446, N37445, N37444, N37443, N37442, N37441, N37440, N37439, N37438, N37437, N37436, N37435, N37434, N37433, N37432, N37431, N37430, N37429, N37428, N37427, N37426, N37425, N37424, N37423, N37422, N37421, N37420, N37419, N37418, N37417, N37416, N37415, N37414, N37413, N37412, N37411, N37410, N37409, N37408, N37407, N37406, N37405, N37404, N37403, N37402, N37401, N37400, N37399, N37398, N37397, N37396, N37395, N37394 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N832)? { N36951, N36950, N36949, N36948, N36947, N36946, N36945, N36944, N36943, N36942, N36941, N36940, N36939, N36938, N36937, N36936, N36935, N36934, N36933, N36932, N36931, N36930, N36929, N36928, N36927, N36926, N36925, N36924, N36923, N36922, N36921, N36920, N36919, N36918, N36917, N36916, N36915, N36914, N36913, N36912, N36911, N36910, N36909, N36908, N36907, N36906, N36905, N36904, N36903, N36902, N36901, N36900, N36899, N36898, N36897, N36896, N36895, N36894, N36893, N36892, N36891, N36890, N36889, N36888 } : 1'b0;
  assign N37526 = (N831)? N37328 : 
                  (N832)? N36952 : 1'b0;
  assign { N37590, N37589, N37588, N37587, N37586, N37585, N37584, N37583, N37582, N37581, N37580, N37579, N37578, N37577, N37576, N37575, N37574, N37573, N37572, N37571, N37570, N37569, N37568, N37567, N37566, N37565, N37564, N37563, N37562, N37561, N37560, N37559, N37558, N37557, N37556, N37555, N37554, N37553, N37552, N37551, N37550, N37549, N37548, N37547, N37546, N37545, N37544, N37543, N37542, N37541, N37540, N37539, N37538, N37537, N37536, N37535, N37534, N37533, N37532, N37531, N37530, N37529, N37528, N37527 } = (N831)? { N37392, N37391, N37390, N37389, N37388, N37387, N37386, N37385, N37384, N37383, N37382, N37381, N37380, N37379, N37378, N37377, N37376, N37375, N37374, N37373, N37372, N37371, N37370, N37369, N37368, N37367, N37366, N37365, N37364, N37363, N37362, N37361, N37360, N37359, N37358, N37357, N37356, N37355, N37354, N37353, N37352, N37351, N37350, N37349, N37348, N37347, N37346, N37345, N37344, N37343, N37342, N37341, N37340, N37339, N37338, N37337, N37336, N37335, N37334, N37333, N37332, N37331, N37330, N37329 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N832)? { N36880, N36879, N36878, N36877, N36876, N36875, N36874, N36873, N36872, N36871, N36870, N36869, N36868, N36867, N36866, N36865, N36864, N36863, N36862, N36861, N36860, N36859, N36858, N36857, N36856, N36855, N36854, N36853, N36852, N36851, N36850, N36849, N36848, N36847, N36846, N36845, N36844, N36843, N36842, N36841, N36840, N36839, N36838, N36837, N36836, N36835, N36834, N36833, N36832, N36831, N36830, N36829, N36828, N36827, N36826, N36825, N36824, N36823, N36822, N36821, N36820, N36819, N36818, N36817 } : 1'b0;
  assign { N37654, N37653, N37652, N37651, N37650, N37649, N37648, N37647, N37646, N37645, N37644, N37643, N37642, N37641, N37640, N37639, N37638, N37637, N37636, N37635, N37634, N37633, N37632, N37631, N37630, N37629, N37628, N37627, N37626, N37625, N37624, N37623, N37622, N37621, N37620, N37619, N37618, N37617, N37616, N37615, N37614, N37613, N37612, N37611, N37610, N37609, N37608, N37607, N37606, N37605, N37604, N37603, N37602, N37601, N37600, N37599, N37598, N37597, N37596, N37595, N37594, N37593, N37592, N37591 } = (N833)? { N37525, N37524, N37523, N37522, N37521, N37520, N37519, N37518, N37517, N37516, N37515, N37514, N37513, N37512, N37511, N37510, N37509, N37508, N37507, N37506, N37505, N37504, N37503, N37502, N37501, N37500, N37499, N37498, N37497, N37496, N37495, N37494, N37493, N37492, N37491, N37490, N37489, N37488, N37487, N37486, N37485, N37484, N37483, N37482, N37481, N37480, N37479, N37478, N37477, N37476, N37475, N37474, N37473, N37472, N37471, N37470, N37469, N37468, N37467, N37466, N37465, N37464, N37463, N37462 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N834)? { N36792, N36791, N36790, N36789, N36788, N36787, N36786, N36785, N36784, N36783, N36782, N36781, N36780, N36779, N36778, N36777, N36776, N36775, N36774, N36773, N36772, N36771, N36770, N36769, N36768, N36767, N36766, N36765, N36764, N36763, N36762, N36761, N36760, N36759, N36758, N36757, N36756, N36755, N36754, N36753, N36752, N36751, N36750, N36749, N36748, N36747, N36746, N36745, N36744, N36743, N36742, N36741, N36740, N36739, N36738, N36737, N36736, N36735, N36734, N36733, N36732, N36731, N36730, N36729 } : 1'b0;
  assign N833 = N36882;
  assign N834 = N36883;
  assign N37655 = (N833)? N37526 : 
                  (N834)? N36793 : 1'b0;
  assign { N37719, N37718, N37717, N37716, N37715, N37714, N37713, N37712, N37711, N37710, N37709, N37708, N37707, N37706, N37705, N37704, N37703, N37702, N37701, N37700, N37699, N37698, N37697, N37696, N37695, N37694, N37693, N37692, N37691, N37690, N37689, N37688, N37687, N37686, N37685, N37684, N37683, N37682, N37681, N37680, N37679, N37678, N37677, N37676, N37675, N37674, N37673, N37672, N37671, N37670, N37669, N37668, N37667, N37666, N37665, N37664, N37663, N37662, N37661, N37660, N37659, N37658, N37657, N37656 } = (N833)? { N37590, N37589, N37588, N37587, N37586, N37585, N37584, N37583, N37582, N37581, N37580, N37579, N37578, N37577, N37576, N37575, N37574, N37573, N37572, N37571, N37570, N37569, N37568, N37567, N37566, N37565, N37564, N37563, N37562, N37561, N37560, N37559, N37558, N37557, N37556, N37555, N37554, N37553, N37552, N37551, N37550, N37549, N37548, N37547, N37546, N37545, N37544, N37543, N37542, N37541, N37540, N37539, N37538, N37537, N37536, N37535, N37534, N37533, N37532, N37531, N37530, N37529, N37528, N37527 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N834)? { N36880, N36879, N36878, N36877, N36876, N36875, N36874, N36873, N36872, N36871, N36870, N36869, N36868, N36867, N36866, N36865, N36864, N36863, N36862, N36861, N36860, N36859, N36858, N36857, N36856, N36855, N36854, N36853, N36852, N36851, N36850, N36849, N36848, N36847, N36846, N36845, N36844, N36843, N36842, N36841, N36840, N36839, N36838, N36837, N36836, N36835, N36834, N36833, N36832, N36831, N36830, N36829, N36828, N36827, N36826, N36825, N36824, N36823, N36822, N36821, N36820, N36819, N36818, N36817 } : 1'b0;
  assign N37720 = (N833)? N37458 : 
                  (N834)? N36881 : 1'b0;
  assign { N37722, N37721 } = (N833)? { N37460, N37459 } : 
                              (N834)? { N36801, N36800 } : 1'b0;
  assign N37723 = (N833)? N37461 : 
                  (N834)? N36802 : 1'b0;
  assign { N37726, N37725 } = (N835)? { N37722, N37721 } : 
                              (N37724)? { N36801, N36800 } : 1'b0;
  assign N835 = N36803;
  assign N37727 = (N835)? N37723 : 
                  (N37724)? N36802 : 1'b0;
  assign N37728 = (N835)? N37655 : 
                  (N37724)? N36793 : 1'b0;
  assign { N37792, N37791, N37790, N37789, N37788, N37787, N37786, N37785, N37784, N37783, N37782, N37781, N37780, N37779, N37778, N37777, N37776, N37775, N37774, N37773, N37772, N37771, N37770, N37769, N37768, N37767, N37766, N37765, N37764, N37763, N37762, N37761, N37760, N37759, N37758, N37757, N37756, N37755, N37754, N37753, N37752, N37751, N37750, N37749, N37748, N37747, N37746, N37745, N37744, N37743, N37742, N37741, N37740, N37739, N37738, N37737, N37736, N37735, N37734, N37733, N37732, N37731, N37730, N37729 } = (N835)? { N37719, N37718, N37717, N37716, N37715, N37714, N37713, N37712, N37711, N37710, N37709, N37708, N37707, N37706, N37705, N37704, N37703, N37702, N37701, N37700, N37699, N37698, N37697, N37696, N37695, N37694, N37693, N37692, N37691, N37690, N37689, N37688, N37687, N37686, N37685, N37684, N37683, N37682, N37681, N37680, N37679, N37678, N37677, N37676, N37675, N37674, N37673, N37672, N37671, N37670, N37669, N37668, N37667, N37666, N37665, N37664, N37663, N37662, N37661, N37660, N37659, N37658, N37657, N37656 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N37724)? { N36721, N36720, N36719, N36718, N36717, N36716, N36715, N36714, N36713, N36712, N36711, N36710, N36709, N36708, N36707, N36706, N36705, N36704, N36703, N36702, N36701, N36700, N36699, N36698, N36697, N36696, N36695, N36694, N36693, N36692, N36691, N36690, N36689, N36688, N36687, N36686, N36685, N36684, N36683, N36682, N36681, N36680, N36679, N36678, N36677, N36676, N36675, N36674, N36673, N36672, N36671, N36670, N36669, N36668, N36667, N36666, N36665, N36664, N36663, N36662, N36661, N36660, N36659, N36658 } : 1'b0;
  assign N37793 = (N835)? N37720 : 
                  (N37724)? N36722 : 1'b0;
  assign { N37857, N37856, N37855, N37854, N37853, N37852, N37851, N37850, N37849, N37848, N37847, N37846, N37845, N37844, N37843, N37842, N37841, N37840, N37839, N37838, N37837, N37836, N37835, N37834, N37833, N37832, N37831, N37830, N37829, N37828, N37827, N37826, N37825, N37824, N37823, N37822, N37821, N37820, N37819, N37818, N37817, N37816, N37815, N37814, N37813, N37812, N37811, N37810, N37809, N37808, N37807, N37806, N37805, N37804, N37803, N37802, N37801, N37800, N37799, N37798, N37797, N37796, N37795, N37794 } = (N835)? { N37654, N37653, N37652, N37651, N37650, N37649, N37648, N37647, N37646, N37645, N37644, N37643, N37642, N37641, N37640, N37639, N37638, N37637, N37636, N37635, N37634, N37633, N37632, N37631, N37630, N37629, N37628, N37627, N37626, N37625, N37624, N37623, N37622, N37621, N37620, N37619, N37618, N37617, N37616, N37615, N37614, N37613, N37612, N37611, N37610, N37609, N37608, N37607, N37606, N37605, N37604, N37603, N37602, N37601, N37600, N37599, N37598, N37597, N37596, N37595, N37594, N37593, N37592, N37591 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N37724)? { N36792, N36791, N36790, N36789, N36788, N36787, N36786, N36785, N36784, N36783, N36782, N36781, N36780, N36779, N36778, N36777, N36776, N36775, N36774, N36773, N36772, N36771, N36770, N36769, N36768, N36767, N36766, N36765, N36764, N36763, N36762, N36761, N36760, N36759, N36758, N36757, N36756, N36755, N36754, N36753, N36752, N36751, N36750, N36749, N36748, N36747, N36746, N36745, N36744, N36743, N36742, N36741, N36740, N36739, N36738, N36737, N36736, N36735, N36734, N36733, N36732, N36731, N36730, N36729 } : 1'b0;
  assign { N37859, N37858 } = (N835)? { N37726, N37725 } : 
                              (N836)? { N36801, N36800 } : 1'b0;
  assign N836 = N36804;
  assign N37860 = (N835)? N37727 : 
                  (N836)? N36802 : 1'b0;
  assign N37861 = (N835)? N37728 : 
                  (N836)? N36793 : 1'b0;
  assign { N37925, N37924, N37923, N37922, N37921, N37920, N37919, N37918, N37917, N37916, N37915, N37914, N37913, N37912, N37911, N37910, N37909, N37908, N37907, N37906, N37905, N37904, N37903, N37902, N37901, N37900, N37899, N37898, N37897, N37896, N37895, N37894, N37893, N37892, N37891, N37890, N37889, N37888, N37887, N37886, N37885, N37884, N37883, N37882, N37881, N37880, N37879, N37878, N37877, N37876, N37875, N37874, N37873, N37872, N37871, N37870, N37869, N37868, N37867, N37866, N37865, N37864, N37863, N37862 } = (N835)? { N37792, N37791, N37790, N37789, N37788, N37787, N37786, N37785, N37784, N37783, N37782, N37781, N37780, N37779, N37778, N37777, N37776, N37775, N37774, N37773, N37772, N37771, N37770, N37769, N37768, N37767, N37766, N37765, N37764, N37763, N37762, N37761, N37760, N37759, N37758, N37757, N37756, N37755, N37754, N37753, N37752, N37751, N37750, N37749, N37748, N37747, N37746, N37745, N37744, N37743, N37742, N37741, N37740, N37739, N37738, N37737, N37736, N37735, N37734, N37733, N37732, N37731, N37730, N37729 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N836)? { N36721, N36720, N36719, N36718, N36717, N36716, N36715, N36714, N36713, N36712, N36711, N36710, N36709, N36708, N36707, N36706, N36705, N36704, N36703, N36702, N36701, N36700, N36699, N36698, N36697, N36696, N36695, N36694, N36693, N36692, N36691, N36690, N36689, N36688, N36687, N36686, N36685, N36684, N36683, N36682, N36681, N36680, N36679, N36678, N36677, N36676, N36675, N36674, N36673, N36672, N36671, N36670, N36669, N36668, N36667, N36666, N36665, N36664, N36663, N36662, N36661, N36660, N36659, N36658 } : 1'b0;
  assign N37926 = (N835)? N37793 : 
                  (N836)? N36722 : 1'b0;
  assign { N37990, N37989, N37988, N37987, N37986, N37985, N37984, N37983, N37982, N37981, N37980, N37979, N37978, N37977, N37976, N37975, N37974, N37973, N37972, N37971, N37970, N37969, N37968, N37967, N37966, N37965, N37964, N37963, N37962, N37961, N37960, N37959, N37958, N37957, N37956, N37955, N37954, N37953, N37952, N37951, N37950, N37949, N37948, N37947, N37946, N37945, N37944, N37943, N37942, N37941, N37940, N37939, N37938, N37937, N37936, N37935, N37934, N37933, N37932, N37931, N37930, N37929, N37928, N37927 } = (N835)? { N37857, N37856, N37855, N37854, N37853, N37852, N37851, N37850, N37849, N37848, N37847, N37846, N37845, N37844, N37843, N37842, N37841, N37840, N37839, N37838, N37837, N37836, N37835, N37834, N37833, N37832, N37831, N37830, N37829, N37828, N37827, N37826, N37825, N37824, N37823, N37822, N37821, N37820, N37819, N37818, N37817, N37816, N37815, N37814, N37813, N37812, N37811, N37810, N37809, N37808, N37807, N37806, N37805, N37804, N37803, N37802, N37801, N37800, N37799, N37798, N37797, N37796, N37795, N37794 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N836)? { N36792, N36791, N36790, N36789, N36788, N36787, N36786, N36785, N36784, N36783, N36782, N36781, N36780, N36779, N36778, N36777, N36776, N36775, N36774, N36773, N36772, N36771, N36770, N36769, N36768, N36767, N36766, N36765, N36764, N36763, N36762, N36761, N36760, N36759, N36758, N36757, N36756, N36755, N36754, N36753, N36752, N36751, N36750, N36749, N36748, N36747, N36746, N36745, N36744, N36743, N36742, N36741, N36740, N36739, N36738, N36737, N36736, N36735, N36734, N36733, N36732, N36731, N36730, N36729 } : 1'b0;
  assign N37991 = (N837)? N37926 : 
                  (N838)? N36722 : 1'b0;
  assign N837 = N36794;
  assign N838 = N36795;
  assign { N37993, N37992 } = (N837)? { N37859, N37858 } : 
                              (N838)? { N36642, N36641 } : 1'b0;
  assign N37994 = (N837)? N37860 : 
                  (N838)? N36643 : 1'b0;
  assign { N38058, N38057, N38056, N38055, N38054, N38053, N38052, N38051, N38050, N38049, N38048, N38047, N38046, N38045, N38044, N38043, N38042, N38041, N38040, N38039, N38038, N38037, N38036, N38035, N38034, N38033, N38032, N38031, N38030, N38029, N38028, N38027, N38026, N38025, N38024, N38023, N38022, N38021, N38020, N38019, N38018, N38017, N38016, N38015, N38014, N38013, N38012, N38011, N38010, N38009, N38008, N38007, N38006, N38005, N38004, N38003, N38002, N38001, N38000, N37999, N37998, N37997, N37996, N37995 } = (N837)? { N37990, N37989, N37988, N37987, N37986, N37985, N37984, N37983, N37982, N37981, N37980, N37979, N37978, N37977, N37976, N37975, N37974, N37973, N37972, N37971, N37970, N37969, N37968, N37967, N37966, N37965, N37964, N37963, N37962, N37961, N37960, N37959, N37958, N37957, N37956, N37955, N37954, N37953, N37952, N37951, N37950, N37949, N37948, N37947, N37946, N37945, N37944, N37943, N37942, N37941, N37940, N37939, N37938, N37937, N37936, N37935, N37934, N37933, N37932, N37931, N37930, N37929, N37928, N37927 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N838)? { N36792, N36791, N36790, N36789, N36788, N36787, N36786, N36785, N36784, N36783, N36782, N36781, N36780, N36779, N36778, N36777, N36776, N36775, N36774, N36773, N36772, N36771, N36770, N36769, N36768, N36767, N36766, N36765, N36764, N36763, N36762, N36761, N36760, N36759, N36758, N36757, N36756, N36755, N36754, N36753, N36752, N36751, N36750, N36749, N36748, N36747, N36746, N36745, N36744, N36743, N36742, N36741, N36740, N36739, N36738, N36737, N36736, N36735, N36734, N36733, N36732, N36731, N36730, N36729 } : 1'b0;
  assign N38059 = (N837)? N37861 : 
                  (N838)? N36793 : 1'b0;
  assign { N38123, N38122, N38121, N38120, N38119, N38118, N38117, N38116, N38115, N38114, N38113, N38112, N38111, N38110, N38109, N38108, N38107, N38106, N38105, N38104, N38103, N38102, N38101, N38100, N38099, N38098, N38097, N38096, N38095, N38094, N38093, N38092, N38091, N38090, N38089, N38088, N38087, N38086, N38085, N38084, N38083, N38082, N38081, N38080, N38079, N38078, N38077, N38076, N38075, N38074, N38073, N38072, N38071, N38070, N38069, N38068, N38067, N38066, N38065, N38064, N38063, N38062, N38061, N38060 } = (N837)? { N37925, N37924, N37923, N37922, N37921, N37920, N37919, N37918, N37917, N37916, N37915, N37914, N37913, N37912, N37911, N37910, N37909, N37908, N37907, N37906, N37905, N37904, N37903, N37902, N37901, N37900, N37899, N37898, N37897, N37896, N37895, N37894, N37893, N37892, N37891, N37890, N37889, N37888, N37887, N37886, N37885, N37884, N37883, N37882, N37881, N37880, N37879, N37878, N37877, N37876, N37875, N37874, N37873, N37872, N37871, N37870, N37869, N37868, N37867, N37866, N37865, N37864, N37863, N37862 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N838)? { N36721, N36720, N36719, N36718, N36717, N36716, N36715, N36714, N36713, N36712, N36711, N36710, N36709, N36708, N36707, N36706, N36705, N36704, N36703, N36702, N36701, N36700, N36699, N36698, N36697, N36696, N36695, N36694, N36693, N36692, N36691, N36690, N36689, N36688, N36687, N36686, N36685, N36684, N36683, N36682, N36681, N36680, N36679, N36678, N36677, N36676, N36675, N36674, N36673, N36672, N36671, N36670, N36669, N36668, N36667, N36666, N36665, N36664, N36663, N36662, N36661, N36660, N36659, N36658 } : 1'b0;
  assign { N38187, N38186, N38185, N38184, N38183, N38182, N38181, N38180, N38179, N38178, N38177, N38176, N38175, N38174, N38173, N38172, N38171, N38170, N38169, N38168, N38167, N38166, N38165, N38164, N38163, N38162, N38161, N38160, N38159, N38158, N38157, N38156, N38155, N38154, N38153, N38152, N38151, N38150, N38149, N38148, N38147, N38146, N38145, N38144, N38143, N38142, N38141, N38140, N38139, N38138, N38137, N38136, N38135, N38134, N38133, N38132, N38131, N38130, N38129, N38128, N38127, N38126, N38125, N38124 } = (N839)? { N38058, N38057, N38056, N38055, N38054, N38053, N38052, N38051, N38050, N38049, N38048, N38047, N38046, N38045, N38044, N38043, N38042, N38041, N38040, N38039, N38038, N38037, N38036, N38035, N38034, N38033, N38032, N38031, N38030, N38029, N38028, N38027, N38026, N38025, N38024, N38023, N38022, N38021, N38020, N38019, N38018, N38017, N38016, N38015, N38014, N38013, N38012, N38011, N38010, N38009, N38008, N38007, N38006, N38005, N38004, N38003, N38002, N38001, N38000, N37999, N37998, N37997, N37996, N37995 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N840)? { N36633, N36632, N36631, N36630, N36629, N36628, N36627, N36626, N36625, N36624, N36623, N36622, N36621, N36620, N36619, N36618, N36617, N36616, N36615, N36614, N36613, N36612, N36611, N36610, N36609, N36608, N36607, N36606, N36605, N36604, N36603, N36602, N36601, N36600, N36599, N36598, N36597, N36596, N36595, N36594, N36593, N36592, N36591, N36590, N36589, N36588, N36587, N36586, N36585, N36584, N36583, N36582, N36581, N36580, N36579, N36578, N36577, N36576, N36575, N36574, N36573, N36572, N36571, N36570 } : 1'b0;
  assign N839 = N36723;
  assign N840 = N36724;
  assign N38188 = (N839)? N38059 : 
                  (N840)? N36634 : 1'b0;
  assign { N38252, N38251, N38250, N38249, N38248, N38247, N38246, N38245, N38244, N38243, N38242, N38241, N38240, N38239, N38238, N38237, N38236, N38235, N38234, N38233, N38232, N38231, N38230, N38229, N38228, N38227, N38226, N38225, N38224, N38223, N38222, N38221, N38220, N38219, N38218, N38217, N38216, N38215, N38214, N38213, N38212, N38211, N38210, N38209, N38208, N38207, N38206, N38205, N38204, N38203, N38202, N38201, N38200, N38199, N38198, N38197, N38196, N38195, N38194, N38193, N38192, N38191, N38190, N38189 } = (N839)? { N38123, N38122, N38121, N38120, N38119, N38118, N38117, N38116, N38115, N38114, N38113, N38112, N38111, N38110, N38109, N38108, N38107, N38106, N38105, N38104, N38103, N38102, N38101, N38100, N38099, N38098, N38097, N38096, N38095, N38094, N38093, N38092, N38091, N38090, N38089, N38088, N38087, N38086, N38085, N38084, N38083, N38082, N38081, N38080, N38079, N38078, N38077, N38076, N38075, N38074, N38073, N38072, N38071, N38070, N38069, N38068, N38067, N38066, N38065, N38064, N38063, N38062, N38061, N38060 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N840)? { N36721, N36720, N36719, N36718, N36717, N36716, N36715, N36714, N36713, N36712, N36711, N36710, N36709, N36708, N36707, N36706, N36705, N36704, N36703, N36702, N36701, N36700, N36699, N36698, N36697, N36696, N36695, N36694, N36693, N36692, N36691, N36690, N36689, N36688, N36687, N36686, N36685, N36684, N36683, N36682, N36681, N36680, N36679, N36678, N36677, N36676, N36675, N36674, N36673, N36672, N36671, N36670, N36669, N36668, N36667, N36666, N36665, N36664, N36663, N36662, N36661, N36660, N36659, N36658 } : 1'b0;
  assign N38253 = (N839)? N37991 : 
                  (N840)? N36722 : 1'b0;
  assign { N38255, N38254 } = (N839)? { N37993, N37992 } : 
                              (N840)? { N36642, N36641 } : 1'b0;
  assign N38256 = (N839)? N37994 : 
                  (N840)? N36643 : 1'b0;
  assign { N38259, N38258 } = (N841)? { N38255, N38254 } : 
                              (N38257)? { N36642, N36641 } : 1'b0;
  assign N841 = N36644;
  assign N38260 = (N841)? N38256 : 
                  (N38257)? N36643 : 1'b0;
  assign N38261 = (N841)? N38188 : 
                  (N38257)? N36634 : 1'b0;
  assign { N38325, N38324, N38323, N38322, N38321, N38320, N38319, N38318, N38317, N38316, N38315, N38314, N38313, N38312, N38311, N38310, N38309, N38308, N38307, N38306, N38305, N38304, N38303, N38302, N38301, N38300, N38299, N38298, N38297, N38296, N38295, N38294, N38293, N38292, N38291, N38290, N38289, N38288, N38287, N38286, N38285, N38284, N38283, N38282, N38281, N38280, N38279, N38278, N38277, N38276, N38275, N38274, N38273, N38272, N38271, N38270, N38269, N38268, N38267, N38266, N38265, N38264, N38263, N38262 } = (N841)? { N38252, N38251, N38250, N38249, N38248, N38247, N38246, N38245, N38244, N38243, N38242, N38241, N38240, N38239, N38238, N38237, N38236, N38235, N38234, N38233, N38232, N38231, N38230, N38229, N38228, N38227, N38226, N38225, N38224, N38223, N38222, N38221, N38220, N38219, N38218, N38217, N38216, N38215, N38214, N38213, N38212, N38211, N38210, N38209, N38208, N38207, N38206, N38205, N38204, N38203, N38202, N38201, N38200, N38199, N38198, N38197, N38196, N38195, N38194, N38193, N38192, N38191, N38190, N38189 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N38257)? { N36564, N36563, N36562, N36561, N36560, N36559, N36558, N36557, N36556, N36555, N36554, N36553, N36552, N36551, N36550, N36549, N36548, N36547, N36546, N36545, N36544, N36543, N36542, N36541, N36540, N36539, N36538, N36537, N36536, N36535, N36534, N36533, N36532, N36531, N36530, N36529, N36528, N36527, N36526, N36525, N36524, N36523, N36522, N36521, N36520, N36519, N36518, N36517, N36516, N36515, N36514, N36513, N36512, N36511, N36510, N36509, N36508, N36507, N36506, N36505, N36504, N36503, N36502, N36501 } : 1'b0;
  assign N38326 = (N841)? N38253 : 
                  (N38257)? N36565 : 1'b0;
  assign { N38390, N38389, N38388, N38387, N38386, N38385, N38384, N38383, N38382, N38381, N38380, N38379, N38378, N38377, N38376, N38375, N38374, N38373, N38372, N38371, N38370, N38369, N38368, N38367, N38366, N38365, N38364, N38363, N38362, N38361, N38360, N38359, N38358, N38357, N38356, N38355, N38354, N38353, N38352, N38351, N38350, N38349, N38348, N38347, N38346, N38345, N38344, N38343, N38342, N38341, N38340, N38339, N38338, N38337, N38336, N38335, N38334, N38333, N38332, N38331, N38330, N38329, N38328, N38327 } = (N841)? { N38187, N38186, N38185, N38184, N38183, N38182, N38181, N38180, N38179, N38178, N38177, N38176, N38175, N38174, N38173, N38172, N38171, N38170, N38169, N38168, N38167, N38166, N38165, N38164, N38163, N38162, N38161, N38160, N38159, N38158, N38157, N38156, N38155, N38154, N38153, N38152, N38151, N38150, N38149, N38148, N38147, N38146, N38145, N38144, N38143, N38142, N38141, N38140, N38139, N38138, N38137, N38136, N38135, N38134, N38133, N38132, N38131, N38130, N38129, N38128, N38127, N38126, N38125, N38124 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N38257)? { N36633, N36632, N36631, N36630, N36629, N36628, N36627, N36626, N36625, N36624, N36623, N36622, N36621, N36620, N36619, N36618, N36617, N36616, N36615, N36614, N36613, N36612, N36611, N36610, N36609, N36608, N36607, N36606, N36605, N36604, N36603, N36602, N36601, N36600, N36599, N36598, N36597, N36596, N36595, N36594, N36593, N36592, N36591, N36590, N36589, N36588, N36587, N36586, N36585, N36584, N36583, N36582, N36581, N36580, N36579, N36578, N36577, N36576, N36575, N36574, N36573, N36572, N36571, N36570 } : 1'b0;
  assign { N38392, N38391 } = (N841)? { N38259, N38258 } : 
                              (N842)? { N36642, N36641 } : 1'b0;
  assign N842 = N36645;
  assign N38393 = (N841)? N38260 : 
                  (N842)? N36643 : 1'b0;
  assign N38394 = (N841)? N38261 : 
                  (N842)? N36634 : 1'b0;
  assign { N38458, N38457, N38456, N38455, N38454, N38453, N38452, N38451, N38450, N38449, N38448, N38447, N38446, N38445, N38444, N38443, N38442, N38441, N38440, N38439, N38438, N38437, N38436, N38435, N38434, N38433, N38432, N38431, N38430, N38429, N38428, N38427, N38426, N38425, N38424, N38423, N38422, N38421, N38420, N38419, N38418, N38417, N38416, N38415, N38414, N38413, N38412, N38411, N38410, N38409, N38408, N38407, N38406, N38405, N38404, N38403, N38402, N38401, N38400, N38399, N38398, N38397, N38396, N38395 } = (N841)? { N38325, N38324, N38323, N38322, N38321, N38320, N38319, N38318, N38317, N38316, N38315, N38314, N38313, N38312, N38311, N38310, N38309, N38308, N38307, N38306, N38305, N38304, N38303, N38302, N38301, N38300, N38299, N38298, N38297, N38296, N38295, N38294, N38293, N38292, N38291, N38290, N38289, N38288, N38287, N38286, N38285, N38284, N38283, N38282, N38281, N38280, N38279, N38278, N38277, N38276, N38275, N38274, N38273, N38272, N38271, N38270, N38269, N38268, N38267, N38266, N38265, N38264, N38263, N38262 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N842)? { N36564, N36563, N36562, N36561, N36560, N36559, N36558, N36557, N36556, N36555, N36554, N36553, N36552, N36551, N36550, N36549, N36548, N36547, N36546, N36545, N36544, N36543, N36542, N36541, N36540, N36539, N36538, N36537, N36536, N36535, N36534, N36533, N36532, N36531, N36530, N36529, N36528, N36527, N36526, N36525, N36524, N36523, N36522, N36521, N36520, N36519, N36518, N36517, N36516, N36515, N36514, N36513, N36512, N36511, N36510, N36509, N36508, N36507, N36506, N36505, N36504, N36503, N36502, N36501 } : 1'b0;
  assign N38459 = (N841)? N38326 : 
                  (N842)? N36565 : 1'b0;
  assign { N38523, N38522, N38521, N38520, N38519, N38518, N38517, N38516, N38515, N38514, N38513, N38512, N38511, N38510, N38509, N38508, N38507, N38506, N38505, N38504, N38503, N38502, N38501, N38500, N38499, N38498, N38497, N38496, N38495, N38494, N38493, N38492, N38491, N38490, N38489, N38488, N38487, N38486, N38485, N38484, N38483, N38482, N38481, N38480, N38479, N38478, N38477, N38476, N38475, N38474, N38473, N38472, N38471, N38470, N38469, N38468, N38467, N38466, N38465, N38464, N38463, N38462, N38461, N38460 } = (N841)? { N38390, N38389, N38388, N38387, N38386, N38385, N38384, N38383, N38382, N38381, N38380, N38379, N38378, N38377, N38376, N38375, N38374, N38373, N38372, N38371, N38370, N38369, N38368, N38367, N38366, N38365, N38364, N38363, N38362, N38361, N38360, N38359, N38358, N38357, N38356, N38355, N38354, N38353, N38352, N38351, N38350, N38349, N38348, N38347, N38346, N38345, N38344, N38343, N38342, N38341, N38340, N38339, N38338, N38337, N38336, N38335, N38334, N38333, N38332, N38331, N38330, N38329, N38328, N38327 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N842)? { N36633, N36632, N36631, N36630, N36629, N36628, N36627, N36626, N36625, N36624, N36623, N36622, N36621, N36620, N36619, N36618, N36617, N36616, N36615, N36614, N36613, N36612, N36611, N36610, N36609, N36608, N36607, N36606, N36605, N36604, N36603, N36602, N36601, N36600, N36599, N36598, N36597, N36596, N36595, N36594, N36593, N36592, N36591, N36590, N36589, N36588, N36587, N36586, N36585, N36584, N36583, N36582, N36581, N36580, N36579, N36578, N36577, N36576, N36575, N36574, N36573, N36572, N36571, N36570 } : 1'b0;
  assign N38524 = (N843)? N38459 : 
                  (N844)? N36565 : 1'b0;
  assign N843 = N36635;
  assign N844 = N36636;
  assign { N38526, N38525 } = (N843)? { N38392, N38391 } : 
                              (N844)? { N36489, N36488 } : 1'b0;
  assign N38527 = (N843)? N38393 : 
                  (N844)? N36490 : 1'b0;
  assign { N38591, N38590, N38589, N38588, N38587, N38586, N38585, N38584, N38583, N38582, N38581, N38580, N38579, N38578, N38577, N38576, N38575, N38574, N38573, N38572, N38571, N38570, N38569, N38568, N38567, N38566, N38565, N38564, N38563, N38562, N38561, N38560, N38559, N38558, N38557, N38556, N38555, N38554, N38553, N38552, N38551, N38550, N38549, N38548, N38547, N38546, N38545, N38544, N38543, N38542, N38541, N38540, N38539, N38538, N38537, N38536, N38535, N38534, N38533, N38532, N38531, N38530, N38529, N38528 } = (N843)? { N38523, N38522, N38521, N38520, N38519, N38518, N38517, N38516, N38515, N38514, N38513, N38512, N38511, N38510, N38509, N38508, N38507, N38506, N38505, N38504, N38503, N38502, N38501, N38500, N38499, N38498, N38497, N38496, N38495, N38494, N38493, N38492, N38491, N38490, N38489, N38488, N38487, N38486, N38485, N38484, N38483, N38482, N38481, N38480, N38479, N38478, N38477, N38476, N38475, N38474, N38473, N38472, N38471, N38470, N38469, N38468, N38467, N38466, N38465, N38464, N38463, N38462, N38461, N38460 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N844)? { N36633, N36632, N36631, N36630, N36629, N36628, N36627, N36626, N36625, N36624, N36623, N36622, N36621, N36620, N36619, N36618, N36617, N36616, N36615, N36614, N36613, N36612, N36611, N36610, N36609, N36608, N36607, N36606, N36605, N36604, N36603, N36602, N36601, N36600, N36599, N36598, N36597, N36596, N36595, N36594, N36593, N36592, N36591, N36590, N36589, N36588, N36587, N36586, N36585, N36584, N36583, N36582, N36581, N36580, N36579, N36578, N36577, N36576, N36575, N36574, N36573, N36572, N36571, N36570 } : 1'b0;
  assign N38592 = (N843)? N38394 : 
                  (N844)? N36634 : 1'b0;
  assign { N38656, N38655, N38654, N38653, N38652, N38651, N38650, N38649, N38648, N38647, N38646, N38645, N38644, N38643, N38642, N38641, N38640, N38639, N38638, N38637, N38636, N38635, N38634, N38633, N38632, N38631, N38630, N38629, N38628, N38627, N38626, N38625, N38624, N38623, N38622, N38621, N38620, N38619, N38618, N38617, N38616, N38615, N38614, N38613, N38612, N38611, N38610, N38609, N38608, N38607, N38606, N38605, N38604, N38603, N38602, N38601, N38600, N38599, N38598, N38597, N38596, N38595, N38594, N38593 } = (N843)? { N38458, N38457, N38456, N38455, N38454, N38453, N38452, N38451, N38450, N38449, N38448, N38447, N38446, N38445, N38444, N38443, N38442, N38441, N38440, N38439, N38438, N38437, N38436, N38435, N38434, N38433, N38432, N38431, N38430, N38429, N38428, N38427, N38426, N38425, N38424, N38423, N38422, N38421, N38420, N38419, N38418, N38417, N38416, N38415, N38414, N38413, N38412, N38411, N38410, N38409, N38408, N38407, N38406, N38405, N38404, N38403, N38402, N38401, N38400, N38399, N38398, N38397, N38396, N38395 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N844)? { N36564, N36563, N36562, N36561, N36560, N36559, N36558, N36557, N36556, N36555, N36554, N36553, N36552, N36551, N36550, N36549, N36548, N36547, N36546, N36545, N36544, N36543, N36542, N36541, N36540, N36539, N36538, N36537, N36536, N36535, N36534, N36533, N36532, N36531, N36530, N36529, N36528, N36527, N36526, N36525, N36524, N36523, N36522, N36521, N36520, N36519, N36518, N36517, N36516, N36515, N36514, N36513, N36512, N36511, N36510, N36509, N36508, N36507, N36506, N36505, N36504, N36503, N36502, N36501 } : 1'b0;
  assign rs2_o = (N802)? { N38591, N38590, N38589, N38588, N38587, N38586, N38585, N38584, N38583, N38582, N38581, N38580, N38579, N38578, N38577, N38576, N38575, N38574, N38573, N38572, N38571, N38570, N38569, N38568, N38567, N38566, N38565, N38564, N38563, N38562, N38561, N38560, N38559, N38558, N38557, N38556, N38555, N38554, N38553, N38552, N38551, N38550, N38549, N38548, N38547, N38546, N38545, N38544, N38543, N38542, N38541, N38540, N38539, N38538, N38537, N38536, N38535, N38534, N38533, N38532, N38531, N38530, N38529, N38528 } : 
                 (N801)? { N36421, N36420, N36419, N36418, N36417, N36416, N36415, N36414, N36413, N36412, N36411, N36410, N36409, N36408, N36407, N36406, N36405, N36404, N36403, N36402, N36401, N36400, N36399, N36398, N36397, N36396, N36395, N36394, N36393, N36392, N36391, N36390, N36389, N36388, N36387, N36386, N36385, N36384, N36383, N36382, N36381, N36380, N36379, N36378, N36377, N36376, N36375, N36374, N36373, N36372, N36371, N36370, N36369, N36368, N36367, N36366, N36365, N36364, N36363, N36362, N36361, N36360, N36359, N36358 } : 1'b0;
  assign N38657 = (N802)? N38592 : 
                  (N801)? N36422 : 1'b0;
  assign rs1_o = (N802)? { N38656, N38655, N38654, N38653, N38652, N38651, N38650, N38649, N38648, N38647, N38646, N38645, N38644, N38643, N38642, N38641, N38640, N38639, N38638, N38637, N38636, N38635, N38634, N38633, N38632, N38631, N38630, N38629, N38628, N38627, N38626, N38625, N38624, N38623, N38622, N38621, N38620, N38619, N38618, N38617, N38616, N38615, N38614, N38613, N38612, N38611, N38610, N38609, N38608, N38607, N38606, N38605, N38604, N38603, N38602, N38601, N38600, N38599, N38598, N38597, N38596, N38595, N38594, N38593 } : 
                 (N801)? { N36564, N36563, N36562, N36561, N36560, N36559, N36558, N36557, N36556, N36555, N36554, N36553, N36552, N36551, N36550, N36549, N36548, N36547, N36546, N36545, N36544, N36543, N36542, N36541, N36540, N36539, N36538, N36537, N36536, N36535, N36534, N36533, N36532, N36531, N36530, N36529, N36528, N36527, N36526, N36525, N36524, N36523, N36522, N36521, N36520, N36519, N36518, N36517, N36516, N36515, N36514, N36513, N36512, N36511, N36510, N36509, N36508, N36507, N36506, N36505, N36504, N36503, N36502, N36501 } : 1'b0;
  assign N38658 = (N802)? N38524 : 
                  (N801)? N36565 : 1'b0;
  assign rs3_o = (N802)? { N38526, N38525 } : 
                 (N801)? { N36489, N36488 } : 1'b0;
  assign rs3_valid_o = (N802)? N38527 : 
                       (N801)? N36490 : 1'b0;
  assign rs1_valid_o = (N845)? 1'b0 : 
                       (N846)? N38658 : 1'b0;
  assign N845 = N38667;
  assign N846 = N38666;
  assign rs2_valid_o = (N847)? 1'b0 : 
                       (N848)? N38657 : 1'b0;
  assign N847 = N38673;
  assign N848 = N38672;
  assign N849 = ~commit_pointer_q[0];
  assign N850 = ~commit_pointer_q[1];
  assign N851 = N849 & N850;
  assign N852 = N849 & commit_pointer_q[1];
  assign N853 = commit_pointer_q[0] & N850;
  assign N854 = commit_pointer_q[0] & commit_pointer_q[1];
  assign N855 = ~commit_pointer_q[2];
  assign N856 = N851 & N855;
  assign N857 = N851 & commit_pointer_q[2];
  assign N858 = N853 & N855;
  assign N859 = N853 & commit_pointer_q[2];
  assign N860 = N852 & N855;
  assign N861 = N852 & commit_pointer_q[2];
  assign N862 = N854 & N855;
  assign N863 = N854 & commit_pointer_q[2];
  assign N867 = ~N864;
  assign N868 = ~N865;
  assign N869 = N867 & N868;
  assign N870 = N867 & N865;
  assign N871 = N864 & N868;
  assign N872 = N864 & N865;
  assign N873 = ~N866;
  assign N874 = N869 & N873;
  assign N875 = N869 & N866;
  assign N876 = N871 & N873;
  assign N877 = N871 & N866;
  assign N878 = N870 & N873;
  assign N879 = N870 & N866;
  assign N880 = N872 & N873;
  assign N881 = N872 & N866;
  assign N882 = ~sb_full_o;
  assign issue_instr_valid_o = N38933 & N882;
  assign N38933 = decoded_instr_valid_i & N38932;
  assign N38932 = ~unresolved_branch_i;
  assign decoded_instr_ack_o = issue_ack_i & N882;
  assign N883 = N38934 & N38935;
  assign N38934 = decoded_instr_valid_i & decoded_instr_ack_o;
  assign N38935 = ~flush_unissued_instr_i;
  assign N884 = ~N883;
  assign N896 = ~N888;
  assign N1260 = ~N889;
  assign N1624 = ~N890;
  assign N1988 = ~N891;
  assign N2352 = ~N892;
  assign N2716 = ~N893;
  assign N3080 = ~N894;
  assign N3444 = ~N895;
  assign N5886 = ~trans_id_i[0];
  assign N5887 = ~trans_id_i[1];
  assign N5888 = N5886 & N5887;
  assign N5889 = N5886 & trans_id_i[1];
  assign N5890 = trans_id_i[0] & N5887;
  assign N5891 = trans_id_i[0] & trans_id_i[1];
  assign N5892 = ~trans_id_i[2];
  assign N5893 = N5888 & N5892;
  assign N5894 = N5888 & trans_id_i[2];
  assign N5895 = N5890 & N5892;
  assign N5896 = N5890 & trans_id_i[2];
  assign N5897 = N5889 & N5892;
  assign N5898 = N5889 & trans_id_i[2];
  assign N5899 = N5891 & N5892;
  assign N5900 = N5891 & trans_id_i[2];
  assign N5902 = wb_valid_i[0] & N5901;
  assign N5903 = ~N5902;
  assign N5920 = ~N5912;
  assign N5985 = ~N5913;
  assign N6050 = ~N5914;
  assign N6115 = ~N5915;
  assign N6180 = ~N5916;
  assign N6245 = ~N5917;
  assign N6310 = ~N5918;
  assign N6375 = ~N5919;
  assign N6956 = ~ex_i[0];
  assign N7989 = ~N6953;
  assign N7990 = ~N6954;
  assign N7991 = ~N6955;
  assign N7995 = ~N6952;
  assign N7999 = N38936 | N38937;
  assign N38936 = ~N7994;
  assign N38937 = ~N7998;
  assign N8000 = ~N7999;
  assign N12121 = ~trans_id_i[3];
  assign N12122 = ~trans_id_i[4];
  assign N12123 = N12121 & N12122;
  assign N12124 = N12121 & trans_id_i[4];
  assign N12125 = trans_id_i[3] & N12122;
  assign N12126 = trans_id_i[3] & trans_id_i[4];
  assign N12127 = ~trans_id_i[5];
  assign N12128 = N12123 & N12127;
  assign N12129 = N12123 & trans_id_i[5];
  assign N12130 = N12125 & N12127;
  assign N12131 = N12125 & trans_id_i[5];
  assign N12132 = N12124 & N12127;
  assign N12133 = N12124 & trans_id_i[5];
  assign N12134 = N12126 & N12127;
  assign N12135 = N12126 & trans_id_i[5];
  assign N12137 = wb_valid_i[1] & N12136;
  assign N12138 = ~N12137;
  assign N12155 = ~N12147;
  assign N12220 = ~N12148;
  assign N12285 = ~N12149;
  assign N12350 = ~N12150;
  assign N12415 = ~N12151;
  assign N12480 = ~N12152;
  assign N12545 = ~N12153;
  assign N12610 = ~N12154;
  assign N13191 = ~ex_i[129];
  assign N14224 = ~N13188;
  assign N14225 = ~N13189;
  assign N14226 = ~N13190;
  assign N14230 = ~N13187;
  assign N14234 = N38938 | N38939;
  assign N38938 = ~N14229;
  assign N38939 = ~N14233;
  assign N14235 = ~N14234;
  assign N18356 = ~trans_id_i[6];
  assign N18357 = ~trans_id_i[7];
  assign N18358 = N18356 & N18357;
  assign N18359 = N18356 & trans_id_i[7];
  assign N18360 = trans_id_i[6] & N18357;
  assign N18361 = trans_id_i[6] & trans_id_i[7];
  assign N18362 = ~trans_id_i[8];
  assign N18363 = N18358 & N18362;
  assign N18364 = N18358 & trans_id_i[8];
  assign N18365 = N18360 & N18362;
  assign N18366 = N18360 & trans_id_i[8];
  assign N18367 = N18359 & N18362;
  assign N18368 = N18359 & trans_id_i[8];
  assign N18369 = N18361 & N18362;
  assign N18370 = N18361 & trans_id_i[8];
  assign N18372 = wb_valid_i[2] & N18371;
  assign N18373 = ~N18372;
  assign N18390 = ~N18382;
  assign N18455 = ~N18383;
  assign N18520 = ~N18384;
  assign N18585 = ~N18385;
  assign N18650 = ~N18386;
  assign N18715 = ~N18387;
  assign N18780 = ~N18388;
  assign N18845 = ~N18389;
  assign N19426 = ~ex_i[258];
  assign N20459 = ~N19423;
  assign N20460 = ~N19424;
  assign N20461 = ~N19425;
  assign N20465 = ~N19422;
  assign N20469 = N38940 | N38941;
  assign N38940 = ~N20464;
  assign N38941 = ~N20468;
  assign N20470 = ~N20469;
  assign N24591 = ~trans_id_i[9];
  assign N24592 = ~trans_id_i[10];
  assign N24593 = N24591 & N24592;
  assign N24594 = N24591 & trans_id_i[10];
  assign N24595 = trans_id_i[9] & N24592;
  assign N24596 = trans_id_i[9] & trans_id_i[10];
  assign N24597 = ~trans_id_i[11];
  assign N24598 = N24593 & N24597;
  assign N24599 = N24593 & trans_id_i[11];
  assign N24600 = N24595 & N24597;
  assign N24601 = N24595 & trans_id_i[11];
  assign N24602 = N24594 & N24597;
  assign N24603 = N24594 & trans_id_i[11];
  assign N24604 = N24596 & N24597;
  assign N24605 = N24596 & trans_id_i[11];
  assign N24607 = wb_valid_i[3] & N24606;
  assign N24608 = ~N24607;
  assign N24625 = ~N24617;
  assign N24690 = ~N24618;
  assign N24755 = ~N24619;
  assign N24820 = ~N24620;
  assign N24885 = ~N24621;
  assign N24950 = ~N24622;
  assign N25015 = ~N24623;
  assign N25080 = ~N24624;
  assign N25661 = ~ex_i[387];
  assign N26694 = ~N25658;
  assign N26695 = ~N25659;
  assign N26696 = ~N25660;
  assign N26700 = ~N25657;
  assign N26704 = N38942 | N38943;
  assign N38942 = ~N26699;
  assign N38943 = ~N26703;
  assign N26705 = ~N26704;
  assign N28778 = ~commit_ack_i[0];
  assign N28779 = commit_ack_i[0];
  assign N28788 = ~N28780;
  assign N28790 = ~N28781;
  assign N28792 = ~N28782;
  assign N28794 = ~N28783;
  assign N28796 = ~N28784;
  assign N28798 = ~N28785;
  assign N28800 = ~N28786;
  assign N28802 = ~N28787;
  assign N28812 = ~N28804;
  assign N28814 = ~N28805;
  assign N28816 = ~N28806;
  assign N28818 = ~N28807;
  assign N28820 = ~N28808;
  assign N28822 = ~N28809;
  assign N28824 = ~N28810;
  assign N28826 = ~N28811;
  assign N28853 = ~commit_ack_i[1];
  assign N28854 = commit_ack_i[1];
  assign N28866 = ~N28858;
  assign N28868 = ~N28859;
  assign N28870 = ~N28860;
  assign N28872 = ~N28861;
  assign N28874 = ~N28862;
  assign N28876 = ~N28863;
  assign N28878 = ~N28864;
  assign N28880 = ~N28865;
  assign N28893 = ~N28885;
  assign N28895 = ~N28886;
  assign N28897 = ~N28887;
  assign N28899 = ~N28888;
  assign N28901 = ~N28889;
  assign N28903 = ~N28890;
  assign N28905 = ~N28891;
  assign N28907 = ~N28892;
  assign N28934 = ~flush_i;
  assign N28935 = ~mem_q[362];
  assign N28999 = ~N28936;
  assign N29004 = ~N28937;
  assign N29009 = ~N28938;
  assign N29014 = ~N28939;
  assign N29019 = ~N28940;
  assign N29024 = ~N28941;
  assign N29029 = ~N28942;
  assign N29034 = ~N28943;
  assign N29039 = ~N28944;
  assign N29044 = ~N28945;
  assign N29049 = ~N28946;
  assign N29054 = ~N28947;
  assign N29059 = ~N28948;
  assign N29064 = ~N28949;
  assign N29069 = ~N28950;
  assign N29074 = ~N28951;
  assign N29079 = ~N28952;
  assign N29084 = ~N28953;
  assign N29089 = ~N28954;
  assign N29094 = ~N28955;
  assign N29099 = ~N28956;
  assign N29104 = ~N28957;
  assign N29109 = ~N28958;
  assign N29114 = ~N28959;
  assign N29119 = ~N28960;
  assign N29124 = ~N28961;
  assign N29129 = ~N28962;
  assign N29134 = ~N28963;
  assign N29139 = ~N28964;
  assign N29144 = ~N28965;
  assign N29149 = ~N28966;
  assign N29154 = ~N28967;
  assign N29159 = ~N28968;
  assign N29164 = ~N28969;
  assign N29169 = ~N28970;
  assign N29174 = ~N28971;
  assign N29179 = ~N28972;
  assign N29184 = ~N28973;
  assign N29189 = ~N28974;
  assign N29194 = ~N28975;
  assign N29199 = ~N28976;
  assign N29204 = ~N28977;
  assign N29209 = ~N28978;
  assign N29214 = ~N28979;
  assign N29219 = ~N28980;
  assign N29224 = ~N28981;
  assign N29229 = ~N28982;
  assign N29234 = ~N28983;
  assign N29239 = ~N28984;
  assign N29244 = ~N28985;
  assign N29249 = ~N28986;
  assign N29254 = ~N28987;
  assign N29259 = ~N28988;
  assign N29264 = ~N28989;
  assign N29269 = ~N28990;
  assign N29274 = ~N28991;
  assign N29279 = ~N28992;
  assign N29284 = ~N28993;
  assign N29289 = ~N28994;
  assign N29294 = ~N28995;
  assign N29299 = ~N28996;
  assign N29304 = ~N28997;
  assign N29309 = ~N28998;
  assign N29566 = ~mem_q[725];
  assign N29630 = ~N29567;
  assign N29635 = ~N29568;
  assign N29640 = ~N29569;
  assign N29645 = ~N29570;
  assign N29650 = ~N29571;
  assign N29655 = ~N29572;
  assign N29660 = ~N29573;
  assign N29665 = ~N29574;
  assign N29670 = ~N29575;
  assign N29675 = ~N29576;
  assign N29680 = ~N29577;
  assign N29685 = ~N29578;
  assign N29690 = ~N29579;
  assign N29695 = ~N29580;
  assign N29700 = ~N29581;
  assign N29705 = ~N29582;
  assign N29710 = ~N29583;
  assign N29715 = ~N29584;
  assign N29720 = ~N29585;
  assign N29725 = ~N29586;
  assign N29730 = ~N29587;
  assign N29735 = ~N29588;
  assign N29740 = ~N29589;
  assign N29745 = ~N29590;
  assign N29750 = ~N29591;
  assign N29755 = ~N29592;
  assign N29760 = ~N29593;
  assign N29765 = ~N29594;
  assign N29770 = ~N29595;
  assign N29775 = ~N29596;
  assign N29780 = ~N29597;
  assign N29785 = ~N29598;
  assign N29790 = ~N29599;
  assign N29795 = ~N29600;
  assign N29800 = ~N29601;
  assign N29805 = ~N29602;
  assign N29810 = ~N29603;
  assign N29815 = ~N29604;
  assign N29820 = ~N29605;
  assign N29825 = ~N29606;
  assign N29830 = ~N29607;
  assign N29835 = ~N29608;
  assign N29840 = ~N29609;
  assign N29845 = ~N29610;
  assign N29850 = ~N29611;
  assign N29855 = ~N29612;
  assign N29860 = ~N29613;
  assign N29865 = ~N29614;
  assign N29870 = ~N29615;
  assign N29875 = ~N29616;
  assign N29880 = ~N29617;
  assign N29885 = ~N29618;
  assign N29890 = ~N29619;
  assign N29895 = ~N29620;
  assign N29900 = ~N29621;
  assign N29905 = ~N29622;
  assign N29910 = ~N29623;
  assign N29915 = ~N29624;
  assign N29920 = ~N29625;
  assign N29925 = ~N29626;
  assign N29930 = ~N29627;
  assign N29935 = ~N29628;
  assign N29940 = ~N29629;
  assign N30197 = ~mem_q[1088];
  assign N30261 = ~N30198;
  assign N30266 = ~N30199;
  assign N30271 = ~N30200;
  assign N30276 = ~N30201;
  assign N30281 = ~N30202;
  assign N30286 = ~N30203;
  assign N30291 = ~N30204;
  assign N30296 = ~N30205;
  assign N30301 = ~N30206;
  assign N30306 = ~N30207;
  assign N30311 = ~N30208;
  assign N30316 = ~N30209;
  assign N30321 = ~N30210;
  assign N30326 = ~N30211;
  assign N30331 = ~N30212;
  assign N30336 = ~N30213;
  assign N30341 = ~N30214;
  assign N30346 = ~N30215;
  assign N30351 = ~N30216;
  assign N30356 = ~N30217;
  assign N30361 = ~N30218;
  assign N30366 = ~N30219;
  assign N30371 = ~N30220;
  assign N30376 = ~N30221;
  assign N30381 = ~N30222;
  assign N30386 = ~N30223;
  assign N30391 = ~N30224;
  assign N30396 = ~N30225;
  assign N30401 = ~N30226;
  assign N30406 = ~N30227;
  assign N30411 = ~N30228;
  assign N30416 = ~N30229;
  assign N30421 = ~N30230;
  assign N30426 = ~N30231;
  assign N30431 = ~N30232;
  assign N30436 = ~N30233;
  assign N30441 = ~N30234;
  assign N30446 = ~N30235;
  assign N30451 = ~N30236;
  assign N30456 = ~N30237;
  assign N30461 = ~N30238;
  assign N30466 = ~N30239;
  assign N30471 = ~N30240;
  assign N30476 = ~N30241;
  assign N30481 = ~N30242;
  assign N30486 = ~N30243;
  assign N30491 = ~N30244;
  assign N30496 = ~N30245;
  assign N30501 = ~N30246;
  assign N30506 = ~N30247;
  assign N30511 = ~N30248;
  assign N30516 = ~N30249;
  assign N30521 = ~N30250;
  assign N30526 = ~N30251;
  assign N30531 = ~N30252;
  assign N30536 = ~N30253;
  assign N30541 = ~N30254;
  assign N30546 = ~N30255;
  assign N30551 = ~N30256;
  assign N30556 = ~N30257;
  assign N30561 = ~N30258;
  assign N30566 = ~N30259;
  assign N30571 = ~N30260;
  assign N30828 = ~mem_q[1451];
  assign N30892 = ~N30829;
  assign N30897 = ~N30830;
  assign N30902 = ~N30831;
  assign N30907 = ~N30832;
  assign N30912 = ~N30833;
  assign N30917 = ~N30834;
  assign N30922 = ~N30835;
  assign N30927 = ~N30836;
  assign N30932 = ~N30837;
  assign N30937 = ~N30838;
  assign N30942 = ~N30839;
  assign N30947 = ~N30840;
  assign N30952 = ~N30841;
  assign N30957 = ~N30842;
  assign N30962 = ~N30843;
  assign N30967 = ~N30844;
  assign N30972 = ~N30845;
  assign N30977 = ~N30846;
  assign N30982 = ~N30847;
  assign N30987 = ~N30848;
  assign N30992 = ~N30849;
  assign N30997 = ~N30850;
  assign N31002 = ~N30851;
  assign N31007 = ~N30852;
  assign N31012 = ~N30853;
  assign N31017 = ~N30854;
  assign N31022 = ~N30855;
  assign N31027 = ~N30856;
  assign N31032 = ~N30857;
  assign N31037 = ~N30858;
  assign N31042 = ~N30859;
  assign N31047 = ~N30860;
  assign N31052 = ~N30861;
  assign N31057 = ~N30862;
  assign N31062 = ~N30863;
  assign N31067 = ~N30864;
  assign N31072 = ~N30865;
  assign N31077 = ~N30866;
  assign N31082 = ~N30867;
  assign N31087 = ~N30868;
  assign N31092 = ~N30869;
  assign N31097 = ~N30870;
  assign N31102 = ~N30871;
  assign N31107 = ~N30872;
  assign N31112 = ~N30873;
  assign N31117 = ~N30874;
  assign N31122 = ~N30875;
  assign N31127 = ~N30876;
  assign N31132 = ~N30877;
  assign N31137 = ~N30878;
  assign N31142 = ~N30879;
  assign N31147 = ~N30880;
  assign N31152 = ~N30881;
  assign N31157 = ~N30882;
  assign N31162 = ~N30883;
  assign N31167 = ~N30884;
  assign N31172 = ~N30885;
  assign N31177 = ~N30886;
  assign N31182 = ~N30887;
  assign N31187 = ~N30888;
  assign N31192 = ~N30889;
  assign N31197 = ~N30890;
  assign N31202 = ~N30891;
  assign N31459 = ~mem_q[1814];
  assign N31523 = ~N31460;
  assign N31528 = ~N31461;
  assign N31533 = ~N31462;
  assign N31538 = ~N31463;
  assign N31543 = ~N31464;
  assign N31548 = ~N31465;
  assign N31553 = ~N31466;
  assign N31558 = ~N31467;
  assign N31563 = ~N31468;
  assign N31568 = ~N31469;
  assign N31573 = ~N31470;
  assign N31578 = ~N31471;
  assign N31583 = ~N31472;
  assign N31588 = ~N31473;
  assign N31593 = ~N31474;
  assign N31598 = ~N31475;
  assign N31603 = ~N31476;
  assign N31608 = ~N31477;
  assign N31613 = ~N31478;
  assign N31618 = ~N31479;
  assign N31623 = ~N31480;
  assign N31628 = ~N31481;
  assign N31633 = ~N31482;
  assign N31638 = ~N31483;
  assign N31643 = ~N31484;
  assign N31648 = ~N31485;
  assign N31653 = ~N31486;
  assign N31658 = ~N31487;
  assign N31663 = ~N31488;
  assign N31668 = ~N31489;
  assign N31673 = ~N31490;
  assign N31678 = ~N31491;
  assign N31683 = ~N31492;
  assign N31688 = ~N31493;
  assign N31693 = ~N31494;
  assign N31698 = ~N31495;
  assign N31703 = ~N31496;
  assign N31708 = ~N31497;
  assign N31713 = ~N31498;
  assign N31718 = ~N31499;
  assign N31723 = ~N31500;
  assign N31728 = ~N31501;
  assign N31733 = ~N31502;
  assign N31738 = ~N31503;
  assign N31743 = ~N31504;
  assign N31748 = ~N31505;
  assign N31753 = ~N31506;
  assign N31758 = ~N31507;
  assign N31763 = ~N31508;
  assign N31768 = ~N31509;
  assign N31773 = ~N31510;
  assign N31778 = ~N31511;
  assign N31783 = ~N31512;
  assign N31788 = ~N31513;
  assign N31793 = ~N31514;
  assign N31798 = ~N31515;
  assign N31803 = ~N31516;
  assign N31808 = ~N31517;
  assign N31813 = ~N31518;
  assign N31818 = ~N31519;
  assign N31823 = ~N31520;
  assign N31828 = ~N31521;
  assign N31833 = ~N31522;
  assign N32090 = ~mem_q[2177];
  assign N32154 = ~N32091;
  assign N32159 = ~N32092;
  assign N32164 = ~N32093;
  assign N32169 = ~N32094;
  assign N32174 = ~N32095;
  assign N32179 = ~N32096;
  assign N32184 = ~N32097;
  assign N32189 = ~N32098;
  assign N32194 = ~N32099;
  assign N32199 = ~N32100;
  assign N32204 = ~N32101;
  assign N32209 = ~N32102;
  assign N32214 = ~N32103;
  assign N32219 = ~N32104;
  assign N32224 = ~N32105;
  assign N32229 = ~N32106;
  assign N32234 = ~N32107;
  assign N32239 = ~N32108;
  assign N32244 = ~N32109;
  assign N32249 = ~N32110;
  assign N32254 = ~N32111;
  assign N32259 = ~N32112;
  assign N32264 = ~N32113;
  assign N32269 = ~N32114;
  assign N32274 = ~N32115;
  assign N32279 = ~N32116;
  assign N32284 = ~N32117;
  assign N32289 = ~N32118;
  assign N32294 = ~N32119;
  assign N32299 = ~N32120;
  assign N32304 = ~N32121;
  assign N32309 = ~N32122;
  assign N32314 = ~N32123;
  assign N32319 = ~N32124;
  assign N32324 = ~N32125;
  assign N32329 = ~N32126;
  assign N32334 = ~N32127;
  assign N32339 = ~N32128;
  assign N32344 = ~N32129;
  assign N32349 = ~N32130;
  assign N32354 = ~N32131;
  assign N32359 = ~N32132;
  assign N32364 = ~N32133;
  assign N32369 = ~N32134;
  assign N32374 = ~N32135;
  assign N32379 = ~N32136;
  assign N32384 = ~N32137;
  assign N32389 = ~N32138;
  assign N32394 = ~N32139;
  assign N32399 = ~N32140;
  assign N32404 = ~N32141;
  assign N32409 = ~N32142;
  assign N32414 = ~N32143;
  assign N32419 = ~N32144;
  assign N32424 = ~N32145;
  assign N32429 = ~N32146;
  assign N32434 = ~N32147;
  assign N32439 = ~N32148;
  assign N32444 = ~N32149;
  assign N32449 = ~N32150;
  assign N32454 = ~N32151;
  assign N32459 = ~N32152;
  assign N32464 = ~N32153;
  assign N32721 = ~mem_q[2540];
  assign N32785 = ~N32722;
  assign N32790 = ~N32723;
  assign N32795 = ~N32724;
  assign N32800 = ~N32725;
  assign N32805 = ~N32726;
  assign N32810 = ~N32727;
  assign N32815 = ~N32728;
  assign N32820 = ~N32729;
  assign N32825 = ~N32730;
  assign N32830 = ~N32731;
  assign N32835 = ~N32732;
  assign N32840 = ~N32733;
  assign N32845 = ~N32734;
  assign N32850 = ~N32735;
  assign N32855 = ~N32736;
  assign N32860 = ~N32737;
  assign N32865 = ~N32738;
  assign N32870 = ~N32739;
  assign N32875 = ~N32740;
  assign N32880 = ~N32741;
  assign N32885 = ~N32742;
  assign N32890 = ~N32743;
  assign N32895 = ~N32744;
  assign N32900 = ~N32745;
  assign N32905 = ~N32746;
  assign N32910 = ~N32747;
  assign N32915 = ~N32748;
  assign N32920 = ~N32749;
  assign N32925 = ~N32750;
  assign N32930 = ~N32751;
  assign N32935 = ~N32752;
  assign N32940 = ~N32753;
  assign N32945 = ~N32754;
  assign N32950 = ~N32755;
  assign N32955 = ~N32756;
  assign N32960 = ~N32757;
  assign N32965 = ~N32758;
  assign N32970 = ~N32759;
  assign N32975 = ~N32760;
  assign N32980 = ~N32761;
  assign N32985 = ~N32762;
  assign N32990 = ~N32763;
  assign N32995 = ~N32764;
  assign N33000 = ~N32765;
  assign N33005 = ~N32766;
  assign N33010 = ~N32767;
  assign N33015 = ~N32768;
  assign N33020 = ~N32769;
  assign N33025 = ~N32770;
  assign N33030 = ~N32771;
  assign N33035 = ~N32772;
  assign N33040 = ~N32773;
  assign N33045 = ~N32774;
  assign N33050 = ~N32775;
  assign N33055 = ~N32776;
  assign N33060 = ~N32777;
  assign N33065 = ~N32778;
  assign N33070 = ~N32779;
  assign N33075 = ~N32780;
  assign N33080 = ~N32781;
  assign N33085 = ~N32782;
  assign N33090 = ~N32783;
  assign N33095 = ~N32784;
  assign N33352 = ~mem_q[2903];
  assign N33416 = ~N33353;
  assign N33421 = ~N33354;
  assign N33426 = ~N33355;
  assign N33431 = ~N33356;
  assign N33436 = ~N33357;
  assign N33441 = ~N33358;
  assign N33446 = ~N33359;
  assign N33451 = ~N33360;
  assign N33456 = ~N33361;
  assign N33461 = ~N33362;
  assign N33466 = ~N33363;
  assign N33471 = ~N33364;
  assign N33476 = ~N33365;
  assign N33481 = ~N33366;
  assign N33486 = ~N33367;
  assign N33491 = ~N33368;
  assign N33496 = ~N33369;
  assign N33501 = ~N33370;
  assign N33506 = ~N33371;
  assign N33511 = ~N33372;
  assign N33516 = ~N33373;
  assign N33521 = ~N33374;
  assign N33526 = ~N33375;
  assign N33531 = ~N33376;
  assign N33536 = ~N33377;
  assign N33541 = ~N33378;
  assign N33546 = ~N33379;
  assign N33551 = ~N33380;
  assign N33556 = ~N33381;
  assign N33561 = ~N33382;
  assign N33566 = ~N33383;
  assign N33571 = ~N33384;
  assign N33576 = ~N33385;
  assign N33581 = ~N33386;
  assign N33586 = ~N33387;
  assign N33591 = ~N33388;
  assign N33596 = ~N33389;
  assign N33601 = ~N33390;
  assign N33606 = ~N33391;
  assign N33611 = ~N33392;
  assign N33616 = ~N33393;
  assign N33621 = ~N33394;
  assign N33626 = ~N33395;
  assign N33631 = ~N33396;
  assign N33636 = ~N33397;
  assign N33641 = ~N33398;
  assign N33646 = ~N33399;
  assign N33651 = ~N33400;
  assign N33656 = ~N33401;
  assign N33661 = ~N33402;
  assign N33666 = ~N33403;
  assign N33671 = ~N33404;
  assign N33676 = ~N33405;
  assign N33681 = ~N33406;
  assign N33686 = ~N33407;
  assign N33691 = ~N33408;
  assign N33696 = ~N33409;
  assign N33701 = ~N33410;
  assign N33706 = ~N33411;
  assign N33711 = ~N33412;
  assign N33716 = ~N33413;
  assign N33721 = ~N33414;
  assign N33726 = ~N33415;
  assign N33731 = mem_q[362];
  assign N33733 = ~N33732;
  assign N33734 = N33731 & N33733;
  assign N33736 = ~N33735;
  assign N33738 = ~N33737;
  assign N34076 = mem_q[725];
  assign N34078 = ~N34077;
  assign N34079 = N34076 & N34078;
  assign N34081 = ~N34080;
  assign N34083 = ~N34082;
  assign N34421 = mem_q[1088];
  assign N34423 = ~N34422;
  assign N34424 = N34421 & N34423;
  assign N34426 = ~N34425;
  assign N34428 = ~N34427;
  assign N34766 = mem_q[1451];
  assign N34768 = ~N34767;
  assign N34769 = N34766 & N34768;
  assign N34771 = ~N34770;
  assign N34773 = ~N34772;
  assign N35111 = mem_q[1814];
  assign N35113 = ~N35112;
  assign N35114 = N35111 & N35113;
  assign N35116 = ~N35115;
  assign N35118 = ~N35117;
  assign N35456 = mem_q[2177];
  assign N35458 = ~N35457;
  assign N35459 = N35456 & N35458;
  assign N35461 = ~N35460;
  assign N35463 = ~N35462;
  assign N35801 = mem_q[2540];
  assign N35803 = ~N35802;
  assign N35804 = N35801 & N35803;
  assign N35806 = ~N35805;
  assign N35808 = ~N35807;
  assign N36146 = mem_q[2903];
  assign N36148 = ~N36147;
  assign N36149 = N36146 & N36148;
  assign N36151 = ~N36150;
  assign N36153 = ~N36152;
  assign N36497 = ~ex_i[0];
  assign N36499 = N38944 & N36497;
  assign N38944 = N36498 & wb_valid_i[0];
  assign N36500 = ~N36499;
  assign N36566 = N36500;
  assign N36568 = N38945 & N36497;
  assign N38945 = N36567 & wb_valid_i[0];
  assign N36569 = ~N36568;
  assign N36636 = ~N36635;
  assign N36637 = N36566 & N36635;
  assign N36639 = N38946 & N36497;
  assign N38946 = N36638 & wb_valid_i[0];
  assign N36640 = ~N36639;
  assign N36645 = ~N36644;
  assign N36646 = N36637 & N36644;
  assign N36647 = N36646 & N36644;
  assign N36654 = ~ex_i[129];
  assign N36656 = N38947 & N36654;
  assign N38947 = N36655 & wb_valid_i[1];
  assign N36657 = ~N36656;
  assign N36724 = ~N36723;
  assign N36725 = N36647 & N36723;
  assign N36727 = N38948 & N36654;
  assign N38948 = N36726 & wb_valid_i[1];
  assign N36728 = ~N36727;
  assign N36795 = ~N36794;
  assign N36796 = N36725 & N36794;
  assign N36798 = N38949 & N36654;
  assign N38949 = N36797 & wb_valid_i[1];
  assign N36799 = ~N36798;
  assign N36804 = ~N36803;
  assign N36805 = N36796 & N36803;
  assign N36806 = N36805 & N36803;
  assign N36813 = ~ex_i[258];
  assign N36815 = N38950 & N36813;
  assign N38950 = N36814 & wb_valid_i[2];
  assign N36816 = ~N36815;
  assign N36883 = ~N36882;
  assign N36884 = N36806 & N36882;
  assign N36886 = N38951 & N36813;
  assign N38951 = N36885 & wb_valid_i[2];
  assign N36887 = ~N36886;
  assign N36954 = ~N36953;
  assign N36955 = N36884 & N36953;
  assign N36957 = N38952 & N36813;
  assign N38952 = N36956 & wb_valid_i[2];
  assign N36958 = ~N36957;
  assign N36963 = ~N36962;
  assign N36964 = N36955 & N36962;
  assign N36965 = N36964 & N36962;
  assign N36972 = ~ex_i[387];
  assign N36974 = N38953 & N36972;
  assign N38953 = N36973 & wb_valid_i[3];
  assign N36975 = ~N36974;
  assign N37042 = ~N37041;
  assign N37043 = N36965 & N37041;
  assign N37045 = N38954 & N36972;
  assign N38954 = N37044 & wb_valid_i[3];
  assign N37046 = ~N37045;
  assign N37113 = ~N37112;
  assign N37115 = N38955 & N36972;
  assign N38955 = N37114 & wb_valid_i[3];
  assign N37116 = ~N37115;
  assign N37191 = ~N36962;
  assign N37724 = ~N36803;
  assign N38257 = ~N36644;
  assign N38659 = ~rst_ni;
  assign N38660 = N884 & N28934;
  assign N38661 = ~N38660;

endmodule