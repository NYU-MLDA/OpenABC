module bsg_mux_one_hot_width_p539_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [2694:0] data_i;
  input [4:0] sel_one_hot_i;
  output [538:0] data_o;
  wire [538:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616;
  wire [2694:0] data_masked;
  assign data_masked[538] = data_i[538] & sel_one_hot_i[0];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[0];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[0];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[0];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[0];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[0];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[0];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[0];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[0];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[0];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[0];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[0];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[0];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[0];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[0];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[0];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[0];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[0];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[0];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[0];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[0];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[0];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[0];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[0];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[0];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[0];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[0];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[0];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[0];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[0];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[0];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[0];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[0];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[0];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[0];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[0];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[0];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[0];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[0];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[0];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[0];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[0];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[0];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[0];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[0];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[0];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[0];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[0];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[0];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[0];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[0];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[0];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[0];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[0];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[0];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[0];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[0];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[0];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[0];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[0];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[0];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[0];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[0];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[0];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[0];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[0];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[0];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[0];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[0];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[0];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[0];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[0];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[0];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[0];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[0];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[0];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[0];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[0];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[0];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[0];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[0];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[0];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[0];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[0];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[0];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[0];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[0];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[0];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[0];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[0];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[0];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[0];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[0];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[0];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[0];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[0];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[0];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[0];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[0];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[0];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[0];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[0];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[0];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[0];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[0];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[0];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[0];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[0];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[0];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[0];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[0];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[0];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[0];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[0];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[0];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[0];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[0];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[0];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[0];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[0];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[0];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[0];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[0];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[0];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[0];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[0];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[0];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[0];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[0];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[0];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[0];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[0];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[0];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[0];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[0];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[0];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[0];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[0];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[0];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[0];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[0];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[0];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[0];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[0];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[0];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[0];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[0];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[0];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[0];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[0];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[0];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[0];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[0];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[0];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[0];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[0];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[0];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[0];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[0];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[0];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[0];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[0];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[0];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[0];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[0];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[0];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[0];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[0];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[0];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[0];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[0];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[0];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[0];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[0];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[0];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[0];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[0];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[0];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[0];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[0];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[0];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[0];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[0];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[0];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[0];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[0];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[0];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[0];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[0];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[0];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[0];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[0];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[0];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[0];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[0];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[0];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[0];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[0];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[0];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[0];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[0];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[0];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[0];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[0];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[0];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[0];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[0];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[0];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[0];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[0];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[0];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[0];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[0];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[0];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[0];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[0];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[0];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[0];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[0];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[0];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[0];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[0];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[0];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[0];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[0];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[0];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[0];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[0];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[0];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[0];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[0];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[0];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[0];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[0];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[0];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[0];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[0];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[0];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[0];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[0];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[0];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[0];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[0];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[0];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[0];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[0];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[0];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[0];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[0];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[0];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[0];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[0];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[0];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[0];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[0];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[0];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[0];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[0];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[0];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[0];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[0];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[0];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[0];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[0];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[0];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[0];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[0];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[0];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[0];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[0];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[0];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[0];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[0];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[0];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[0];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[0];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[0];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[0];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[0];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[0];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[0];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[0];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[0];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[0];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[0];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[0];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[0];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[0];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[0];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[0];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[0];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[0];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[0];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[0];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[0];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[0];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[0];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[0];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[0];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[0];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[0];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[0];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[0];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[0];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[0];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[0];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[0];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[0];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[0];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[0];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[0];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[0];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[0];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[0];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[0];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[0];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[0];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[0];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[0];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[0];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[0];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[0];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[0];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[0];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[0];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[0];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[0];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[0];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[0];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[0];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[0];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[0];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[0];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[0];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[0];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[0];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[0];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[0];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[0];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[0];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[0];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[0];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[0];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[0];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[0];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[0];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[0];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[0];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[0];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[0];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[0];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[0];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[0];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[0];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[0];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[0];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[0];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[0];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[0];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[0];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[0];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[0];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[0];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[0];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[0];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[0];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[0];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[0];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[0];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[0];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[0];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[0];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[0];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[0];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[0];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[0];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[0];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[0];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[0];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[0];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[0];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[0];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[0];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[0];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[0];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[0];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[0];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[0];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[0];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[0];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[0];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[0];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[0];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[0];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[0];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[0];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[0];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[0];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[0];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[0];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[0];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[0];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[0];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[0];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[0];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[0];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[0];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[0];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[0];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[1077] = data_i[1077] & sel_one_hot_i[1];
  assign data_masked[1076] = data_i[1076] & sel_one_hot_i[1];
  assign data_masked[1075] = data_i[1075] & sel_one_hot_i[1];
  assign data_masked[1074] = data_i[1074] & sel_one_hot_i[1];
  assign data_masked[1073] = data_i[1073] & sel_one_hot_i[1];
  assign data_masked[1072] = data_i[1072] & sel_one_hot_i[1];
  assign data_masked[1071] = data_i[1071] & sel_one_hot_i[1];
  assign data_masked[1070] = data_i[1070] & sel_one_hot_i[1];
  assign data_masked[1069] = data_i[1069] & sel_one_hot_i[1];
  assign data_masked[1068] = data_i[1068] & sel_one_hot_i[1];
  assign data_masked[1067] = data_i[1067] & sel_one_hot_i[1];
  assign data_masked[1066] = data_i[1066] & sel_one_hot_i[1];
  assign data_masked[1065] = data_i[1065] & sel_one_hot_i[1];
  assign data_masked[1064] = data_i[1064] & sel_one_hot_i[1];
  assign data_masked[1063] = data_i[1063] & sel_one_hot_i[1];
  assign data_masked[1062] = data_i[1062] & sel_one_hot_i[1];
  assign data_masked[1061] = data_i[1061] & sel_one_hot_i[1];
  assign data_masked[1060] = data_i[1060] & sel_one_hot_i[1];
  assign data_masked[1059] = data_i[1059] & sel_one_hot_i[1];
  assign data_masked[1058] = data_i[1058] & sel_one_hot_i[1];
  assign data_masked[1057] = data_i[1057] & sel_one_hot_i[1];
  assign data_masked[1056] = data_i[1056] & sel_one_hot_i[1];
  assign data_masked[1055] = data_i[1055] & sel_one_hot_i[1];
  assign data_masked[1054] = data_i[1054] & sel_one_hot_i[1];
  assign data_masked[1053] = data_i[1053] & sel_one_hot_i[1];
  assign data_masked[1052] = data_i[1052] & sel_one_hot_i[1];
  assign data_masked[1051] = data_i[1051] & sel_one_hot_i[1];
  assign data_masked[1050] = data_i[1050] & sel_one_hot_i[1];
  assign data_masked[1049] = data_i[1049] & sel_one_hot_i[1];
  assign data_masked[1048] = data_i[1048] & sel_one_hot_i[1];
  assign data_masked[1047] = data_i[1047] & sel_one_hot_i[1];
  assign data_masked[1046] = data_i[1046] & sel_one_hot_i[1];
  assign data_masked[1045] = data_i[1045] & sel_one_hot_i[1];
  assign data_masked[1044] = data_i[1044] & sel_one_hot_i[1];
  assign data_masked[1043] = data_i[1043] & sel_one_hot_i[1];
  assign data_masked[1042] = data_i[1042] & sel_one_hot_i[1];
  assign data_masked[1041] = data_i[1041] & sel_one_hot_i[1];
  assign data_masked[1040] = data_i[1040] & sel_one_hot_i[1];
  assign data_masked[1039] = data_i[1039] & sel_one_hot_i[1];
  assign data_masked[1038] = data_i[1038] & sel_one_hot_i[1];
  assign data_masked[1037] = data_i[1037] & sel_one_hot_i[1];
  assign data_masked[1036] = data_i[1036] & sel_one_hot_i[1];
  assign data_masked[1035] = data_i[1035] & sel_one_hot_i[1];
  assign data_masked[1034] = data_i[1034] & sel_one_hot_i[1];
  assign data_masked[1033] = data_i[1033] & sel_one_hot_i[1];
  assign data_masked[1032] = data_i[1032] & sel_one_hot_i[1];
  assign data_masked[1031] = data_i[1031] & sel_one_hot_i[1];
  assign data_masked[1030] = data_i[1030] & sel_one_hot_i[1];
  assign data_masked[1029] = data_i[1029] & sel_one_hot_i[1];
  assign data_masked[1028] = data_i[1028] & sel_one_hot_i[1];
  assign data_masked[1027] = data_i[1027] & sel_one_hot_i[1];
  assign data_masked[1026] = data_i[1026] & sel_one_hot_i[1];
  assign data_masked[1025] = data_i[1025] & sel_one_hot_i[1];
  assign data_masked[1024] = data_i[1024] & sel_one_hot_i[1];
  assign data_masked[1023] = data_i[1023] & sel_one_hot_i[1];
  assign data_masked[1022] = data_i[1022] & sel_one_hot_i[1];
  assign data_masked[1021] = data_i[1021] & sel_one_hot_i[1];
  assign data_masked[1020] = data_i[1020] & sel_one_hot_i[1];
  assign data_masked[1019] = data_i[1019] & sel_one_hot_i[1];
  assign data_masked[1018] = data_i[1018] & sel_one_hot_i[1];
  assign data_masked[1017] = data_i[1017] & sel_one_hot_i[1];
  assign data_masked[1016] = data_i[1016] & sel_one_hot_i[1];
  assign data_masked[1015] = data_i[1015] & sel_one_hot_i[1];
  assign data_masked[1014] = data_i[1014] & sel_one_hot_i[1];
  assign data_masked[1013] = data_i[1013] & sel_one_hot_i[1];
  assign data_masked[1012] = data_i[1012] & sel_one_hot_i[1];
  assign data_masked[1011] = data_i[1011] & sel_one_hot_i[1];
  assign data_masked[1010] = data_i[1010] & sel_one_hot_i[1];
  assign data_masked[1009] = data_i[1009] & sel_one_hot_i[1];
  assign data_masked[1008] = data_i[1008] & sel_one_hot_i[1];
  assign data_masked[1007] = data_i[1007] & sel_one_hot_i[1];
  assign data_masked[1006] = data_i[1006] & sel_one_hot_i[1];
  assign data_masked[1005] = data_i[1005] & sel_one_hot_i[1];
  assign data_masked[1004] = data_i[1004] & sel_one_hot_i[1];
  assign data_masked[1003] = data_i[1003] & sel_one_hot_i[1];
  assign data_masked[1002] = data_i[1002] & sel_one_hot_i[1];
  assign data_masked[1001] = data_i[1001] & sel_one_hot_i[1];
  assign data_masked[1000] = data_i[1000] & sel_one_hot_i[1];
  assign data_masked[999] = data_i[999] & sel_one_hot_i[1];
  assign data_masked[998] = data_i[998] & sel_one_hot_i[1];
  assign data_masked[997] = data_i[997] & sel_one_hot_i[1];
  assign data_masked[996] = data_i[996] & sel_one_hot_i[1];
  assign data_masked[995] = data_i[995] & sel_one_hot_i[1];
  assign data_masked[994] = data_i[994] & sel_one_hot_i[1];
  assign data_masked[993] = data_i[993] & sel_one_hot_i[1];
  assign data_masked[992] = data_i[992] & sel_one_hot_i[1];
  assign data_masked[991] = data_i[991] & sel_one_hot_i[1];
  assign data_masked[990] = data_i[990] & sel_one_hot_i[1];
  assign data_masked[989] = data_i[989] & sel_one_hot_i[1];
  assign data_masked[988] = data_i[988] & sel_one_hot_i[1];
  assign data_masked[987] = data_i[987] & sel_one_hot_i[1];
  assign data_masked[986] = data_i[986] & sel_one_hot_i[1];
  assign data_masked[985] = data_i[985] & sel_one_hot_i[1];
  assign data_masked[984] = data_i[984] & sel_one_hot_i[1];
  assign data_masked[983] = data_i[983] & sel_one_hot_i[1];
  assign data_masked[982] = data_i[982] & sel_one_hot_i[1];
  assign data_masked[981] = data_i[981] & sel_one_hot_i[1];
  assign data_masked[980] = data_i[980] & sel_one_hot_i[1];
  assign data_masked[979] = data_i[979] & sel_one_hot_i[1];
  assign data_masked[978] = data_i[978] & sel_one_hot_i[1];
  assign data_masked[977] = data_i[977] & sel_one_hot_i[1];
  assign data_masked[976] = data_i[976] & sel_one_hot_i[1];
  assign data_masked[975] = data_i[975] & sel_one_hot_i[1];
  assign data_masked[974] = data_i[974] & sel_one_hot_i[1];
  assign data_masked[973] = data_i[973] & sel_one_hot_i[1];
  assign data_masked[972] = data_i[972] & sel_one_hot_i[1];
  assign data_masked[971] = data_i[971] & sel_one_hot_i[1];
  assign data_masked[970] = data_i[970] & sel_one_hot_i[1];
  assign data_masked[969] = data_i[969] & sel_one_hot_i[1];
  assign data_masked[968] = data_i[968] & sel_one_hot_i[1];
  assign data_masked[967] = data_i[967] & sel_one_hot_i[1];
  assign data_masked[966] = data_i[966] & sel_one_hot_i[1];
  assign data_masked[965] = data_i[965] & sel_one_hot_i[1];
  assign data_masked[964] = data_i[964] & sel_one_hot_i[1];
  assign data_masked[963] = data_i[963] & sel_one_hot_i[1];
  assign data_masked[962] = data_i[962] & sel_one_hot_i[1];
  assign data_masked[961] = data_i[961] & sel_one_hot_i[1];
  assign data_masked[960] = data_i[960] & sel_one_hot_i[1];
  assign data_masked[959] = data_i[959] & sel_one_hot_i[1];
  assign data_masked[958] = data_i[958] & sel_one_hot_i[1];
  assign data_masked[957] = data_i[957] & sel_one_hot_i[1];
  assign data_masked[956] = data_i[956] & sel_one_hot_i[1];
  assign data_masked[955] = data_i[955] & sel_one_hot_i[1];
  assign data_masked[954] = data_i[954] & sel_one_hot_i[1];
  assign data_masked[953] = data_i[953] & sel_one_hot_i[1];
  assign data_masked[952] = data_i[952] & sel_one_hot_i[1];
  assign data_masked[951] = data_i[951] & sel_one_hot_i[1];
  assign data_masked[950] = data_i[950] & sel_one_hot_i[1];
  assign data_masked[949] = data_i[949] & sel_one_hot_i[1];
  assign data_masked[948] = data_i[948] & sel_one_hot_i[1];
  assign data_masked[947] = data_i[947] & sel_one_hot_i[1];
  assign data_masked[946] = data_i[946] & sel_one_hot_i[1];
  assign data_masked[945] = data_i[945] & sel_one_hot_i[1];
  assign data_masked[944] = data_i[944] & sel_one_hot_i[1];
  assign data_masked[943] = data_i[943] & sel_one_hot_i[1];
  assign data_masked[942] = data_i[942] & sel_one_hot_i[1];
  assign data_masked[941] = data_i[941] & sel_one_hot_i[1];
  assign data_masked[940] = data_i[940] & sel_one_hot_i[1];
  assign data_masked[939] = data_i[939] & sel_one_hot_i[1];
  assign data_masked[938] = data_i[938] & sel_one_hot_i[1];
  assign data_masked[937] = data_i[937] & sel_one_hot_i[1];
  assign data_masked[936] = data_i[936] & sel_one_hot_i[1];
  assign data_masked[935] = data_i[935] & sel_one_hot_i[1];
  assign data_masked[934] = data_i[934] & sel_one_hot_i[1];
  assign data_masked[933] = data_i[933] & sel_one_hot_i[1];
  assign data_masked[932] = data_i[932] & sel_one_hot_i[1];
  assign data_masked[931] = data_i[931] & sel_one_hot_i[1];
  assign data_masked[930] = data_i[930] & sel_one_hot_i[1];
  assign data_masked[929] = data_i[929] & sel_one_hot_i[1];
  assign data_masked[928] = data_i[928] & sel_one_hot_i[1];
  assign data_masked[927] = data_i[927] & sel_one_hot_i[1];
  assign data_masked[926] = data_i[926] & sel_one_hot_i[1];
  assign data_masked[925] = data_i[925] & sel_one_hot_i[1];
  assign data_masked[924] = data_i[924] & sel_one_hot_i[1];
  assign data_masked[923] = data_i[923] & sel_one_hot_i[1];
  assign data_masked[922] = data_i[922] & sel_one_hot_i[1];
  assign data_masked[921] = data_i[921] & sel_one_hot_i[1];
  assign data_masked[920] = data_i[920] & sel_one_hot_i[1];
  assign data_masked[919] = data_i[919] & sel_one_hot_i[1];
  assign data_masked[918] = data_i[918] & sel_one_hot_i[1];
  assign data_masked[917] = data_i[917] & sel_one_hot_i[1];
  assign data_masked[916] = data_i[916] & sel_one_hot_i[1];
  assign data_masked[915] = data_i[915] & sel_one_hot_i[1];
  assign data_masked[914] = data_i[914] & sel_one_hot_i[1];
  assign data_masked[913] = data_i[913] & sel_one_hot_i[1];
  assign data_masked[912] = data_i[912] & sel_one_hot_i[1];
  assign data_masked[911] = data_i[911] & sel_one_hot_i[1];
  assign data_masked[910] = data_i[910] & sel_one_hot_i[1];
  assign data_masked[909] = data_i[909] & sel_one_hot_i[1];
  assign data_masked[908] = data_i[908] & sel_one_hot_i[1];
  assign data_masked[907] = data_i[907] & sel_one_hot_i[1];
  assign data_masked[906] = data_i[906] & sel_one_hot_i[1];
  assign data_masked[905] = data_i[905] & sel_one_hot_i[1];
  assign data_masked[904] = data_i[904] & sel_one_hot_i[1];
  assign data_masked[903] = data_i[903] & sel_one_hot_i[1];
  assign data_masked[902] = data_i[902] & sel_one_hot_i[1];
  assign data_masked[901] = data_i[901] & sel_one_hot_i[1];
  assign data_masked[900] = data_i[900] & sel_one_hot_i[1];
  assign data_masked[899] = data_i[899] & sel_one_hot_i[1];
  assign data_masked[898] = data_i[898] & sel_one_hot_i[1];
  assign data_masked[897] = data_i[897] & sel_one_hot_i[1];
  assign data_masked[896] = data_i[896] & sel_one_hot_i[1];
  assign data_masked[895] = data_i[895] & sel_one_hot_i[1];
  assign data_masked[894] = data_i[894] & sel_one_hot_i[1];
  assign data_masked[893] = data_i[893] & sel_one_hot_i[1];
  assign data_masked[892] = data_i[892] & sel_one_hot_i[1];
  assign data_masked[891] = data_i[891] & sel_one_hot_i[1];
  assign data_masked[890] = data_i[890] & sel_one_hot_i[1];
  assign data_masked[889] = data_i[889] & sel_one_hot_i[1];
  assign data_masked[888] = data_i[888] & sel_one_hot_i[1];
  assign data_masked[887] = data_i[887] & sel_one_hot_i[1];
  assign data_masked[886] = data_i[886] & sel_one_hot_i[1];
  assign data_masked[885] = data_i[885] & sel_one_hot_i[1];
  assign data_masked[884] = data_i[884] & sel_one_hot_i[1];
  assign data_masked[883] = data_i[883] & sel_one_hot_i[1];
  assign data_masked[882] = data_i[882] & sel_one_hot_i[1];
  assign data_masked[881] = data_i[881] & sel_one_hot_i[1];
  assign data_masked[880] = data_i[880] & sel_one_hot_i[1];
  assign data_masked[879] = data_i[879] & sel_one_hot_i[1];
  assign data_masked[878] = data_i[878] & sel_one_hot_i[1];
  assign data_masked[877] = data_i[877] & sel_one_hot_i[1];
  assign data_masked[876] = data_i[876] & sel_one_hot_i[1];
  assign data_masked[875] = data_i[875] & sel_one_hot_i[1];
  assign data_masked[874] = data_i[874] & sel_one_hot_i[1];
  assign data_masked[873] = data_i[873] & sel_one_hot_i[1];
  assign data_masked[872] = data_i[872] & sel_one_hot_i[1];
  assign data_masked[871] = data_i[871] & sel_one_hot_i[1];
  assign data_masked[870] = data_i[870] & sel_one_hot_i[1];
  assign data_masked[869] = data_i[869] & sel_one_hot_i[1];
  assign data_masked[868] = data_i[868] & sel_one_hot_i[1];
  assign data_masked[867] = data_i[867] & sel_one_hot_i[1];
  assign data_masked[866] = data_i[866] & sel_one_hot_i[1];
  assign data_masked[865] = data_i[865] & sel_one_hot_i[1];
  assign data_masked[864] = data_i[864] & sel_one_hot_i[1];
  assign data_masked[863] = data_i[863] & sel_one_hot_i[1];
  assign data_masked[862] = data_i[862] & sel_one_hot_i[1];
  assign data_masked[861] = data_i[861] & sel_one_hot_i[1];
  assign data_masked[860] = data_i[860] & sel_one_hot_i[1];
  assign data_masked[859] = data_i[859] & sel_one_hot_i[1];
  assign data_masked[858] = data_i[858] & sel_one_hot_i[1];
  assign data_masked[857] = data_i[857] & sel_one_hot_i[1];
  assign data_masked[856] = data_i[856] & sel_one_hot_i[1];
  assign data_masked[855] = data_i[855] & sel_one_hot_i[1];
  assign data_masked[854] = data_i[854] & sel_one_hot_i[1];
  assign data_masked[853] = data_i[853] & sel_one_hot_i[1];
  assign data_masked[852] = data_i[852] & sel_one_hot_i[1];
  assign data_masked[851] = data_i[851] & sel_one_hot_i[1];
  assign data_masked[850] = data_i[850] & sel_one_hot_i[1];
  assign data_masked[849] = data_i[849] & sel_one_hot_i[1];
  assign data_masked[848] = data_i[848] & sel_one_hot_i[1];
  assign data_masked[847] = data_i[847] & sel_one_hot_i[1];
  assign data_masked[846] = data_i[846] & sel_one_hot_i[1];
  assign data_masked[845] = data_i[845] & sel_one_hot_i[1];
  assign data_masked[844] = data_i[844] & sel_one_hot_i[1];
  assign data_masked[843] = data_i[843] & sel_one_hot_i[1];
  assign data_masked[842] = data_i[842] & sel_one_hot_i[1];
  assign data_masked[841] = data_i[841] & sel_one_hot_i[1];
  assign data_masked[840] = data_i[840] & sel_one_hot_i[1];
  assign data_masked[839] = data_i[839] & sel_one_hot_i[1];
  assign data_masked[838] = data_i[838] & sel_one_hot_i[1];
  assign data_masked[837] = data_i[837] & sel_one_hot_i[1];
  assign data_masked[836] = data_i[836] & sel_one_hot_i[1];
  assign data_masked[835] = data_i[835] & sel_one_hot_i[1];
  assign data_masked[834] = data_i[834] & sel_one_hot_i[1];
  assign data_masked[833] = data_i[833] & sel_one_hot_i[1];
  assign data_masked[832] = data_i[832] & sel_one_hot_i[1];
  assign data_masked[831] = data_i[831] & sel_one_hot_i[1];
  assign data_masked[830] = data_i[830] & sel_one_hot_i[1];
  assign data_masked[829] = data_i[829] & sel_one_hot_i[1];
  assign data_masked[828] = data_i[828] & sel_one_hot_i[1];
  assign data_masked[827] = data_i[827] & sel_one_hot_i[1];
  assign data_masked[826] = data_i[826] & sel_one_hot_i[1];
  assign data_masked[825] = data_i[825] & sel_one_hot_i[1];
  assign data_masked[824] = data_i[824] & sel_one_hot_i[1];
  assign data_masked[823] = data_i[823] & sel_one_hot_i[1];
  assign data_masked[822] = data_i[822] & sel_one_hot_i[1];
  assign data_masked[821] = data_i[821] & sel_one_hot_i[1];
  assign data_masked[820] = data_i[820] & sel_one_hot_i[1];
  assign data_masked[819] = data_i[819] & sel_one_hot_i[1];
  assign data_masked[818] = data_i[818] & sel_one_hot_i[1];
  assign data_masked[817] = data_i[817] & sel_one_hot_i[1];
  assign data_masked[816] = data_i[816] & sel_one_hot_i[1];
  assign data_masked[815] = data_i[815] & sel_one_hot_i[1];
  assign data_masked[814] = data_i[814] & sel_one_hot_i[1];
  assign data_masked[813] = data_i[813] & sel_one_hot_i[1];
  assign data_masked[812] = data_i[812] & sel_one_hot_i[1];
  assign data_masked[811] = data_i[811] & sel_one_hot_i[1];
  assign data_masked[810] = data_i[810] & sel_one_hot_i[1];
  assign data_masked[809] = data_i[809] & sel_one_hot_i[1];
  assign data_masked[808] = data_i[808] & sel_one_hot_i[1];
  assign data_masked[807] = data_i[807] & sel_one_hot_i[1];
  assign data_masked[806] = data_i[806] & sel_one_hot_i[1];
  assign data_masked[805] = data_i[805] & sel_one_hot_i[1];
  assign data_masked[804] = data_i[804] & sel_one_hot_i[1];
  assign data_masked[803] = data_i[803] & sel_one_hot_i[1];
  assign data_masked[802] = data_i[802] & sel_one_hot_i[1];
  assign data_masked[801] = data_i[801] & sel_one_hot_i[1];
  assign data_masked[800] = data_i[800] & sel_one_hot_i[1];
  assign data_masked[799] = data_i[799] & sel_one_hot_i[1];
  assign data_masked[798] = data_i[798] & sel_one_hot_i[1];
  assign data_masked[797] = data_i[797] & sel_one_hot_i[1];
  assign data_masked[796] = data_i[796] & sel_one_hot_i[1];
  assign data_masked[795] = data_i[795] & sel_one_hot_i[1];
  assign data_masked[794] = data_i[794] & sel_one_hot_i[1];
  assign data_masked[793] = data_i[793] & sel_one_hot_i[1];
  assign data_masked[792] = data_i[792] & sel_one_hot_i[1];
  assign data_masked[791] = data_i[791] & sel_one_hot_i[1];
  assign data_masked[790] = data_i[790] & sel_one_hot_i[1];
  assign data_masked[789] = data_i[789] & sel_one_hot_i[1];
  assign data_masked[788] = data_i[788] & sel_one_hot_i[1];
  assign data_masked[787] = data_i[787] & sel_one_hot_i[1];
  assign data_masked[786] = data_i[786] & sel_one_hot_i[1];
  assign data_masked[785] = data_i[785] & sel_one_hot_i[1];
  assign data_masked[784] = data_i[784] & sel_one_hot_i[1];
  assign data_masked[783] = data_i[783] & sel_one_hot_i[1];
  assign data_masked[782] = data_i[782] & sel_one_hot_i[1];
  assign data_masked[781] = data_i[781] & sel_one_hot_i[1];
  assign data_masked[780] = data_i[780] & sel_one_hot_i[1];
  assign data_masked[779] = data_i[779] & sel_one_hot_i[1];
  assign data_masked[778] = data_i[778] & sel_one_hot_i[1];
  assign data_masked[777] = data_i[777] & sel_one_hot_i[1];
  assign data_masked[776] = data_i[776] & sel_one_hot_i[1];
  assign data_masked[775] = data_i[775] & sel_one_hot_i[1];
  assign data_masked[774] = data_i[774] & sel_one_hot_i[1];
  assign data_masked[773] = data_i[773] & sel_one_hot_i[1];
  assign data_masked[772] = data_i[772] & sel_one_hot_i[1];
  assign data_masked[771] = data_i[771] & sel_one_hot_i[1];
  assign data_masked[770] = data_i[770] & sel_one_hot_i[1];
  assign data_masked[769] = data_i[769] & sel_one_hot_i[1];
  assign data_masked[768] = data_i[768] & sel_one_hot_i[1];
  assign data_masked[767] = data_i[767] & sel_one_hot_i[1];
  assign data_masked[766] = data_i[766] & sel_one_hot_i[1];
  assign data_masked[765] = data_i[765] & sel_one_hot_i[1];
  assign data_masked[764] = data_i[764] & sel_one_hot_i[1];
  assign data_masked[763] = data_i[763] & sel_one_hot_i[1];
  assign data_masked[762] = data_i[762] & sel_one_hot_i[1];
  assign data_masked[761] = data_i[761] & sel_one_hot_i[1];
  assign data_masked[760] = data_i[760] & sel_one_hot_i[1];
  assign data_masked[759] = data_i[759] & sel_one_hot_i[1];
  assign data_masked[758] = data_i[758] & sel_one_hot_i[1];
  assign data_masked[757] = data_i[757] & sel_one_hot_i[1];
  assign data_masked[756] = data_i[756] & sel_one_hot_i[1];
  assign data_masked[755] = data_i[755] & sel_one_hot_i[1];
  assign data_masked[754] = data_i[754] & sel_one_hot_i[1];
  assign data_masked[753] = data_i[753] & sel_one_hot_i[1];
  assign data_masked[752] = data_i[752] & sel_one_hot_i[1];
  assign data_masked[751] = data_i[751] & sel_one_hot_i[1];
  assign data_masked[750] = data_i[750] & sel_one_hot_i[1];
  assign data_masked[749] = data_i[749] & sel_one_hot_i[1];
  assign data_masked[748] = data_i[748] & sel_one_hot_i[1];
  assign data_masked[747] = data_i[747] & sel_one_hot_i[1];
  assign data_masked[746] = data_i[746] & sel_one_hot_i[1];
  assign data_masked[745] = data_i[745] & sel_one_hot_i[1];
  assign data_masked[744] = data_i[744] & sel_one_hot_i[1];
  assign data_masked[743] = data_i[743] & sel_one_hot_i[1];
  assign data_masked[742] = data_i[742] & sel_one_hot_i[1];
  assign data_masked[741] = data_i[741] & sel_one_hot_i[1];
  assign data_masked[740] = data_i[740] & sel_one_hot_i[1];
  assign data_masked[739] = data_i[739] & sel_one_hot_i[1];
  assign data_masked[738] = data_i[738] & sel_one_hot_i[1];
  assign data_masked[737] = data_i[737] & sel_one_hot_i[1];
  assign data_masked[736] = data_i[736] & sel_one_hot_i[1];
  assign data_masked[735] = data_i[735] & sel_one_hot_i[1];
  assign data_masked[734] = data_i[734] & sel_one_hot_i[1];
  assign data_masked[733] = data_i[733] & sel_one_hot_i[1];
  assign data_masked[732] = data_i[732] & sel_one_hot_i[1];
  assign data_masked[731] = data_i[731] & sel_one_hot_i[1];
  assign data_masked[730] = data_i[730] & sel_one_hot_i[1];
  assign data_masked[729] = data_i[729] & sel_one_hot_i[1];
  assign data_masked[728] = data_i[728] & sel_one_hot_i[1];
  assign data_masked[727] = data_i[727] & sel_one_hot_i[1];
  assign data_masked[726] = data_i[726] & sel_one_hot_i[1];
  assign data_masked[725] = data_i[725] & sel_one_hot_i[1];
  assign data_masked[724] = data_i[724] & sel_one_hot_i[1];
  assign data_masked[723] = data_i[723] & sel_one_hot_i[1];
  assign data_masked[722] = data_i[722] & sel_one_hot_i[1];
  assign data_masked[721] = data_i[721] & sel_one_hot_i[1];
  assign data_masked[720] = data_i[720] & sel_one_hot_i[1];
  assign data_masked[719] = data_i[719] & sel_one_hot_i[1];
  assign data_masked[718] = data_i[718] & sel_one_hot_i[1];
  assign data_masked[717] = data_i[717] & sel_one_hot_i[1];
  assign data_masked[716] = data_i[716] & sel_one_hot_i[1];
  assign data_masked[715] = data_i[715] & sel_one_hot_i[1];
  assign data_masked[714] = data_i[714] & sel_one_hot_i[1];
  assign data_masked[713] = data_i[713] & sel_one_hot_i[1];
  assign data_masked[712] = data_i[712] & sel_one_hot_i[1];
  assign data_masked[711] = data_i[711] & sel_one_hot_i[1];
  assign data_masked[710] = data_i[710] & sel_one_hot_i[1];
  assign data_masked[709] = data_i[709] & sel_one_hot_i[1];
  assign data_masked[708] = data_i[708] & sel_one_hot_i[1];
  assign data_masked[707] = data_i[707] & sel_one_hot_i[1];
  assign data_masked[706] = data_i[706] & sel_one_hot_i[1];
  assign data_masked[705] = data_i[705] & sel_one_hot_i[1];
  assign data_masked[704] = data_i[704] & sel_one_hot_i[1];
  assign data_masked[703] = data_i[703] & sel_one_hot_i[1];
  assign data_masked[702] = data_i[702] & sel_one_hot_i[1];
  assign data_masked[701] = data_i[701] & sel_one_hot_i[1];
  assign data_masked[700] = data_i[700] & sel_one_hot_i[1];
  assign data_masked[699] = data_i[699] & sel_one_hot_i[1];
  assign data_masked[698] = data_i[698] & sel_one_hot_i[1];
  assign data_masked[697] = data_i[697] & sel_one_hot_i[1];
  assign data_masked[696] = data_i[696] & sel_one_hot_i[1];
  assign data_masked[695] = data_i[695] & sel_one_hot_i[1];
  assign data_masked[694] = data_i[694] & sel_one_hot_i[1];
  assign data_masked[693] = data_i[693] & sel_one_hot_i[1];
  assign data_masked[692] = data_i[692] & sel_one_hot_i[1];
  assign data_masked[691] = data_i[691] & sel_one_hot_i[1];
  assign data_masked[690] = data_i[690] & sel_one_hot_i[1];
  assign data_masked[689] = data_i[689] & sel_one_hot_i[1];
  assign data_masked[688] = data_i[688] & sel_one_hot_i[1];
  assign data_masked[687] = data_i[687] & sel_one_hot_i[1];
  assign data_masked[686] = data_i[686] & sel_one_hot_i[1];
  assign data_masked[685] = data_i[685] & sel_one_hot_i[1];
  assign data_masked[684] = data_i[684] & sel_one_hot_i[1];
  assign data_masked[683] = data_i[683] & sel_one_hot_i[1];
  assign data_masked[682] = data_i[682] & sel_one_hot_i[1];
  assign data_masked[681] = data_i[681] & sel_one_hot_i[1];
  assign data_masked[680] = data_i[680] & sel_one_hot_i[1];
  assign data_masked[679] = data_i[679] & sel_one_hot_i[1];
  assign data_masked[678] = data_i[678] & sel_one_hot_i[1];
  assign data_masked[677] = data_i[677] & sel_one_hot_i[1];
  assign data_masked[676] = data_i[676] & sel_one_hot_i[1];
  assign data_masked[675] = data_i[675] & sel_one_hot_i[1];
  assign data_masked[674] = data_i[674] & sel_one_hot_i[1];
  assign data_masked[673] = data_i[673] & sel_one_hot_i[1];
  assign data_masked[672] = data_i[672] & sel_one_hot_i[1];
  assign data_masked[671] = data_i[671] & sel_one_hot_i[1];
  assign data_masked[670] = data_i[670] & sel_one_hot_i[1];
  assign data_masked[669] = data_i[669] & sel_one_hot_i[1];
  assign data_masked[668] = data_i[668] & sel_one_hot_i[1];
  assign data_masked[667] = data_i[667] & sel_one_hot_i[1];
  assign data_masked[666] = data_i[666] & sel_one_hot_i[1];
  assign data_masked[665] = data_i[665] & sel_one_hot_i[1];
  assign data_masked[664] = data_i[664] & sel_one_hot_i[1];
  assign data_masked[663] = data_i[663] & sel_one_hot_i[1];
  assign data_masked[662] = data_i[662] & sel_one_hot_i[1];
  assign data_masked[661] = data_i[661] & sel_one_hot_i[1];
  assign data_masked[660] = data_i[660] & sel_one_hot_i[1];
  assign data_masked[659] = data_i[659] & sel_one_hot_i[1];
  assign data_masked[658] = data_i[658] & sel_one_hot_i[1];
  assign data_masked[657] = data_i[657] & sel_one_hot_i[1];
  assign data_masked[656] = data_i[656] & sel_one_hot_i[1];
  assign data_masked[655] = data_i[655] & sel_one_hot_i[1];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[1];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[1];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[1];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[1];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[1];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[1];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[1];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[1];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[1];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[1];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[1];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[1];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[1];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[1];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[1];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[1];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[1];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[1];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[1];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[1];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[1];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[1];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[1];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[1];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[1];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[1];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[1];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[1];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[1];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[1];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[1];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[1];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[1];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[1];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[1];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[1];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[1];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[1];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[1];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[1];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[1];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[1];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[1];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[1];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[1];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[1];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[1];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[1];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[1];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[1];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[1];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[1];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[1];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[1];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[1];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[1];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[1];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[1];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[1];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[1];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[1];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[1];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[1];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[1];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[1];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[1];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[1];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[1];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[1];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[1];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[1];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[1];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[1];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[1];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[1];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[1];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[1];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[1];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[1];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[1];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[1];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[1];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[1];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[1];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[1];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[1];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[1];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[1];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[1];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[1];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[1];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[1];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[1];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[1];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[1];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[1];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[1];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[1];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[1];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[1];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[1];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[1];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[1];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[1];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[1];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[1];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[1];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[1];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[1];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[1];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[1];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[1];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[1];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[1];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[1];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[1];
  assign data_masked[1616] = data_i[1616] & sel_one_hot_i[2];
  assign data_masked[1615] = data_i[1615] & sel_one_hot_i[2];
  assign data_masked[1614] = data_i[1614] & sel_one_hot_i[2];
  assign data_masked[1613] = data_i[1613] & sel_one_hot_i[2];
  assign data_masked[1612] = data_i[1612] & sel_one_hot_i[2];
  assign data_masked[1611] = data_i[1611] & sel_one_hot_i[2];
  assign data_masked[1610] = data_i[1610] & sel_one_hot_i[2];
  assign data_masked[1609] = data_i[1609] & sel_one_hot_i[2];
  assign data_masked[1608] = data_i[1608] & sel_one_hot_i[2];
  assign data_masked[1607] = data_i[1607] & sel_one_hot_i[2];
  assign data_masked[1606] = data_i[1606] & sel_one_hot_i[2];
  assign data_masked[1605] = data_i[1605] & sel_one_hot_i[2];
  assign data_masked[1604] = data_i[1604] & sel_one_hot_i[2];
  assign data_masked[1603] = data_i[1603] & sel_one_hot_i[2];
  assign data_masked[1602] = data_i[1602] & sel_one_hot_i[2];
  assign data_masked[1601] = data_i[1601] & sel_one_hot_i[2];
  assign data_masked[1600] = data_i[1600] & sel_one_hot_i[2];
  assign data_masked[1599] = data_i[1599] & sel_one_hot_i[2];
  assign data_masked[1598] = data_i[1598] & sel_one_hot_i[2];
  assign data_masked[1597] = data_i[1597] & sel_one_hot_i[2];
  assign data_masked[1596] = data_i[1596] & sel_one_hot_i[2];
  assign data_masked[1595] = data_i[1595] & sel_one_hot_i[2];
  assign data_masked[1594] = data_i[1594] & sel_one_hot_i[2];
  assign data_masked[1593] = data_i[1593] & sel_one_hot_i[2];
  assign data_masked[1592] = data_i[1592] & sel_one_hot_i[2];
  assign data_masked[1591] = data_i[1591] & sel_one_hot_i[2];
  assign data_masked[1590] = data_i[1590] & sel_one_hot_i[2];
  assign data_masked[1589] = data_i[1589] & sel_one_hot_i[2];
  assign data_masked[1588] = data_i[1588] & sel_one_hot_i[2];
  assign data_masked[1587] = data_i[1587] & sel_one_hot_i[2];
  assign data_masked[1586] = data_i[1586] & sel_one_hot_i[2];
  assign data_masked[1585] = data_i[1585] & sel_one_hot_i[2];
  assign data_masked[1584] = data_i[1584] & sel_one_hot_i[2];
  assign data_masked[1583] = data_i[1583] & sel_one_hot_i[2];
  assign data_masked[1582] = data_i[1582] & sel_one_hot_i[2];
  assign data_masked[1581] = data_i[1581] & sel_one_hot_i[2];
  assign data_masked[1580] = data_i[1580] & sel_one_hot_i[2];
  assign data_masked[1579] = data_i[1579] & sel_one_hot_i[2];
  assign data_masked[1578] = data_i[1578] & sel_one_hot_i[2];
  assign data_masked[1577] = data_i[1577] & sel_one_hot_i[2];
  assign data_masked[1576] = data_i[1576] & sel_one_hot_i[2];
  assign data_masked[1575] = data_i[1575] & sel_one_hot_i[2];
  assign data_masked[1574] = data_i[1574] & sel_one_hot_i[2];
  assign data_masked[1573] = data_i[1573] & sel_one_hot_i[2];
  assign data_masked[1572] = data_i[1572] & sel_one_hot_i[2];
  assign data_masked[1571] = data_i[1571] & sel_one_hot_i[2];
  assign data_masked[1570] = data_i[1570] & sel_one_hot_i[2];
  assign data_masked[1569] = data_i[1569] & sel_one_hot_i[2];
  assign data_masked[1568] = data_i[1568] & sel_one_hot_i[2];
  assign data_masked[1567] = data_i[1567] & sel_one_hot_i[2];
  assign data_masked[1566] = data_i[1566] & sel_one_hot_i[2];
  assign data_masked[1565] = data_i[1565] & sel_one_hot_i[2];
  assign data_masked[1564] = data_i[1564] & sel_one_hot_i[2];
  assign data_masked[1563] = data_i[1563] & sel_one_hot_i[2];
  assign data_masked[1562] = data_i[1562] & sel_one_hot_i[2];
  assign data_masked[1561] = data_i[1561] & sel_one_hot_i[2];
  assign data_masked[1560] = data_i[1560] & sel_one_hot_i[2];
  assign data_masked[1559] = data_i[1559] & sel_one_hot_i[2];
  assign data_masked[1558] = data_i[1558] & sel_one_hot_i[2];
  assign data_masked[1557] = data_i[1557] & sel_one_hot_i[2];
  assign data_masked[1556] = data_i[1556] & sel_one_hot_i[2];
  assign data_masked[1555] = data_i[1555] & sel_one_hot_i[2];
  assign data_masked[1554] = data_i[1554] & sel_one_hot_i[2];
  assign data_masked[1553] = data_i[1553] & sel_one_hot_i[2];
  assign data_masked[1552] = data_i[1552] & sel_one_hot_i[2];
  assign data_masked[1551] = data_i[1551] & sel_one_hot_i[2];
  assign data_masked[1550] = data_i[1550] & sel_one_hot_i[2];
  assign data_masked[1549] = data_i[1549] & sel_one_hot_i[2];
  assign data_masked[1548] = data_i[1548] & sel_one_hot_i[2];
  assign data_masked[1547] = data_i[1547] & sel_one_hot_i[2];
  assign data_masked[1546] = data_i[1546] & sel_one_hot_i[2];
  assign data_masked[1545] = data_i[1545] & sel_one_hot_i[2];
  assign data_masked[1544] = data_i[1544] & sel_one_hot_i[2];
  assign data_masked[1543] = data_i[1543] & sel_one_hot_i[2];
  assign data_masked[1542] = data_i[1542] & sel_one_hot_i[2];
  assign data_masked[1541] = data_i[1541] & sel_one_hot_i[2];
  assign data_masked[1540] = data_i[1540] & sel_one_hot_i[2];
  assign data_masked[1539] = data_i[1539] & sel_one_hot_i[2];
  assign data_masked[1538] = data_i[1538] & sel_one_hot_i[2];
  assign data_masked[1537] = data_i[1537] & sel_one_hot_i[2];
  assign data_masked[1536] = data_i[1536] & sel_one_hot_i[2];
  assign data_masked[1535] = data_i[1535] & sel_one_hot_i[2];
  assign data_masked[1534] = data_i[1534] & sel_one_hot_i[2];
  assign data_masked[1533] = data_i[1533] & sel_one_hot_i[2];
  assign data_masked[1532] = data_i[1532] & sel_one_hot_i[2];
  assign data_masked[1531] = data_i[1531] & sel_one_hot_i[2];
  assign data_masked[1530] = data_i[1530] & sel_one_hot_i[2];
  assign data_masked[1529] = data_i[1529] & sel_one_hot_i[2];
  assign data_masked[1528] = data_i[1528] & sel_one_hot_i[2];
  assign data_masked[1527] = data_i[1527] & sel_one_hot_i[2];
  assign data_masked[1526] = data_i[1526] & sel_one_hot_i[2];
  assign data_masked[1525] = data_i[1525] & sel_one_hot_i[2];
  assign data_masked[1524] = data_i[1524] & sel_one_hot_i[2];
  assign data_masked[1523] = data_i[1523] & sel_one_hot_i[2];
  assign data_masked[1522] = data_i[1522] & sel_one_hot_i[2];
  assign data_masked[1521] = data_i[1521] & sel_one_hot_i[2];
  assign data_masked[1520] = data_i[1520] & sel_one_hot_i[2];
  assign data_masked[1519] = data_i[1519] & sel_one_hot_i[2];
  assign data_masked[1518] = data_i[1518] & sel_one_hot_i[2];
  assign data_masked[1517] = data_i[1517] & sel_one_hot_i[2];
  assign data_masked[1516] = data_i[1516] & sel_one_hot_i[2];
  assign data_masked[1515] = data_i[1515] & sel_one_hot_i[2];
  assign data_masked[1514] = data_i[1514] & sel_one_hot_i[2];
  assign data_masked[1513] = data_i[1513] & sel_one_hot_i[2];
  assign data_masked[1512] = data_i[1512] & sel_one_hot_i[2];
  assign data_masked[1511] = data_i[1511] & sel_one_hot_i[2];
  assign data_masked[1510] = data_i[1510] & sel_one_hot_i[2];
  assign data_masked[1509] = data_i[1509] & sel_one_hot_i[2];
  assign data_masked[1508] = data_i[1508] & sel_one_hot_i[2];
  assign data_masked[1507] = data_i[1507] & sel_one_hot_i[2];
  assign data_masked[1506] = data_i[1506] & sel_one_hot_i[2];
  assign data_masked[1505] = data_i[1505] & sel_one_hot_i[2];
  assign data_masked[1504] = data_i[1504] & sel_one_hot_i[2];
  assign data_masked[1503] = data_i[1503] & sel_one_hot_i[2];
  assign data_masked[1502] = data_i[1502] & sel_one_hot_i[2];
  assign data_masked[1501] = data_i[1501] & sel_one_hot_i[2];
  assign data_masked[1500] = data_i[1500] & sel_one_hot_i[2];
  assign data_masked[1499] = data_i[1499] & sel_one_hot_i[2];
  assign data_masked[1498] = data_i[1498] & sel_one_hot_i[2];
  assign data_masked[1497] = data_i[1497] & sel_one_hot_i[2];
  assign data_masked[1496] = data_i[1496] & sel_one_hot_i[2];
  assign data_masked[1495] = data_i[1495] & sel_one_hot_i[2];
  assign data_masked[1494] = data_i[1494] & sel_one_hot_i[2];
  assign data_masked[1493] = data_i[1493] & sel_one_hot_i[2];
  assign data_masked[1492] = data_i[1492] & sel_one_hot_i[2];
  assign data_masked[1491] = data_i[1491] & sel_one_hot_i[2];
  assign data_masked[1490] = data_i[1490] & sel_one_hot_i[2];
  assign data_masked[1489] = data_i[1489] & sel_one_hot_i[2];
  assign data_masked[1488] = data_i[1488] & sel_one_hot_i[2];
  assign data_masked[1487] = data_i[1487] & sel_one_hot_i[2];
  assign data_masked[1486] = data_i[1486] & sel_one_hot_i[2];
  assign data_masked[1485] = data_i[1485] & sel_one_hot_i[2];
  assign data_masked[1484] = data_i[1484] & sel_one_hot_i[2];
  assign data_masked[1483] = data_i[1483] & sel_one_hot_i[2];
  assign data_masked[1482] = data_i[1482] & sel_one_hot_i[2];
  assign data_masked[1481] = data_i[1481] & sel_one_hot_i[2];
  assign data_masked[1480] = data_i[1480] & sel_one_hot_i[2];
  assign data_masked[1479] = data_i[1479] & sel_one_hot_i[2];
  assign data_masked[1478] = data_i[1478] & sel_one_hot_i[2];
  assign data_masked[1477] = data_i[1477] & sel_one_hot_i[2];
  assign data_masked[1476] = data_i[1476] & sel_one_hot_i[2];
  assign data_masked[1475] = data_i[1475] & sel_one_hot_i[2];
  assign data_masked[1474] = data_i[1474] & sel_one_hot_i[2];
  assign data_masked[1473] = data_i[1473] & sel_one_hot_i[2];
  assign data_masked[1472] = data_i[1472] & sel_one_hot_i[2];
  assign data_masked[1471] = data_i[1471] & sel_one_hot_i[2];
  assign data_masked[1470] = data_i[1470] & sel_one_hot_i[2];
  assign data_masked[1469] = data_i[1469] & sel_one_hot_i[2];
  assign data_masked[1468] = data_i[1468] & sel_one_hot_i[2];
  assign data_masked[1467] = data_i[1467] & sel_one_hot_i[2];
  assign data_masked[1466] = data_i[1466] & sel_one_hot_i[2];
  assign data_masked[1465] = data_i[1465] & sel_one_hot_i[2];
  assign data_masked[1464] = data_i[1464] & sel_one_hot_i[2];
  assign data_masked[1463] = data_i[1463] & sel_one_hot_i[2];
  assign data_masked[1462] = data_i[1462] & sel_one_hot_i[2];
  assign data_masked[1461] = data_i[1461] & sel_one_hot_i[2];
  assign data_masked[1460] = data_i[1460] & sel_one_hot_i[2];
  assign data_masked[1459] = data_i[1459] & sel_one_hot_i[2];
  assign data_masked[1458] = data_i[1458] & sel_one_hot_i[2];
  assign data_masked[1457] = data_i[1457] & sel_one_hot_i[2];
  assign data_masked[1456] = data_i[1456] & sel_one_hot_i[2];
  assign data_masked[1455] = data_i[1455] & sel_one_hot_i[2];
  assign data_masked[1454] = data_i[1454] & sel_one_hot_i[2];
  assign data_masked[1453] = data_i[1453] & sel_one_hot_i[2];
  assign data_masked[1452] = data_i[1452] & sel_one_hot_i[2];
  assign data_masked[1451] = data_i[1451] & sel_one_hot_i[2];
  assign data_masked[1450] = data_i[1450] & sel_one_hot_i[2];
  assign data_masked[1449] = data_i[1449] & sel_one_hot_i[2];
  assign data_masked[1448] = data_i[1448] & sel_one_hot_i[2];
  assign data_masked[1447] = data_i[1447] & sel_one_hot_i[2];
  assign data_masked[1446] = data_i[1446] & sel_one_hot_i[2];
  assign data_masked[1445] = data_i[1445] & sel_one_hot_i[2];
  assign data_masked[1444] = data_i[1444] & sel_one_hot_i[2];
  assign data_masked[1443] = data_i[1443] & sel_one_hot_i[2];
  assign data_masked[1442] = data_i[1442] & sel_one_hot_i[2];
  assign data_masked[1441] = data_i[1441] & sel_one_hot_i[2];
  assign data_masked[1440] = data_i[1440] & sel_one_hot_i[2];
  assign data_masked[1439] = data_i[1439] & sel_one_hot_i[2];
  assign data_masked[1438] = data_i[1438] & sel_one_hot_i[2];
  assign data_masked[1437] = data_i[1437] & sel_one_hot_i[2];
  assign data_masked[1436] = data_i[1436] & sel_one_hot_i[2];
  assign data_masked[1435] = data_i[1435] & sel_one_hot_i[2];
  assign data_masked[1434] = data_i[1434] & sel_one_hot_i[2];
  assign data_masked[1433] = data_i[1433] & sel_one_hot_i[2];
  assign data_masked[1432] = data_i[1432] & sel_one_hot_i[2];
  assign data_masked[1431] = data_i[1431] & sel_one_hot_i[2];
  assign data_masked[1430] = data_i[1430] & sel_one_hot_i[2];
  assign data_masked[1429] = data_i[1429] & sel_one_hot_i[2];
  assign data_masked[1428] = data_i[1428] & sel_one_hot_i[2];
  assign data_masked[1427] = data_i[1427] & sel_one_hot_i[2];
  assign data_masked[1426] = data_i[1426] & sel_one_hot_i[2];
  assign data_masked[1425] = data_i[1425] & sel_one_hot_i[2];
  assign data_masked[1424] = data_i[1424] & sel_one_hot_i[2];
  assign data_masked[1423] = data_i[1423] & sel_one_hot_i[2];
  assign data_masked[1422] = data_i[1422] & sel_one_hot_i[2];
  assign data_masked[1421] = data_i[1421] & sel_one_hot_i[2];
  assign data_masked[1420] = data_i[1420] & sel_one_hot_i[2];
  assign data_masked[1419] = data_i[1419] & sel_one_hot_i[2];
  assign data_masked[1418] = data_i[1418] & sel_one_hot_i[2];
  assign data_masked[1417] = data_i[1417] & sel_one_hot_i[2];
  assign data_masked[1416] = data_i[1416] & sel_one_hot_i[2];
  assign data_masked[1415] = data_i[1415] & sel_one_hot_i[2];
  assign data_masked[1414] = data_i[1414] & sel_one_hot_i[2];
  assign data_masked[1413] = data_i[1413] & sel_one_hot_i[2];
  assign data_masked[1412] = data_i[1412] & sel_one_hot_i[2];
  assign data_masked[1411] = data_i[1411] & sel_one_hot_i[2];
  assign data_masked[1410] = data_i[1410] & sel_one_hot_i[2];
  assign data_masked[1409] = data_i[1409] & sel_one_hot_i[2];
  assign data_masked[1408] = data_i[1408] & sel_one_hot_i[2];
  assign data_masked[1407] = data_i[1407] & sel_one_hot_i[2];
  assign data_masked[1406] = data_i[1406] & sel_one_hot_i[2];
  assign data_masked[1405] = data_i[1405] & sel_one_hot_i[2];
  assign data_masked[1404] = data_i[1404] & sel_one_hot_i[2];
  assign data_masked[1403] = data_i[1403] & sel_one_hot_i[2];
  assign data_masked[1402] = data_i[1402] & sel_one_hot_i[2];
  assign data_masked[1401] = data_i[1401] & sel_one_hot_i[2];
  assign data_masked[1400] = data_i[1400] & sel_one_hot_i[2];
  assign data_masked[1399] = data_i[1399] & sel_one_hot_i[2];
  assign data_masked[1398] = data_i[1398] & sel_one_hot_i[2];
  assign data_masked[1397] = data_i[1397] & sel_one_hot_i[2];
  assign data_masked[1396] = data_i[1396] & sel_one_hot_i[2];
  assign data_masked[1395] = data_i[1395] & sel_one_hot_i[2];
  assign data_masked[1394] = data_i[1394] & sel_one_hot_i[2];
  assign data_masked[1393] = data_i[1393] & sel_one_hot_i[2];
  assign data_masked[1392] = data_i[1392] & sel_one_hot_i[2];
  assign data_masked[1391] = data_i[1391] & sel_one_hot_i[2];
  assign data_masked[1390] = data_i[1390] & sel_one_hot_i[2];
  assign data_masked[1389] = data_i[1389] & sel_one_hot_i[2];
  assign data_masked[1388] = data_i[1388] & sel_one_hot_i[2];
  assign data_masked[1387] = data_i[1387] & sel_one_hot_i[2];
  assign data_masked[1386] = data_i[1386] & sel_one_hot_i[2];
  assign data_masked[1385] = data_i[1385] & sel_one_hot_i[2];
  assign data_masked[1384] = data_i[1384] & sel_one_hot_i[2];
  assign data_masked[1383] = data_i[1383] & sel_one_hot_i[2];
  assign data_masked[1382] = data_i[1382] & sel_one_hot_i[2];
  assign data_masked[1381] = data_i[1381] & sel_one_hot_i[2];
  assign data_masked[1380] = data_i[1380] & sel_one_hot_i[2];
  assign data_masked[1379] = data_i[1379] & sel_one_hot_i[2];
  assign data_masked[1378] = data_i[1378] & sel_one_hot_i[2];
  assign data_masked[1377] = data_i[1377] & sel_one_hot_i[2];
  assign data_masked[1376] = data_i[1376] & sel_one_hot_i[2];
  assign data_masked[1375] = data_i[1375] & sel_one_hot_i[2];
  assign data_masked[1374] = data_i[1374] & sel_one_hot_i[2];
  assign data_masked[1373] = data_i[1373] & sel_one_hot_i[2];
  assign data_masked[1372] = data_i[1372] & sel_one_hot_i[2];
  assign data_masked[1371] = data_i[1371] & sel_one_hot_i[2];
  assign data_masked[1370] = data_i[1370] & sel_one_hot_i[2];
  assign data_masked[1369] = data_i[1369] & sel_one_hot_i[2];
  assign data_masked[1368] = data_i[1368] & sel_one_hot_i[2];
  assign data_masked[1367] = data_i[1367] & sel_one_hot_i[2];
  assign data_masked[1366] = data_i[1366] & sel_one_hot_i[2];
  assign data_masked[1365] = data_i[1365] & sel_one_hot_i[2];
  assign data_masked[1364] = data_i[1364] & sel_one_hot_i[2];
  assign data_masked[1363] = data_i[1363] & sel_one_hot_i[2];
  assign data_masked[1362] = data_i[1362] & sel_one_hot_i[2];
  assign data_masked[1361] = data_i[1361] & sel_one_hot_i[2];
  assign data_masked[1360] = data_i[1360] & sel_one_hot_i[2];
  assign data_masked[1359] = data_i[1359] & sel_one_hot_i[2];
  assign data_masked[1358] = data_i[1358] & sel_one_hot_i[2];
  assign data_masked[1357] = data_i[1357] & sel_one_hot_i[2];
  assign data_masked[1356] = data_i[1356] & sel_one_hot_i[2];
  assign data_masked[1355] = data_i[1355] & sel_one_hot_i[2];
  assign data_masked[1354] = data_i[1354] & sel_one_hot_i[2];
  assign data_masked[1353] = data_i[1353] & sel_one_hot_i[2];
  assign data_masked[1352] = data_i[1352] & sel_one_hot_i[2];
  assign data_masked[1351] = data_i[1351] & sel_one_hot_i[2];
  assign data_masked[1350] = data_i[1350] & sel_one_hot_i[2];
  assign data_masked[1349] = data_i[1349] & sel_one_hot_i[2];
  assign data_masked[1348] = data_i[1348] & sel_one_hot_i[2];
  assign data_masked[1347] = data_i[1347] & sel_one_hot_i[2];
  assign data_masked[1346] = data_i[1346] & sel_one_hot_i[2];
  assign data_masked[1345] = data_i[1345] & sel_one_hot_i[2];
  assign data_masked[1344] = data_i[1344] & sel_one_hot_i[2];
  assign data_masked[1343] = data_i[1343] & sel_one_hot_i[2];
  assign data_masked[1342] = data_i[1342] & sel_one_hot_i[2];
  assign data_masked[1341] = data_i[1341] & sel_one_hot_i[2];
  assign data_masked[1340] = data_i[1340] & sel_one_hot_i[2];
  assign data_masked[1339] = data_i[1339] & sel_one_hot_i[2];
  assign data_masked[1338] = data_i[1338] & sel_one_hot_i[2];
  assign data_masked[1337] = data_i[1337] & sel_one_hot_i[2];
  assign data_masked[1336] = data_i[1336] & sel_one_hot_i[2];
  assign data_masked[1335] = data_i[1335] & sel_one_hot_i[2];
  assign data_masked[1334] = data_i[1334] & sel_one_hot_i[2];
  assign data_masked[1333] = data_i[1333] & sel_one_hot_i[2];
  assign data_masked[1332] = data_i[1332] & sel_one_hot_i[2];
  assign data_masked[1331] = data_i[1331] & sel_one_hot_i[2];
  assign data_masked[1330] = data_i[1330] & sel_one_hot_i[2];
  assign data_masked[1329] = data_i[1329] & sel_one_hot_i[2];
  assign data_masked[1328] = data_i[1328] & sel_one_hot_i[2];
  assign data_masked[1327] = data_i[1327] & sel_one_hot_i[2];
  assign data_masked[1326] = data_i[1326] & sel_one_hot_i[2];
  assign data_masked[1325] = data_i[1325] & sel_one_hot_i[2];
  assign data_masked[1324] = data_i[1324] & sel_one_hot_i[2];
  assign data_masked[1323] = data_i[1323] & sel_one_hot_i[2];
  assign data_masked[1322] = data_i[1322] & sel_one_hot_i[2];
  assign data_masked[1321] = data_i[1321] & sel_one_hot_i[2];
  assign data_masked[1320] = data_i[1320] & sel_one_hot_i[2];
  assign data_masked[1319] = data_i[1319] & sel_one_hot_i[2];
  assign data_masked[1318] = data_i[1318] & sel_one_hot_i[2];
  assign data_masked[1317] = data_i[1317] & sel_one_hot_i[2];
  assign data_masked[1316] = data_i[1316] & sel_one_hot_i[2];
  assign data_masked[1315] = data_i[1315] & sel_one_hot_i[2];
  assign data_masked[1314] = data_i[1314] & sel_one_hot_i[2];
  assign data_masked[1313] = data_i[1313] & sel_one_hot_i[2];
  assign data_masked[1312] = data_i[1312] & sel_one_hot_i[2];
  assign data_masked[1311] = data_i[1311] & sel_one_hot_i[2];
  assign data_masked[1310] = data_i[1310] & sel_one_hot_i[2];
  assign data_masked[1309] = data_i[1309] & sel_one_hot_i[2];
  assign data_masked[1308] = data_i[1308] & sel_one_hot_i[2];
  assign data_masked[1307] = data_i[1307] & sel_one_hot_i[2];
  assign data_masked[1306] = data_i[1306] & sel_one_hot_i[2];
  assign data_masked[1305] = data_i[1305] & sel_one_hot_i[2];
  assign data_masked[1304] = data_i[1304] & sel_one_hot_i[2];
  assign data_masked[1303] = data_i[1303] & sel_one_hot_i[2];
  assign data_masked[1302] = data_i[1302] & sel_one_hot_i[2];
  assign data_masked[1301] = data_i[1301] & sel_one_hot_i[2];
  assign data_masked[1300] = data_i[1300] & sel_one_hot_i[2];
  assign data_masked[1299] = data_i[1299] & sel_one_hot_i[2];
  assign data_masked[1298] = data_i[1298] & sel_one_hot_i[2];
  assign data_masked[1297] = data_i[1297] & sel_one_hot_i[2];
  assign data_masked[1296] = data_i[1296] & sel_one_hot_i[2];
  assign data_masked[1295] = data_i[1295] & sel_one_hot_i[2];
  assign data_masked[1294] = data_i[1294] & sel_one_hot_i[2];
  assign data_masked[1293] = data_i[1293] & sel_one_hot_i[2];
  assign data_masked[1292] = data_i[1292] & sel_one_hot_i[2];
  assign data_masked[1291] = data_i[1291] & sel_one_hot_i[2];
  assign data_masked[1290] = data_i[1290] & sel_one_hot_i[2];
  assign data_masked[1289] = data_i[1289] & sel_one_hot_i[2];
  assign data_masked[1288] = data_i[1288] & sel_one_hot_i[2];
  assign data_masked[1287] = data_i[1287] & sel_one_hot_i[2];
  assign data_masked[1286] = data_i[1286] & sel_one_hot_i[2];
  assign data_masked[1285] = data_i[1285] & sel_one_hot_i[2];
  assign data_masked[1284] = data_i[1284] & sel_one_hot_i[2];
  assign data_masked[1283] = data_i[1283] & sel_one_hot_i[2];
  assign data_masked[1282] = data_i[1282] & sel_one_hot_i[2];
  assign data_masked[1281] = data_i[1281] & sel_one_hot_i[2];
  assign data_masked[1280] = data_i[1280] & sel_one_hot_i[2];
  assign data_masked[1279] = data_i[1279] & sel_one_hot_i[2];
  assign data_masked[1278] = data_i[1278] & sel_one_hot_i[2];
  assign data_masked[1277] = data_i[1277] & sel_one_hot_i[2];
  assign data_masked[1276] = data_i[1276] & sel_one_hot_i[2];
  assign data_masked[1275] = data_i[1275] & sel_one_hot_i[2];
  assign data_masked[1274] = data_i[1274] & sel_one_hot_i[2];
  assign data_masked[1273] = data_i[1273] & sel_one_hot_i[2];
  assign data_masked[1272] = data_i[1272] & sel_one_hot_i[2];
  assign data_masked[1271] = data_i[1271] & sel_one_hot_i[2];
  assign data_masked[1270] = data_i[1270] & sel_one_hot_i[2];
  assign data_masked[1269] = data_i[1269] & sel_one_hot_i[2];
  assign data_masked[1268] = data_i[1268] & sel_one_hot_i[2];
  assign data_masked[1267] = data_i[1267] & sel_one_hot_i[2];
  assign data_masked[1266] = data_i[1266] & sel_one_hot_i[2];
  assign data_masked[1265] = data_i[1265] & sel_one_hot_i[2];
  assign data_masked[1264] = data_i[1264] & sel_one_hot_i[2];
  assign data_masked[1263] = data_i[1263] & sel_one_hot_i[2];
  assign data_masked[1262] = data_i[1262] & sel_one_hot_i[2];
  assign data_masked[1261] = data_i[1261] & sel_one_hot_i[2];
  assign data_masked[1260] = data_i[1260] & sel_one_hot_i[2];
  assign data_masked[1259] = data_i[1259] & sel_one_hot_i[2];
  assign data_masked[1258] = data_i[1258] & sel_one_hot_i[2];
  assign data_masked[1257] = data_i[1257] & sel_one_hot_i[2];
  assign data_masked[1256] = data_i[1256] & sel_one_hot_i[2];
  assign data_masked[1255] = data_i[1255] & sel_one_hot_i[2];
  assign data_masked[1254] = data_i[1254] & sel_one_hot_i[2];
  assign data_masked[1253] = data_i[1253] & sel_one_hot_i[2];
  assign data_masked[1252] = data_i[1252] & sel_one_hot_i[2];
  assign data_masked[1251] = data_i[1251] & sel_one_hot_i[2];
  assign data_masked[1250] = data_i[1250] & sel_one_hot_i[2];
  assign data_masked[1249] = data_i[1249] & sel_one_hot_i[2];
  assign data_masked[1248] = data_i[1248] & sel_one_hot_i[2];
  assign data_masked[1247] = data_i[1247] & sel_one_hot_i[2];
  assign data_masked[1246] = data_i[1246] & sel_one_hot_i[2];
  assign data_masked[1245] = data_i[1245] & sel_one_hot_i[2];
  assign data_masked[1244] = data_i[1244] & sel_one_hot_i[2];
  assign data_masked[1243] = data_i[1243] & sel_one_hot_i[2];
  assign data_masked[1242] = data_i[1242] & sel_one_hot_i[2];
  assign data_masked[1241] = data_i[1241] & sel_one_hot_i[2];
  assign data_masked[1240] = data_i[1240] & sel_one_hot_i[2];
  assign data_masked[1239] = data_i[1239] & sel_one_hot_i[2];
  assign data_masked[1238] = data_i[1238] & sel_one_hot_i[2];
  assign data_masked[1237] = data_i[1237] & sel_one_hot_i[2];
  assign data_masked[1236] = data_i[1236] & sel_one_hot_i[2];
  assign data_masked[1235] = data_i[1235] & sel_one_hot_i[2];
  assign data_masked[1234] = data_i[1234] & sel_one_hot_i[2];
  assign data_masked[1233] = data_i[1233] & sel_one_hot_i[2];
  assign data_masked[1232] = data_i[1232] & sel_one_hot_i[2];
  assign data_masked[1231] = data_i[1231] & sel_one_hot_i[2];
  assign data_masked[1230] = data_i[1230] & sel_one_hot_i[2];
  assign data_masked[1229] = data_i[1229] & sel_one_hot_i[2];
  assign data_masked[1228] = data_i[1228] & sel_one_hot_i[2];
  assign data_masked[1227] = data_i[1227] & sel_one_hot_i[2];
  assign data_masked[1226] = data_i[1226] & sel_one_hot_i[2];
  assign data_masked[1225] = data_i[1225] & sel_one_hot_i[2];
  assign data_masked[1224] = data_i[1224] & sel_one_hot_i[2];
  assign data_masked[1223] = data_i[1223] & sel_one_hot_i[2];
  assign data_masked[1222] = data_i[1222] & sel_one_hot_i[2];
  assign data_masked[1221] = data_i[1221] & sel_one_hot_i[2];
  assign data_masked[1220] = data_i[1220] & sel_one_hot_i[2];
  assign data_masked[1219] = data_i[1219] & sel_one_hot_i[2];
  assign data_masked[1218] = data_i[1218] & sel_one_hot_i[2];
  assign data_masked[1217] = data_i[1217] & sel_one_hot_i[2];
  assign data_masked[1216] = data_i[1216] & sel_one_hot_i[2];
  assign data_masked[1215] = data_i[1215] & sel_one_hot_i[2];
  assign data_masked[1214] = data_i[1214] & sel_one_hot_i[2];
  assign data_masked[1213] = data_i[1213] & sel_one_hot_i[2];
  assign data_masked[1212] = data_i[1212] & sel_one_hot_i[2];
  assign data_masked[1211] = data_i[1211] & sel_one_hot_i[2];
  assign data_masked[1210] = data_i[1210] & sel_one_hot_i[2];
  assign data_masked[1209] = data_i[1209] & sel_one_hot_i[2];
  assign data_masked[1208] = data_i[1208] & sel_one_hot_i[2];
  assign data_masked[1207] = data_i[1207] & sel_one_hot_i[2];
  assign data_masked[1206] = data_i[1206] & sel_one_hot_i[2];
  assign data_masked[1205] = data_i[1205] & sel_one_hot_i[2];
  assign data_masked[1204] = data_i[1204] & sel_one_hot_i[2];
  assign data_masked[1203] = data_i[1203] & sel_one_hot_i[2];
  assign data_masked[1202] = data_i[1202] & sel_one_hot_i[2];
  assign data_masked[1201] = data_i[1201] & sel_one_hot_i[2];
  assign data_masked[1200] = data_i[1200] & sel_one_hot_i[2];
  assign data_masked[1199] = data_i[1199] & sel_one_hot_i[2];
  assign data_masked[1198] = data_i[1198] & sel_one_hot_i[2];
  assign data_masked[1197] = data_i[1197] & sel_one_hot_i[2];
  assign data_masked[1196] = data_i[1196] & sel_one_hot_i[2];
  assign data_masked[1195] = data_i[1195] & sel_one_hot_i[2];
  assign data_masked[1194] = data_i[1194] & sel_one_hot_i[2];
  assign data_masked[1193] = data_i[1193] & sel_one_hot_i[2];
  assign data_masked[1192] = data_i[1192] & sel_one_hot_i[2];
  assign data_masked[1191] = data_i[1191] & sel_one_hot_i[2];
  assign data_masked[1190] = data_i[1190] & sel_one_hot_i[2];
  assign data_masked[1189] = data_i[1189] & sel_one_hot_i[2];
  assign data_masked[1188] = data_i[1188] & sel_one_hot_i[2];
  assign data_masked[1187] = data_i[1187] & sel_one_hot_i[2];
  assign data_masked[1186] = data_i[1186] & sel_one_hot_i[2];
  assign data_masked[1185] = data_i[1185] & sel_one_hot_i[2];
  assign data_masked[1184] = data_i[1184] & sel_one_hot_i[2];
  assign data_masked[1183] = data_i[1183] & sel_one_hot_i[2];
  assign data_masked[1182] = data_i[1182] & sel_one_hot_i[2];
  assign data_masked[1181] = data_i[1181] & sel_one_hot_i[2];
  assign data_masked[1180] = data_i[1180] & sel_one_hot_i[2];
  assign data_masked[1179] = data_i[1179] & sel_one_hot_i[2];
  assign data_masked[1178] = data_i[1178] & sel_one_hot_i[2];
  assign data_masked[1177] = data_i[1177] & sel_one_hot_i[2];
  assign data_masked[1176] = data_i[1176] & sel_one_hot_i[2];
  assign data_masked[1175] = data_i[1175] & sel_one_hot_i[2];
  assign data_masked[1174] = data_i[1174] & sel_one_hot_i[2];
  assign data_masked[1173] = data_i[1173] & sel_one_hot_i[2];
  assign data_masked[1172] = data_i[1172] & sel_one_hot_i[2];
  assign data_masked[1171] = data_i[1171] & sel_one_hot_i[2];
  assign data_masked[1170] = data_i[1170] & sel_one_hot_i[2];
  assign data_masked[1169] = data_i[1169] & sel_one_hot_i[2];
  assign data_masked[1168] = data_i[1168] & sel_one_hot_i[2];
  assign data_masked[1167] = data_i[1167] & sel_one_hot_i[2];
  assign data_masked[1166] = data_i[1166] & sel_one_hot_i[2];
  assign data_masked[1165] = data_i[1165] & sel_one_hot_i[2];
  assign data_masked[1164] = data_i[1164] & sel_one_hot_i[2];
  assign data_masked[1163] = data_i[1163] & sel_one_hot_i[2];
  assign data_masked[1162] = data_i[1162] & sel_one_hot_i[2];
  assign data_masked[1161] = data_i[1161] & sel_one_hot_i[2];
  assign data_masked[1160] = data_i[1160] & sel_one_hot_i[2];
  assign data_masked[1159] = data_i[1159] & sel_one_hot_i[2];
  assign data_masked[1158] = data_i[1158] & sel_one_hot_i[2];
  assign data_masked[1157] = data_i[1157] & sel_one_hot_i[2];
  assign data_masked[1156] = data_i[1156] & sel_one_hot_i[2];
  assign data_masked[1155] = data_i[1155] & sel_one_hot_i[2];
  assign data_masked[1154] = data_i[1154] & sel_one_hot_i[2];
  assign data_masked[1153] = data_i[1153] & sel_one_hot_i[2];
  assign data_masked[1152] = data_i[1152] & sel_one_hot_i[2];
  assign data_masked[1151] = data_i[1151] & sel_one_hot_i[2];
  assign data_masked[1150] = data_i[1150] & sel_one_hot_i[2];
  assign data_masked[1149] = data_i[1149] & sel_one_hot_i[2];
  assign data_masked[1148] = data_i[1148] & sel_one_hot_i[2];
  assign data_masked[1147] = data_i[1147] & sel_one_hot_i[2];
  assign data_masked[1146] = data_i[1146] & sel_one_hot_i[2];
  assign data_masked[1145] = data_i[1145] & sel_one_hot_i[2];
  assign data_masked[1144] = data_i[1144] & sel_one_hot_i[2];
  assign data_masked[1143] = data_i[1143] & sel_one_hot_i[2];
  assign data_masked[1142] = data_i[1142] & sel_one_hot_i[2];
  assign data_masked[1141] = data_i[1141] & sel_one_hot_i[2];
  assign data_masked[1140] = data_i[1140] & sel_one_hot_i[2];
  assign data_masked[1139] = data_i[1139] & sel_one_hot_i[2];
  assign data_masked[1138] = data_i[1138] & sel_one_hot_i[2];
  assign data_masked[1137] = data_i[1137] & sel_one_hot_i[2];
  assign data_masked[1136] = data_i[1136] & sel_one_hot_i[2];
  assign data_masked[1135] = data_i[1135] & sel_one_hot_i[2];
  assign data_masked[1134] = data_i[1134] & sel_one_hot_i[2];
  assign data_masked[1133] = data_i[1133] & sel_one_hot_i[2];
  assign data_masked[1132] = data_i[1132] & sel_one_hot_i[2];
  assign data_masked[1131] = data_i[1131] & sel_one_hot_i[2];
  assign data_masked[1130] = data_i[1130] & sel_one_hot_i[2];
  assign data_masked[1129] = data_i[1129] & sel_one_hot_i[2];
  assign data_masked[1128] = data_i[1128] & sel_one_hot_i[2];
  assign data_masked[1127] = data_i[1127] & sel_one_hot_i[2];
  assign data_masked[1126] = data_i[1126] & sel_one_hot_i[2];
  assign data_masked[1125] = data_i[1125] & sel_one_hot_i[2];
  assign data_masked[1124] = data_i[1124] & sel_one_hot_i[2];
  assign data_masked[1123] = data_i[1123] & sel_one_hot_i[2];
  assign data_masked[1122] = data_i[1122] & sel_one_hot_i[2];
  assign data_masked[1121] = data_i[1121] & sel_one_hot_i[2];
  assign data_masked[1120] = data_i[1120] & sel_one_hot_i[2];
  assign data_masked[1119] = data_i[1119] & sel_one_hot_i[2];
  assign data_masked[1118] = data_i[1118] & sel_one_hot_i[2];
  assign data_masked[1117] = data_i[1117] & sel_one_hot_i[2];
  assign data_masked[1116] = data_i[1116] & sel_one_hot_i[2];
  assign data_masked[1115] = data_i[1115] & sel_one_hot_i[2];
  assign data_masked[1114] = data_i[1114] & sel_one_hot_i[2];
  assign data_masked[1113] = data_i[1113] & sel_one_hot_i[2];
  assign data_masked[1112] = data_i[1112] & sel_one_hot_i[2];
  assign data_masked[1111] = data_i[1111] & sel_one_hot_i[2];
  assign data_masked[1110] = data_i[1110] & sel_one_hot_i[2];
  assign data_masked[1109] = data_i[1109] & sel_one_hot_i[2];
  assign data_masked[1108] = data_i[1108] & sel_one_hot_i[2];
  assign data_masked[1107] = data_i[1107] & sel_one_hot_i[2];
  assign data_masked[1106] = data_i[1106] & sel_one_hot_i[2];
  assign data_masked[1105] = data_i[1105] & sel_one_hot_i[2];
  assign data_masked[1104] = data_i[1104] & sel_one_hot_i[2];
  assign data_masked[1103] = data_i[1103] & sel_one_hot_i[2];
  assign data_masked[1102] = data_i[1102] & sel_one_hot_i[2];
  assign data_masked[1101] = data_i[1101] & sel_one_hot_i[2];
  assign data_masked[1100] = data_i[1100] & sel_one_hot_i[2];
  assign data_masked[1099] = data_i[1099] & sel_one_hot_i[2];
  assign data_masked[1098] = data_i[1098] & sel_one_hot_i[2];
  assign data_masked[1097] = data_i[1097] & sel_one_hot_i[2];
  assign data_masked[1096] = data_i[1096] & sel_one_hot_i[2];
  assign data_masked[1095] = data_i[1095] & sel_one_hot_i[2];
  assign data_masked[1094] = data_i[1094] & sel_one_hot_i[2];
  assign data_masked[1093] = data_i[1093] & sel_one_hot_i[2];
  assign data_masked[1092] = data_i[1092] & sel_one_hot_i[2];
  assign data_masked[1091] = data_i[1091] & sel_one_hot_i[2];
  assign data_masked[1090] = data_i[1090] & sel_one_hot_i[2];
  assign data_masked[1089] = data_i[1089] & sel_one_hot_i[2];
  assign data_masked[1088] = data_i[1088] & sel_one_hot_i[2];
  assign data_masked[1087] = data_i[1087] & sel_one_hot_i[2];
  assign data_masked[1086] = data_i[1086] & sel_one_hot_i[2];
  assign data_masked[1085] = data_i[1085] & sel_one_hot_i[2];
  assign data_masked[1084] = data_i[1084] & sel_one_hot_i[2];
  assign data_masked[1083] = data_i[1083] & sel_one_hot_i[2];
  assign data_masked[1082] = data_i[1082] & sel_one_hot_i[2];
  assign data_masked[1081] = data_i[1081] & sel_one_hot_i[2];
  assign data_masked[1080] = data_i[1080] & sel_one_hot_i[2];
  assign data_masked[1079] = data_i[1079] & sel_one_hot_i[2];
  assign data_masked[1078] = data_i[1078] & sel_one_hot_i[2];
  assign data_masked[2155] = data_i[2155] & sel_one_hot_i[3];
  assign data_masked[2154] = data_i[2154] & sel_one_hot_i[3];
  assign data_masked[2153] = data_i[2153] & sel_one_hot_i[3];
  assign data_masked[2152] = data_i[2152] & sel_one_hot_i[3];
  assign data_masked[2151] = data_i[2151] & sel_one_hot_i[3];
  assign data_masked[2150] = data_i[2150] & sel_one_hot_i[3];
  assign data_masked[2149] = data_i[2149] & sel_one_hot_i[3];
  assign data_masked[2148] = data_i[2148] & sel_one_hot_i[3];
  assign data_masked[2147] = data_i[2147] & sel_one_hot_i[3];
  assign data_masked[2146] = data_i[2146] & sel_one_hot_i[3];
  assign data_masked[2145] = data_i[2145] & sel_one_hot_i[3];
  assign data_masked[2144] = data_i[2144] & sel_one_hot_i[3];
  assign data_masked[2143] = data_i[2143] & sel_one_hot_i[3];
  assign data_masked[2142] = data_i[2142] & sel_one_hot_i[3];
  assign data_masked[2141] = data_i[2141] & sel_one_hot_i[3];
  assign data_masked[2140] = data_i[2140] & sel_one_hot_i[3];
  assign data_masked[2139] = data_i[2139] & sel_one_hot_i[3];
  assign data_masked[2138] = data_i[2138] & sel_one_hot_i[3];
  assign data_masked[2137] = data_i[2137] & sel_one_hot_i[3];
  assign data_masked[2136] = data_i[2136] & sel_one_hot_i[3];
  assign data_masked[2135] = data_i[2135] & sel_one_hot_i[3];
  assign data_masked[2134] = data_i[2134] & sel_one_hot_i[3];
  assign data_masked[2133] = data_i[2133] & sel_one_hot_i[3];
  assign data_masked[2132] = data_i[2132] & sel_one_hot_i[3];
  assign data_masked[2131] = data_i[2131] & sel_one_hot_i[3];
  assign data_masked[2130] = data_i[2130] & sel_one_hot_i[3];
  assign data_masked[2129] = data_i[2129] & sel_one_hot_i[3];
  assign data_masked[2128] = data_i[2128] & sel_one_hot_i[3];
  assign data_masked[2127] = data_i[2127] & sel_one_hot_i[3];
  assign data_masked[2126] = data_i[2126] & sel_one_hot_i[3];
  assign data_masked[2125] = data_i[2125] & sel_one_hot_i[3];
  assign data_masked[2124] = data_i[2124] & sel_one_hot_i[3];
  assign data_masked[2123] = data_i[2123] & sel_one_hot_i[3];
  assign data_masked[2122] = data_i[2122] & sel_one_hot_i[3];
  assign data_masked[2121] = data_i[2121] & sel_one_hot_i[3];
  assign data_masked[2120] = data_i[2120] & sel_one_hot_i[3];
  assign data_masked[2119] = data_i[2119] & sel_one_hot_i[3];
  assign data_masked[2118] = data_i[2118] & sel_one_hot_i[3];
  assign data_masked[2117] = data_i[2117] & sel_one_hot_i[3];
  assign data_masked[2116] = data_i[2116] & sel_one_hot_i[3];
  assign data_masked[2115] = data_i[2115] & sel_one_hot_i[3];
  assign data_masked[2114] = data_i[2114] & sel_one_hot_i[3];
  assign data_masked[2113] = data_i[2113] & sel_one_hot_i[3];
  assign data_masked[2112] = data_i[2112] & sel_one_hot_i[3];
  assign data_masked[2111] = data_i[2111] & sel_one_hot_i[3];
  assign data_masked[2110] = data_i[2110] & sel_one_hot_i[3];
  assign data_masked[2109] = data_i[2109] & sel_one_hot_i[3];
  assign data_masked[2108] = data_i[2108] & sel_one_hot_i[3];
  assign data_masked[2107] = data_i[2107] & sel_one_hot_i[3];
  assign data_masked[2106] = data_i[2106] & sel_one_hot_i[3];
  assign data_masked[2105] = data_i[2105] & sel_one_hot_i[3];
  assign data_masked[2104] = data_i[2104] & sel_one_hot_i[3];
  assign data_masked[2103] = data_i[2103] & sel_one_hot_i[3];
  assign data_masked[2102] = data_i[2102] & sel_one_hot_i[3];
  assign data_masked[2101] = data_i[2101] & sel_one_hot_i[3];
  assign data_masked[2100] = data_i[2100] & sel_one_hot_i[3];
  assign data_masked[2099] = data_i[2099] & sel_one_hot_i[3];
  assign data_masked[2098] = data_i[2098] & sel_one_hot_i[3];
  assign data_masked[2097] = data_i[2097] & sel_one_hot_i[3];
  assign data_masked[2096] = data_i[2096] & sel_one_hot_i[3];
  assign data_masked[2095] = data_i[2095] & sel_one_hot_i[3];
  assign data_masked[2094] = data_i[2094] & sel_one_hot_i[3];
  assign data_masked[2093] = data_i[2093] & sel_one_hot_i[3];
  assign data_masked[2092] = data_i[2092] & sel_one_hot_i[3];
  assign data_masked[2091] = data_i[2091] & sel_one_hot_i[3];
  assign data_masked[2090] = data_i[2090] & sel_one_hot_i[3];
  assign data_masked[2089] = data_i[2089] & sel_one_hot_i[3];
  assign data_masked[2088] = data_i[2088] & sel_one_hot_i[3];
  assign data_masked[2087] = data_i[2087] & sel_one_hot_i[3];
  assign data_masked[2086] = data_i[2086] & sel_one_hot_i[3];
  assign data_masked[2085] = data_i[2085] & sel_one_hot_i[3];
  assign data_masked[2084] = data_i[2084] & sel_one_hot_i[3];
  assign data_masked[2083] = data_i[2083] & sel_one_hot_i[3];
  assign data_masked[2082] = data_i[2082] & sel_one_hot_i[3];
  assign data_masked[2081] = data_i[2081] & sel_one_hot_i[3];
  assign data_masked[2080] = data_i[2080] & sel_one_hot_i[3];
  assign data_masked[2079] = data_i[2079] & sel_one_hot_i[3];
  assign data_masked[2078] = data_i[2078] & sel_one_hot_i[3];
  assign data_masked[2077] = data_i[2077] & sel_one_hot_i[3];
  assign data_masked[2076] = data_i[2076] & sel_one_hot_i[3];
  assign data_masked[2075] = data_i[2075] & sel_one_hot_i[3];
  assign data_masked[2074] = data_i[2074] & sel_one_hot_i[3];
  assign data_masked[2073] = data_i[2073] & sel_one_hot_i[3];
  assign data_masked[2072] = data_i[2072] & sel_one_hot_i[3];
  assign data_masked[2071] = data_i[2071] & sel_one_hot_i[3];
  assign data_masked[2070] = data_i[2070] & sel_one_hot_i[3];
  assign data_masked[2069] = data_i[2069] & sel_one_hot_i[3];
  assign data_masked[2068] = data_i[2068] & sel_one_hot_i[3];
  assign data_masked[2067] = data_i[2067] & sel_one_hot_i[3];
  assign data_masked[2066] = data_i[2066] & sel_one_hot_i[3];
  assign data_masked[2065] = data_i[2065] & sel_one_hot_i[3];
  assign data_masked[2064] = data_i[2064] & sel_one_hot_i[3];
  assign data_masked[2063] = data_i[2063] & sel_one_hot_i[3];
  assign data_masked[2062] = data_i[2062] & sel_one_hot_i[3];
  assign data_masked[2061] = data_i[2061] & sel_one_hot_i[3];
  assign data_masked[2060] = data_i[2060] & sel_one_hot_i[3];
  assign data_masked[2059] = data_i[2059] & sel_one_hot_i[3];
  assign data_masked[2058] = data_i[2058] & sel_one_hot_i[3];
  assign data_masked[2057] = data_i[2057] & sel_one_hot_i[3];
  assign data_masked[2056] = data_i[2056] & sel_one_hot_i[3];
  assign data_masked[2055] = data_i[2055] & sel_one_hot_i[3];
  assign data_masked[2054] = data_i[2054] & sel_one_hot_i[3];
  assign data_masked[2053] = data_i[2053] & sel_one_hot_i[3];
  assign data_masked[2052] = data_i[2052] & sel_one_hot_i[3];
  assign data_masked[2051] = data_i[2051] & sel_one_hot_i[3];
  assign data_masked[2050] = data_i[2050] & sel_one_hot_i[3];
  assign data_masked[2049] = data_i[2049] & sel_one_hot_i[3];
  assign data_masked[2048] = data_i[2048] & sel_one_hot_i[3];
  assign data_masked[2047] = data_i[2047] & sel_one_hot_i[3];
  assign data_masked[2046] = data_i[2046] & sel_one_hot_i[3];
  assign data_masked[2045] = data_i[2045] & sel_one_hot_i[3];
  assign data_masked[2044] = data_i[2044] & sel_one_hot_i[3];
  assign data_masked[2043] = data_i[2043] & sel_one_hot_i[3];
  assign data_masked[2042] = data_i[2042] & sel_one_hot_i[3];
  assign data_masked[2041] = data_i[2041] & sel_one_hot_i[3];
  assign data_masked[2040] = data_i[2040] & sel_one_hot_i[3];
  assign data_masked[2039] = data_i[2039] & sel_one_hot_i[3];
  assign data_masked[2038] = data_i[2038] & sel_one_hot_i[3];
  assign data_masked[2037] = data_i[2037] & sel_one_hot_i[3];
  assign data_masked[2036] = data_i[2036] & sel_one_hot_i[3];
  assign data_masked[2035] = data_i[2035] & sel_one_hot_i[3];
  assign data_masked[2034] = data_i[2034] & sel_one_hot_i[3];
  assign data_masked[2033] = data_i[2033] & sel_one_hot_i[3];
  assign data_masked[2032] = data_i[2032] & sel_one_hot_i[3];
  assign data_masked[2031] = data_i[2031] & sel_one_hot_i[3];
  assign data_masked[2030] = data_i[2030] & sel_one_hot_i[3];
  assign data_masked[2029] = data_i[2029] & sel_one_hot_i[3];
  assign data_masked[2028] = data_i[2028] & sel_one_hot_i[3];
  assign data_masked[2027] = data_i[2027] & sel_one_hot_i[3];
  assign data_masked[2026] = data_i[2026] & sel_one_hot_i[3];
  assign data_masked[2025] = data_i[2025] & sel_one_hot_i[3];
  assign data_masked[2024] = data_i[2024] & sel_one_hot_i[3];
  assign data_masked[2023] = data_i[2023] & sel_one_hot_i[3];
  assign data_masked[2022] = data_i[2022] & sel_one_hot_i[3];
  assign data_masked[2021] = data_i[2021] & sel_one_hot_i[3];
  assign data_masked[2020] = data_i[2020] & sel_one_hot_i[3];
  assign data_masked[2019] = data_i[2019] & sel_one_hot_i[3];
  assign data_masked[2018] = data_i[2018] & sel_one_hot_i[3];
  assign data_masked[2017] = data_i[2017] & sel_one_hot_i[3];
  assign data_masked[2016] = data_i[2016] & sel_one_hot_i[3];
  assign data_masked[2015] = data_i[2015] & sel_one_hot_i[3];
  assign data_masked[2014] = data_i[2014] & sel_one_hot_i[3];
  assign data_masked[2013] = data_i[2013] & sel_one_hot_i[3];
  assign data_masked[2012] = data_i[2012] & sel_one_hot_i[3];
  assign data_masked[2011] = data_i[2011] & sel_one_hot_i[3];
  assign data_masked[2010] = data_i[2010] & sel_one_hot_i[3];
  assign data_masked[2009] = data_i[2009] & sel_one_hot_i[3];
  assign data_masked[2008] = data_i[2008] & sel_one_hot_i[3];
  assign data_masked[2007] = data_i[2007] & sel_one_hot_i[3];
  assign data_masked[2006] = data_i[2006] & sel_one_hot_i[3];
  assign data_masked[2005] = data_i[2005] & sel_one_hot_i[3];
  assign data_masked[2004] = data_i[2004] & sel_one_hot_i[3];
  assign data_masked[2003] = data_i[2003] & sel_one_hot_i[3];
  assign data_masked[2002] = data_i[2002] & sel_one_hot_i[3];
  assign data_masked[2001] = data_i[2001] & sel_one_hot_i[3];
  assign data_masked[2000] = data_i[2000] & sel_one_hot_i[3];
  assign data_masked[1999] = data_i[1999] & sel_one_hot_i[3];
  assign data_masked[1998] = data_i[1998] & sel_one_hot_i[3];
  assign data_masked[1997] = data_i[1997] & sel_one_hot_i[3];
  assign data_masked[1996] = data_i[1996] & sel_one_hot_i[3];
  assign data_masked[1995] = data_i[1995] & sel_one_hot_i[3];
  assign data_masked[1994] = data_i[1994] & sel_one_hot_i[3];
  assign data_masked[1993] = data_i[1993] & sel_one_hot_i[3];
  assign data_masked[1992] = data_i[1992] & sel_one_hot_i[3];
  assign data_masked[1991] = data_i[1991] & sel_one_hot_i[3];
  assign data_masked[1990] = data_i[1990] & sel_one_hot_i[3];
  assign data_masked[1989] = data_i[1989] & sel_one_hot_i[3];
  assign data_masked[1988] = data_i[1988] & sel_one_hot_i[3];
  assign data_masked[1987] = data_i[1987] & sel_one_hot_i[3];
  assign data_masked[1986] = data_i[1986] & sel_one_hot_i[3];
  assign data_masked[1985] = data_i[1985] & sel_one_hot_i[3];
  assign data_masked[1984] = data_i[1984] & sel_one_hot_i[3];
  assign data_masked[1983] = data_i[1983] & sel_one_hot_i[3];
  assign data_masked[1982] = data_i[1982] & sel_one_hot_i[3];
  assign data_masked[1981] = data_i[1981] & sel_one_hot_i[3];
  assign data_masked[1980] = data_i[1980] & sel_one_hot_i[3];
  assign data_masked[1979] = data_i[1979] & sel_one_hot_i[3];
  assign data_masked[1978] = data_i[1978] & sel_one_hot_i[3];
  assign data_masked[1977] = data_i[1977] & sel_one_hot_i[3];
  assign data_masked[1976] = data_i[1976] & sel_one_hot_i[3];
  assign data_masked[1975] = data_i[1975] & sel_one_hot_i[3];
  assign data_masked[1974] = data_i[1974] & sel_one_hot_i[3];
  assign data_masked[1973] = data_i[1973] & sel_one_hot_i[3];
  assign data_masked[1972] = data_i[1972] & sel_one_hot_i[3];
  assign data_masked[1971] = data_i[1971] & sel_one_hot_i[3];
  assign data_masked[1970] = data_i[1970] & sel_one_hot_i[3];
  assign data_masked[1969] = data_i[1969] & sel_one_hot_i[3];
  assign data_masked[1968] = data_i[1968] & sel_one_hot_i[3];
  assign data_masked[1967] = data_i[1967] & sel_one_hot_i[3];
  assign data_masked[1966] = data_i[1966] & sel_one_hot_i[3];
  assign data_masked[1965] = data_i[1965] & sel_one_hot_i[3];
  assign data_masked[1964] = data_i[1964] & sel_one_hot_i[3];
  assign data_masked[1963] = data_i[1963] & sel_one_hot_i[3];
  assign data_masked[1962] = data_i[1962] & sel_one_hot_i[3];
  assign data_masked[1961] = data_i[1961] & sel_one_hot_i[3];
  assign data_masked[1960] = data_i[1960] & sel_one_hot_i[3];
  assign data_masked[1959] = data_i[1959] & sel_one_hot_i[3];
  assign data_masked[1958] = data_i[1958] & sel_one_hot_i[3];
  assign data_masked[1957] = data_i[1957] & sel_one_hot_i[3];
  assign data_masked[1956] = data_i[1956] & sel_one_hot_i[3];
  assign data_masked[1955] = data_i[1955] & sel_one_hot_i[3];
  assign data_masked[1954] = data_i[1954] & sel_one_hot_i[3];
  assign data_masked[1953] = data_i[1953] & sel_one_hot_i[3];
  assign data_masked[1952] = data_i[1952] & sel_one_hot_i[3];
  assign data_masked[1951] = data_i[1951] & sel_one_hot_i[3];
  assign data_masked[1950] = data_i[1950] & sel_one_hot_i[3];
  assign data_masked[1949] = data_i[1949] & sel_one_hot_i[3];
  assign data_masked[1948] = data_i[1948] & sel_one_hot_i[3];
  assign data_masked[1947] = data_i[1947] & sel_one_hot_i[3];
  assign data_masked[1946] = data_i[1946] & sel_one_hot_i[3];
  assign data_masked[1945] = data_i[1945] & sel_one_hot_i[3];
  assign data_masked[1944] = data_i[1944] & sel_one_hot_i[3];
  assign data_masked[1943] = data_i[1943] & sel_one_hot_i[3];
  assign data_masked[1942] = data_i[1942] & sel_one_hot_i[3];
  assign data_masked[1941] = data_i[1941] & sel_one_hot_i[3];
  assign data_masked[1940] = data_i[1940] & sel_one_hot_i[3];
  assign data_masked[1939] = data_i[1939] & sel_one_hot_i[3];
  assign data_masked[1938] = data_i[1938] & sel_one_hot_i[3];
  assign data_masked[1937] = data_i[1937] & sel_one_hot_i[3];
  assign data_masked[1936] = data_i[1936] & sel_one_hot_i[3];
  assign data_masked[1935] = data_i[1935] & sel_one_hot_i[3];
  assign data_masked[1934] = data_i[1934] & sel_one_hot_i[3];
  assign data_masked[1933] = data_i[1933] & sel_one_hot_i[3];
  assign data_masked[1932] = data_i[1932] & sel_one_hot_i[3];
  assign data_masked[1931] = data_i[1931] & sel_one_hot_i[3];
  assign data_masked[1930] = data_i[1930] & sel_one_hot_i[3];
  assign data_masked[1929] = data_i[1929] & sel_one_hot_i[3];
  assign data_masked[1928] = data_i[1928] & sel_one_hot_i[3];
  assign data_masked[1927] = data_i[1927] & sel_one_hot_i[3];
  assign data_masked[1926] = data_i[1926] & sel_one_hot_i[3];
  assign data_masked[1925] = data_i[1925] & sel_one_hot_i[3];
  assign data_masked[1924] = data_i[1924] & sel_one_hot_i[3];
  assign data_masked[1923] = data_i[1923] & sel_one_hot_i[3];
  assign data_masked[1922] = data_i[1922] & sel_one_hot_i[3];
  assign data_masked[1921] = data_i[1921] & sel_one_hot_i[3];
  assign data_masked[1920] = data_i[1920] & sel_one_hot_i[3];
  assign data_masked[1919] = data_i[1919] & sel_one_hot_i[3];
  assign data_masked[1918] = data_i[1918] & sel_one_hot_i[3];
  assign data_masked[1917] = data_i[1917] & sel_one_hot_i[3];
  assign data_masked[1916] = data_i[1916] & sel_one_hot_i[3];
  assign data_masked[1915] = data_i[1915] & sel_one_hot_i[3];
  assign data_masked[1914] = data_i[1914] & sel_one_hot_i[3];
  assign data_masked[1913] = data_i[1913] & sel_one_hot_i[3];
  assign data_masked[1912] = data_i[1912] & sel_one_hot_i[3];
  assign data_masked[1911] = data_i[1911] & sel_one_hot_i[3];
  assign data_masked[1910] = data_i[1910] & sel_one_hot_i[3];
  assign data_masked[1909] = data_i[1909] & sel_one_hot_i[3];
  assign data_masked[1908] = data_i[1908] & sel_one_hot_i[3];
  assign data_masked[1907] = data_i[1907] & sel_one_hot_i[3];
  assign data_masked[1906] = data_i[1906] & sel_one_hot_i[3];
  assign data_masked[1905] = data_i[1905] & sel_one_hot_i[3];
  assign data_masked[1904] = data_i[1904] & sel_one_hot_i[3];
  assign data_masked[1903] = data_i[1903] & sel_one_hot_i[3];
  assign data_masked[1902] = data_i[1902] & sel_one_hot_i[3];
  assign data_masked[1901] = data_i[1901] & sel_one_hot_i[3];
  assign data_masked[1900] = data_i[1900] & sel_one_hot_i[3];
  assign data_masked[1899] = data_i[1899] & sel_one_hot_i[3];
  assign data_masked[1898] = data_i[1898] & sel_one_hot_i[3];
  assign data_masked[1897] = data_i[1897] & sel_one_hot_i[3];
  assign data_masked[1896] = data_i[1896] & sel_one_hot_i[3];
  assign data_masked[1895] = data_i[1895] & sel_one_hot_i[3];
  assign data_masked[1894] = data_i[1894] & sel_one_hot_i[3];
  assign data_masked[1893] = data_i[1893] & sel_one_hot_i[3];
  assign data_masked[1892] = data_i[1892] & sel_one_hot_i[3];
  assign data_masked[1891] = data_i[1891] & sel_one_hot_i[3];
  assign data_masked[1890] = data_i[1890] & sel_one_hot_i[3];
  assign data_masked[1889] = data_i[1889] & sel_one_hot_i[3];
  assign data_masked[1888] = data_i[1888] & sel_one_hot_i[3];
  assign data_masked[1887] = data_i[1887] & sel_one_hot_i[3];
  assign data_masked[1886] = data_i[1886] & sel_one_hot_i[3];
  assign data_masked[1885] = data_i[1885] & sel_one_hot_i[3];
  assign data_masked[1884] = data_i[1884] & sel_one_hot_i[3];
  assign data_masked[1883] = data_i[1883] & sel_one_hot_i[3];
  assign data_masked[1882] = data_i[1882] & sel_one_hot_i[3];
  assign data_masked[1881] = data_i[1881] & sel_one_hot_i[3];
  assign data_masked[1880] = data_i[1880] & sel_one_hot_i[3];
  assign data_masked[1879] = data_i[1879] & sel_one_hot_i[3];
  assign data_masked[1878] = data_i[1878] & sel_one_hot_i[3];
  assign data_masked[1877] = data_i[1877] & sel_one_hot_i[3];
  assign data_masked[1876] = data_i[1876] & sel_one_hot_i[3];
  assign data_masked[1875] = data_i[1875] & sel_one_hot_i[3];
  assign data_masked[1874] = data_i[1874] & sel_one_hot_i[3];
  assign data_masked[1873] = data_i[1873] & sel_one_hot_i[3];
  assign data_masked[1872] = data_i[1872] & sel_one_hot_i[3];
  assign data_masked[1871] = data_i[1871] & sel_one_hot_i[3];
  assign data_masked[1870] = data_i[1870] & sel_one_hot_i[3];
  assign data_masked[1869] = data_i[1869] & sel_one_hot_i[3];
  assign data_masked[1868] = data_i[1868] & sel_one_hot_i[3];
  assign data_masked[1867] = data_i[1867] & sel_one_hot_i[3];
  assign data_masked[1866] = data_i[1866] & sel_one_hot_i[3];
  assign data_masked[1865] = data_i[1865] & sel_one_hot_i[3];
  assign data_masked[1864] = data_i[1864] & sel_one_hot_i[3];
  assign data_masked[1863] = data_i[1863] & sel_one_hot_i[3];
  assign data_masked[1862] = data_i[1862] & sel_one_hot_i[3];
  assign data_masked[1861] = data_i[1861] & sel_one_hot_i[3];
  assign data_masked[1860] = data_i[1860] & sel_one_hot_i[3];
  assign data_masked[1859] = data_i[1859] & sel_one_hot_i[3];
  assign data_masked[1858] = data_i[1858] & sel_one_hot_i[3];
  assign data_masked[1857] = data_i[1857] & sel_one_hot_i[3];
  assign data_masked[1856] = data_i[1856] & sel_one_hot_i[3];
  assign data_masked[1855] = data_i[1855] & sel_one_hot_i[3];
  assign data_masked[1854] = data_i[1854] & sel_one_hot_i[3];
  assign data_masked[1853] = data_i[1853] & sel_one_hot_i[3];
  assign data_masked[1852] = data_i[1852] & sel_one_hot_i[3];
  assign data_masked[1851] = data_i[1851] & sel_one_hot_i[3];
  assign data_masked[1850] = data_i[1850] & sel_one_hot_i[3];
  assign data_masked[1849] = data_i[1849] & sel_one_hot_i[3];
  assign data_masked[1848] = data_i[1848] & sel_one_hot_i[3];
  assign data_masked[1847] = data_i[1847] & sel_one_hot_i[3];
  assign data_masked[1846] = data_i[1846] & sel_one_hot_i[3];
  assign data_masked[1845] = data_i[1845] & sel_one_hot_i[3];
  assign data_masked[1844] = data_i[1844] & sel_one_hot_i[3];
  assign data_masked[1843] = data_i[1843] & sel_one_hot_i[3];
  assign data_masked[1842] = data_i[1842] & sel_one_hot_i[3];
  assign data_masked[1841] = data_i[1841] & sel_one_hot_i[3];
  assign data_masked[1840] = data_i[1840] & sel_one_hot_i[3];
  assign data_masked[1839] = data_i[1839] & sel_one_hot_i[3];
  assign data_masked[1838] = data_i[1838] & sel_one_hot_i[3];
  assign data_masked[1837] = data_i[1837] & sel_one_hot_i[3];
  assign data_masked[1836] = data_i[1836] & sel_one_hot_i[3];
  assign data_masked[1835] = data_i[1835] & sel_one_hot_i[3];
  assign data_masked[1834] = data_i[1834] & sel_one_hot_i[3];
  assign data_masked[1833] = data_i[1833] & sel_one_hot_i[3];
  assign data_masked[1832] = data_i[1832] & sel_one_hot_i[3];
  assign data_masked[1831] = data_i[1831] & sel_one_hot_i[3];
  assign data_masked[1830] = data_i[1830] & sel_one_hot_i[3];
  assign data_masked[1829] = data_i[1829] & sel_one_hot_i[3];
  assign data_masked[1828] = data_i[1828] & sel_one_hot_i[3];
  assign data_masked[1827] = data_i[1827] & sel_one_hot_i[3];
  assign data_masked[1826] = data_i[1826] & sel_one_hot_i[3];
  assign data_masked[1825] = data_i[1825] & sel_one_hot_i[3];
  assign data_masked[1824] = data_i[1824] & sel_one_hot_i[3];
  assign data_masked[1823] = data_i[1823] & sel_one_hot_i[3];
  assign data_masked[1822] = data_i[1822] & sel_one_hot_i[3];
  assign data_masked[1821] = data_i[1821] & sel_one_hot_i[3];
  assign data_masked[1820] = data_i[1820] & sel_one_hot_i[3];
  assign data_masked[1819] = data_i[1819] & sel_one_hot_i[3];
  assign data_masked[1818] = data_i[1818] & sel_one_hot_i[3];
  assign data_masked[1817] = data_i[1817] & sel_one_hot_i[3];
  assign data_masked[1816] = data_i[1816] & sel_one_hot_i[3];
  assign data_masked[1815] = data_i[1815] & sel_one_hot_i[3];
  assign data_masked[1814] = data_i[1814] & sel_one_hot_i[3];
  assign data_masked[1813] = data_i[1813] & sel_one_hot_i[3];
  assign data_masked[1812] = data_i[1812] & sel_one_hot_i[3];
  assign data_masked[1811] = data_i[1811] & sel_one_hot_i[3];
  assign data_masked[1810] = data_i[1810] & sel_one_hot_i[3];
  assign data_masked[1809] = data_i[1809] & sel_one_hot_i[3];
  assign data_masked[1808] = data_i[1808] & sel_one_hot_i[3];
  assign data_masked[1807] = data_i[1807] & sel_one_hot_i[3];
  assign data_masked[1806] = data_i[1806] & sel_one_hot_i[3];
  assign data_masked[1805] = data_i[1805] & sel_one_hot_i[3];
  assign data_masked[1804] = data_i[1804] & sel_one_hot_i[3];
  assign data_masked[1803] = data_i[1803] & sel_one_hot_i[3];
  assign data_masked[1802] = data_i[1802] & sel_one_hot_i[3];
  assign data_masked[1801] = data_i[1801] & sel_one_hot_i[3];
  assign data_masked[1800] = data_i[1800] & sel_one_hot_i[3];
  assign data_masked[1799] = data_i[1799] & sel_one_hot_i[3];
  assign data_masked[1798] = data_i[1798] & sel_one_hot_i[3];
  assign data_masked[1797] = data_i[1797] & sel_one_hot_i[3];
  assign data_masked[1796] = data_i[1796] & sel_one_hot_i[3];
  assign data_masked[1795] = data_i[1795] & sel_one_hot_i[3];
  assign data_masked[1794] = data_i[1794] & sel_one_hot_i[3];
  assign data_masked[1793] = data_i[1793] & sel_one_hot_i[3];
  assign data_masked[1792] = data_i[1792] & sel_one_hot_i[3];
  assign data_masked[1791] = data_i[1791] & sel_one_hot_i[3];
  assign data_masked[1790] = data_i[1790] & sel_one_hot_i[3];
  assign data_masked[1789] = data_i[1789] & sel_one_hot_i[3];
  assign data_masked[1788] = data_i[1788] & sel_one_hot_i[3];
  assign data_masked[1787] = data_i[1787] & sel_one_hot_i[3];
  assign data_masked[1786] = data_i[1786] & sel_one_hot_i[3];
  assign data_masked[1785] = data_i[1785] & sel_one_hot_i[3];
  assign data_masked[1784] = data_i[1784] & sel_one_hot_i[3];
  assign data_masked[1783] = data_i[1783] & sel_one_hot_i[3];
  assign data_masked[1782] = data_i[1782] & sel_one_hot_i[3];
  assign data_masked[1781] = data_i[1781] & sel_one_hot_i[3];
  assign data_masked[1780] = data_i[1780] & sel_one_hot_i[3];
  assign data_masked[1779] = data_i[1779] & sel_one_hot_i[3];
  assign data_masked[1778] = data_i[1778] & sel_one_hot_i[3];
  assign data_masked[1777] = data_i[1777] & sel_one_hot_i[3];
  assign data_masked[1776] = data_i[1776] & sel_one_hot_i[3];
  assign data_masked[1775] = data_i[1775] & sel_one_hot_i[3];
  assign data_masked[1774] = data_i[1774] & sel_one_hot_i[3];
  assign data_masked[1773] = data_i[1773] & sel_one_hot_i[3];
  assign data_masked[1772] = data_i[1772] & sel_one_hot_i[3];
  assign data_masked[1771] = data_i[1771] & sel_one_hot_i[3];
  assign data_masked[1770] = data_i[1770] & sel_one_hot_i[3];
  assign data_masked[1769] = data_i[1769] & sel_one_hot_i[3];
  assign data_masked[1768] = data_i[1768] & sel_one_hot_i[3];
  assign data_masked[1767] = data_i[1767] & sel_one_hot_i[3];
  assign data_masked[1766] = data_i[1766] & sel_one_hot_i[3];
  assign data_masked[1765] = data_i[1765] & sel_one_hot_i[3];
  assign data_masked[1764] = data_i[1764] & sel_one_hot_i[3];
  assign data_masked[1763] = data_i[1763] & sel_one_hot_i[3];
  assign data_masked[1762] = data_i[1762] & sel_one_hot_i[3];
  assign data_masked[1761] = data_i[1761] & sel_one_hot_i[3];
  assign data_masked[1760] = data_i[1760] & sel_one_hot_i[3];
  assign data_masked[1759] = data_i[1759] & sel_one_hot_i[3];
  assign data_masked[1758] = data_i[1758] & sel_one_hot_i[3];
  assign data_masked[1757] = data_i[1757] & sel_one_hot_i[3];
  assign data_masked[1756] = data_i[1756] & sel_one_hot_i[3];
  assign data_masked[1755] = data_i[1755] & sel_one_hot_i[3];
  assign data_masked[1754] = data_i[1754] & sel_one_hot_i[3];
  assign data_masked[1753] = data_i[1753] & sel_one_hot_i[3];
  assign data_masked[1752] = data_i[1752] & sel_one_hot_i[3];
  assign data_masked[1751] = data_i[1751] & sel_one_hot_i[3];
  assign data_masked[1750] = data_i[1750] & sel_one_hot_i[3];
  assign data_masked[1749] = data_i[1749] & sel_one_hot_i[3];
  assign data_masked[1748] = data_i[1748] & sel_one_hot_i[3];
  assign data_masked[1747] = data_i[1747] & sel_one_hot_i[3];
  assign data_masked[1746] = data_i[1746] & sel_one_hot_i[3];
  assign data_masked[1745] = data_i[1745] & sel_one_hot_i[3];
  assign data_masked[1744] = data_i[1744] & sel_one_hot_i[3];
  assign data_masked[1743] = data_i[1743] & sel_one_hot_i[3];
  assign data_masked[1742] = data_i[1742] & sel_one_hot_i[3];
  assign data_masked[1741] = data_i[1741] & sel_one_hot_i[3];
  assign data_masked[1740] = data_i[1740] & sel_one_hot_i[3];
  assign data_masked[1739] = data_i[1739] & sel_one_hot_i[3];
  assign data_masked[1738] = data_i[1738] & sel_one_hot_i[3];
  assign data_masked[1737] = data_i[1737] & sel_one_hot_i[3];
  assign data_masked[1736] = data_i[1736] & sel_one_hot_i[3];
  assign data_masked[1735] = data_i[1735] & sel_one_hot_i[3];
  assign data_masked[1734] = data_i[1734] & sel_one_hot_i[3];
  assign data_masked[1733] = data_i[1733] & sel_one_hot_i[3];
  assign data_masked[1732] = data_i[1732] & sel_one_hot_i[3];
  assign data_masked[1731] = data_i[1731] & sel_one_hot_i[3];
  assign data_masked[1730] = data_i[1730] & sel_one_hot_i[3];
  assign data_masked[1729] = data_i[1729] & sel_one_hot_i[3];
  assign data_masked[1728] = data_i[1728] & sel_one_hot_i[3];
  assign data_masked[1727] = data_i[1727] & sel_one_hot_i[3];
  assign data_masked[1726] = data_i[1726] & sel_one_hot_i[3];
  assign data_masked[1725] = data_i[1725] & sel_one_hot_i[3];
  assign data_masked[1724] = data_i[1724] & sel_one_hot_i[3];
  assign data_masked[1723] = data_i[1723] & sel_one_hot_i[3];
  assign data_masked[1722] = data_i[1722] & sel_one_hot_i[3];
  assign data_masked[1721] = data_i[1721] & sel_one_hot_i[3];
  assign data_masked[1720] = data_i[1720] & sel_one_hot_i[3];
  assign data_masked[1719] = data_i[1719] & sel_one_hot_i[3];
  assign data_masked[1718] = data_i[1718] & sel_one_hot_i[3];
  assign data_masked[1717] = data_i[1717] & sel_one_hot_i[3];
  assign data_masked[1716] = data_i[1716] & sel_one_hot_i[3];
  assign data_masked[1715] = data_i[1715] & sel_one_hot_i[3];
  assign data_masked[1714] = data_i[1714] & sel_one_hot_i[3];
  assign data_masked[1713] = data_i[1713] & sel_one_hot_i[3];
  assign data_masked[1712] = data_i[1712] & sel_one_hot_i[3];
  assign data_masked[1711] = data_i[1711] & sel_one_hot_i[3];
  assign data_masked[1710] = data_i[1710] & sel_one_hot_i[3];
  assign data_masked[1709] = data_i[1709] & sel_one_hot_i[3];
  assign data_masked[1708] = data_i[1708] & sel_one_hot_i[3];
  assign data_masked[1707] = data_i[1707] & sel_one_hot_i[3];
  assign data_masked[1706] = data_i[1706] & sel_one_hot_i[3];
  assign data_masked[1705] = data_i[1705] & sel_one_hot_i[3];
  assign data_masked[1704] = data_i[1704] & sel_one_hot_i[3];
  assign data_masked[1703] = data_i[1703] & sel_one_hot_i[3];
  assign data_masked[1702] = data_i[1702] & sel_one_hot_i[3];
  assign data_masked[1701] = data_i[1701] & sel_one_hot_i[3];
  assign data_masked[1700] = data_i[1700] & sel_one_hot_i[3];
  assign data_masked[1699] = data_i[1699] & sel_one_hot_i[3];
  assign data_masked[1698] = data_i[1698] & sel_one_hot_i[3];
  assign data_masked[1697] = data_i[1697] & sel_one_hot_i[3];
  assign data_masked[1696] = data_i[1696] & sel_one_hot_i[3];
  assign data_masked[1695] = data_i[1695] & sel_one_hot_i[3];
  assign data_masked[1694] = data_i[1694] & sel_one_hot_i[3];
  assign data_masked[1693] = data_i[1693] & sel_one_hot_i[3];
  assign data_masked[1692] = data_i[1692] & sel_one_hot_i[3];
  assign data_masked[1691] = data_i[1691] & sel_one_hot_i[3];
  assign data_masked[1690] = data_i[1690] & sel_one_hot_i[3];
  assign data_masked[1689] = data_i[1689] & sel_one_hot_i[3];
  assign data_masked[1688] = data_i[1688] & sel_one_hot_i[3];
  assign data_masked[1687] = data_i[1687] & sel_one_hot_i[3];
  assign data_masked[1686] = data_i[1686] & sel_one_hot_i[3];
  assign data_masked[1685] = data_i[1685] & sel_one_hot_i[3];
  assign data_masked[1684] = data_i[1684] & sel_one_hot_i[3];
  assign data_masked[1683] = data_i[1683] & sel_one_hot_i[3];
  assign data_masked[1682] = data_i[1682] & sel_one_hot_i[3];
  assign data_masked[1681] = data_i[1681] & sel_one_hot_i[3];
  assign data_masked[1680] = data_i[1680] & sel_one_hot_i[3];
  assign data_masked[1679] = data_i[1679] & sel_one_hot_i[3];
  assign data_masked[1678] = data_i[1678] & sel_one_hot_i[3];
  assign data_masked[1677] = data_i[1677] & sel_one_hot_i[3];
  assign data_masked[1676] = data_i[1676] & sel_one_hot_i[3];
  assign data_masked[1675] = data_i[1675] & sel_one_hot_i[3];
  assign data_masked[1674] = data_i[1674] & sel_one_hot_i[3];
  assign data_masked[1673] = data_i[1673] & sel_one_hot_i[3];
  assign data_masked[1672] = data_i[1672] & sel_one_hot_i[3];
  assign data_masked[1671] = data_i[1671] & sel_one_hot_i[3];
  assign data_masked[1670] = data_i[1670] & sel_one_hot_i[3];
  assign data_masked[1669] = data_i[1669] & sel_one_hot_i[3];
  assign data_masked[1668] = data_i[1668] & sel_one_hot_i[3];
  assign data_masked[1667] = data_i[1667] & sel_one_hot_i[3];
  assign data_masked[1666] = data_i[1666] & sel_one_hot_i[3];
  assign data_masked[1665] = data_i[1665] & sel_one_hot_i[3];
  assign data_masked[1664] = data_i[1664] & sel_one_hot_i[3];
  assign data_masked[1663] = data_i[1663] & sel_one_hot_i[3];
  assign data_masked[1662] = data_i[1662] & sel_one_hot_i[3];
  assign data_masked[1661] = data_i[1661] & sel_one_hot_i[3];
  assign data_masked[1660] = data_i[1660] & sel_one_hot_i[3];
  assign data_masked[1659] = data_i[1659] & sel_one_hot_i[3];
  assign data_masked[1658] = data_i[1658] & sel_one_hot_i[3];
  assign data_masked[1657] = data_i[1657] & sel_one_hot_i[3];
  assign data_masked[1656] = data_i[1656] & sel_one_hot_i[3];
  assign data_masked[1655] = data_i[1655] & sel_one_hot_i[3];
  assign data_masked[1654] = data_i[1654] & sel_one_hot_i[3];
  assign data_masked[1653] = data_i[1653] & sel_one_hot_i[3];
  assign data_masked[1652] = data_i[1652] & sel_one_hot_i[3];
  assign data_masked[1651] = data_i[1651] & sel_one_hot_i[3];
  assign data_masked[1650] = data_i[1650] & sel_one_hot_i[3];
  assign data_masked[1649] = data_i[1649] & sel_one_hot_i[3];
  assign data_masked[1648] = data_i[1648] & sel_one_hot_i[3];
  assign data_masked[1647] = data_i[1647] & sel_one_hot_i[3];
  assign data_masked[1646] = data_i[1646] & sel_one_hot_i[3];
  assign data_masked[1645] = data_i[1645] & sel_one_hot_i[3];
  assign data_masked[1644] = data_i[1644] & sel_one_hot_i[3];
  assign data_masked[1643] = data_i[1643] & sel_one_hot_i[3];
  assign data_masked[1642] = data_i[1642] & sel_one_hot_i[3];
  assign data_masked[1641] = data_i[1641] & sel_one_hot_i[3];
  assign data_masked[1640] = data_i[1640] & sel_one_hot_i[3];
  assign data_masked[1639] = data_i[1639] & sel_one_hot_i[3];
  assign data_masked[1638] = data_i[1638] & sel_one_hot_i[3];
  assign data_masked[1637] = data_i[1637] & sel_one_hot_i[3];
  assign data_masked[1636] = data_i[1636] & sel_one_hot_i[3];
  assign data_masked[1635] = data_i[1635] & sel_one_hot_i[3];
  assign data_masked[1634] = data_i[1634] & sel_one_hot_i[3];
  assign data_masked[1633] = data_i[1633] & sel_one_hot_i[3];
  assign data_masked[1632] = data_i[1632] & sel_one_hot_i[3];
  assign data_masked[1631] = data_i[1631] & sel_one_hot_i[3];
  assign data_masked[1630] = data_i[1630] & sel_one_hot_i[3];
  assign data_masked[1629] = data_i[1629] & sel_one_hot_i[3];
  assign data_masked[1628] = data_i[1628] & sel_one_hot_i[3];
  assign data_masked[1627] = data_i[1627] & sel_one_hot_i[3];
  assign data_masked[1626] = data_i[1626] & sel_one_hot_i[3];
  assign data_masked[1625] = data_i[1625] & sel_one_hot_i[3];
  assign data_masked[1624] = data_i[1624] & sel_one_hot_i[3];
  assign data_masked[1623] = data_i[1623] & sel_one_hot_i[3];
  assign data_masked[1622] = data_i[1622] & sel_one_hot_i[3];
  assign data_masked[1621] = data_i[1621] & sel_one_hot_i[3];
  assign data_masked[1620] = data_i[1620] & sel_one_hot_i[3];
  assign data_masked[1619] = data_i[1619] & sel_one_hot_i[3];
  assign data_masked[1618] = data_i[1618] & sel_one_hot_i[3];
  assign data_masked[1617] = data_i[1617] & sel_one_hot_i[3];
  assign data_masked[2694] = data_i[2694] & sel_one_hot_i[4];
  assign data_masked[2693] = data_i[2693] & sel_one_hot_i[4];
  assign data_masked[2692] = data_i[2692] & sel_one_hot_i[4];
  assign data_masked[2691] = data_i[2691] & sel_one_hot_i[4];
  assign data_masked[2690] = data_i[2690] & sel_one_hot_i[4];
  assign data_masked[2689] = data_i[2689] & sel_one_hot_i[4];
  assign data_masked[2688] = data_i[2688] & sel_one_hot_i[4];
  assign data_masked[2687] = data_i[2687] & sel_one_hot_i[4];
  assign data_masked[2686] = data_i[2686] & sel_one_hot_i[4];
  assign data_masked[2685] = data_i[2685] & sel_one_hot_i[4];
  assign data_masked[2684] = data_i[2684] & sel_one_hot_i[4];
  assign data_masked[2683] = data_i[2683] & sel_one_hot_i[4];
  assign data_masked[2682] = data_i[2682] & sel_one_hot_i[4];
  assign data_masked[2681] = data_i[2681] & sel_one_hot_i[4];
  assign data_masked[2680] = data_i[2680] & sel_one_hot_i[4];
  assign data_masked[2679] = data_i[2679] & sel_one_hot_i[4];
  assign data_masked[2678] = data_i[2678] & sel_one_hot_i[4];
  assign data_masked[2677] = data_i[2677] & sel_one_hot_i[4];
  assign data_masked[2676] = data_i[2676] & sel_one_hot_i[4];
  assign data_masked[2675] = data_i[2675] & sel_one_hot_i[4];
  assign data_masked[2674] = data_i[2674] & sel_one_hot_i[4];
  assign data_masked[2673] = data_i[2673] & sel_one_hot_i[4];
  assign data_masked[2672] = data_i[2672] & sel_one_hot_i[4];
  assign data_masked[2671] = data_i[2671] & sel_one_hot_i[4];
  assign data_masked[2670] = data_i[2670] & sel_one_hot_i[4];
  assign data_masked[2669] = data_i[2669] & sel_one_hot_i[4];
  assign data_masked[2668] = data_i[2668] & sel_one_hot_i[4];
  assign data_masked[2667] = data_i[2667] & sel_one_hot_i[4];
  assign data_masked[2666] = data_i[2666] & sel_one_hot_i[4];
  assign data_masked[2665] = data_i[2665] & sel_one_hot_i[4];
  assign data_masked[2664] = data_i[2664] & sel_one_hot_i[4];
  assign data_masked[2663] = data_i[2663] & sel_one_hot_i[4];
  assign data_masked[2662] = data_i[2662] & sel_one_hot_i[4];
  assign data_masked[2661] = data_i[2661] & sel_one_hot_i[4];
  assign data_masked[2660] = data_i[2660] & sel_one_hot_i[4];
  assign data_masked[2659] = data_i[2659] & sel_one_hot_i[4];
  assign data_masked[2658] = data_i[2658] & sel_one_hot_i[4];
  assign data_masked[2657] = data_i[2657] & sel_one_hot_i[4];
  assign data_masked[2656] = data_i[2656] & sel_one_hot_i[4];
  assign data_masked[2655] = data_i[2655] & sel_one_hot_i[4];
  assign data_masked[2654] = data_i[2654] & sel_one_hot_i[4];
  assign data_masked[2653] = data_i[2653] & sel_one_hot_i[4];
  assign data_masked[2652] = data_i[2652] & sel_one_hot_i[4];
  assign data_masked[2651] = data_i[2651] & sel_one_hot_i[4];
  assign data_masked[2650] = data_i[2650] & sel_one_hot_i[4];
  assign data_masked[2649] = data_i[2649] & sel_one_hot_i[4];
  assign data_masked[2648] = data_i[2648] & sel_one_hot_i[4];
  assign data_masked[2647] = data_i[2647] & sel_one_hot_i[4];
  assign data_masked[2646] = data_i[2646] & sel_one_hot_i[4];
  assign data_masked[2645] = data_i[2645] & sel_one_hot_i[4];
  assign data_masked[2644] = data_i[2644] & sel_one_hot_i[4];
  assign data_masked[2643] = data_i[2643] & sel_one_hot_i[4];
  assign data_masked[2642] = data_i[2642] & sel_one_hot_i[4];
  assign data_masked[2641] = data_i[2641] & sel_one_hot_i[4];
  assign data_masked[2640] = data_i[2640] & sel_one_hot_i[4];
  assign data_masked[2639] = data_i[2639] & sel_one_hot_i[4];
  assign data_masked[2638] = data_i[2638] & sel_one_hot_i[4];
  assign data_masked[2637] = data_i[2637] & sel_one_hot_i[4];
  assign data_masked[2636] = data_i[2636] & sel_one_hot_i[4];
  assign data_masked[2635] = data_i[2635] & sel_one_hot_i[4];
  assign data_masked[2634] = data_i[2634] & sel_one_hot_i[4];
  assign data_masked[2633] = data_i[2633] & sel_one_hot_i[4];
  assign data_masked[2632] = data_i[2632] & sel_one_hot_i[4];
  assign data_masked[2631] = data_i[2631] & sel_one_hot_i[4];
  assign data_masked[2630] = data_i[2630] & sel_one_hot_i[4];
  assign data_masked[2629] = data_i[2629] & sel_one_hot_i[4];
  assign data_masked[2628] = data_i[2628] & sel_one_hot_i[4];
  assign data_masked[2627] = data_i[2627] & sel_one_hot_i[4];
  assign data_masked[2626] = data_i[2626] & sel_one_hot_i[4];
  assign data_masked[2625] = data_i[2625] & sel_one_hot_i[4];
  assign data_masked[2624] = data_i[2624] & sel_one_hot_i[4];
  assign data_masked[2623] = data_i[2623] & sel_one_hot_i[4];
  assign data_masked[2622] = data_i[2622] & sel_one_hot_i[4];
  assign data_masked[2621] = data_i[2621] & sel_one_hot_i[4];
  assign data_masked[2620] = data_i[2620] & sel_one_hot_i[4];
  assign data_masked[2619] = data_i[2619] & sel_one_hot_i[4];
  assign data_masked[2618] = data_i[2618] & sel_one_hot_i[4];
  assign data_masked[2617] = data_i[2617] & sel_one_hot_i[4];
  assign data_masked[2616] = data_i[2616] & sel_one_hot_i[4];
  assign data_masked[2615] = data_i[2615] & sel_one_hot_i[4];
  assign data_masked[2614] = data_i[2614] & sel_one_hot_i[4];
  assign data_masked[2613] = data_i[2613] & sel_one_hot_i[4];
  assign data_masked[2612] = data_i[2612] & sel_one_hot_i[4];
  assign data_masked[2611] = data_i[2611] & sel_one_hot_i[4];
  assign data_masked[2610] = data_i[2610] & sel_one_hot_i[4];
  assign data_masked[2609] = data_i[2609] & sel_one_hot_i[4];
  assign data_masked[2608] = data_i[2608] & sel_one_hot_i[4];
  assign data_masked[2607] = data_i[2607] & sel_one_hot_i[4];
  assign data_masked[2606] = data_i[2606] & sel_one_hot_i[4];
  assign data_masked[2605] = data_i[2605] & sel_one_hot_i[4];
  assign data_masked[2604] = data_i[2604] & sel_one_hot_i[4];
  assign data_masked[2603] = data_i[2603] & sel_one_hot_i[4];
  assign data_masked[2602] = data_i[2602] & sel_one_hot_i[4];
  assign data_masked[2601] = data_i[2601] & sel_one_hot_i[4];
  assign data_masked[2600] = data_i[2600] & sel_one_hot_i[4];
  assign data_masked[2599] = data_i[2599] & sel_one_hot_i[4];
  assign data_masked[2598] = data_i[2598] & sel_one_hot_i[4];
  assign data_masked[2597] = data_i[2597] & sel_one_hot_i[4];
  assign data_masked[2596] = data_i[2596] & sel_one_hot_i[4];
  assign data_masked[2595] = data_i[2595] & sel_one_hot_i[4];
  assign data_masked[2594] = data_i[2594] & sel_one_hot_i[4];
  assign data_masked[2593] = data_i[2593] & sel_one_hot_i[4];
  assign data_masked[2592] = data_i[2592] & sel_one_hot_i[4];
  assign data_masked[2591] = data_i[2591] & sel_one_hot_i[4];
  assign data_masked[2590] = data_i[2590] & sel_one_hot_i[4];
  assign data_masked[2589] = data_i[2589] & sel_one_hot_i[4];
  assign data_masked[2588] = data_i[2588] & sel_one_hot_i[4];
  assign data_masked[2587] = data_i[2587] & sel_one_hot_i[4];
  assign data_masked[2586] = data_i[2586] & sel_one_hot_i[4];
  assign data_masked[2585] = data_i[2585] & sel_one_hot_i[4];
  assign data_masked[2584] = data_i[2584] & sel_one_hot_i[4];
  assign data_masked[2583] = data_i[2583] & sel_one_hot_i[4];
  assign data_masked[2582] = data_i[2582] & sel_one_hot_i[4];
  assign data_masked[2581] = data_i[2581] & sel_one_hot_i[4];
  assign data_masked[2580] = data_i[2580] & sel_one_hot_i[4];
  assign data_masked[2579] = data_i[2579] & sel_one_hot_i[4];
  assign data_masked[2578] = data_i[2578] & sel_one_hot_i[4];
  assign data_masked[2577] = data_i[2577] & sel_one_hot_i[4];
  assign data_masked[2576] = data_i[2576] & sel_one_hot_i[4];
  assign data_masked[2575] = data_i[2575] & sel_one_hot_i[4];
  assign data_masked[2574] = data_i[2574] & sel_one_hot_i[4];
  assign data_masked[2573] = data_i[2573] & sel_one_hot_i[4];
  assign data_masked[2572] = data_i[2572] & sel_one_hot_i[4];
  assign data_masked[2571] = data_i[2571] & sel_one_hot_i[4];
  assign data_masked[2570] = data_i[2570] & sel_one_hot_i[4];
  assign data_masked[2569] = data_i[2569] & sel_one_hot_i[4];
  assign data_masked[2568] = data_i[2568] & sel_one_hot_i[4];
  assign data_masked[2567] = data_i[2567] & sel_one_hot_i[4];
  assign data_masked[2566] = data_i[2566] & sel_one_hot_i[4];
  assign data_masked[2565] = data_i[2565] & sel_one_hot_i[4];
  assign data_masked[2564] = data_i[2564] & sel_one_hot_i[4];
  assign data_masked[2563] = data_i[2563] & sel_one_hot_i[4];
  assign data_masked[2562] = data_i[2562] & sel_one_hot_i[4];
  assign data_masked[2561] = data_i[2561] & sel_one_hot_i[4];
  assign data_masked[2560] = data_i[2560] & sel_one_hot_i[4];
  assign data_masked[2559] = data_i[2559] & sel_one_hot_i[4];
  assign data_masked[2558] = data_i[2558] & sel_one_hot_i[4];
  assign data_masked[2557] = data_i[2557] & sel_one_hot_i[4];
  assign data_masked[2556] = data_i[2556] & sel_one_hot_i[4];
  assign data_masked[2555] = data_i[2555] & sel_one_hot_i[4];
  assign data_masked[2554] = data_i[2554] & sel_one_hot_i[4];
  assign data_masked[2553] = data_i[2553] & sel_one_hot_i[4];
  assign data_masked[2552] = data_i[2552] & sel_one_hot_i[4];
  assign data_masked[2551] = data_i[2551] & sel_one_hot_i[4];
  assign data_masked[2550] = data_i[2550] & sel_one_hot_i[4];
  assign data_masked[2549] = data_i[2549] & sel_one_hot_i[4];
  assign data_masked[2548] = data_i[2548] & sel_one_hot_i[4];
  assign data_masked[2547] = data_i[2547] & sel_one_hot_i[4];
  assign data_masked[2546] = data_i[2546] & sel_one_hot_i[4];
  assign data_masked[2545] = data_i[2545] & sel_one_hot_i[4];
  assign data_masked[2544] = data_i[2544] & sel_one_hot_i[4];
  assign data_masked[2543] = data_i[2543] & sel_one_hot_i[4];
  assign data_masked[2542] = data_i[2542] & sel_one_hot_i[4];
  assign data_masked[2541] = data_i[2541] & sel_one_hot_i[4];
  assign data_masked[2540] = data_i[2540] & sel_one_hot_i[4];
  assign data_masked[2539] = data_i[2539] & sel_one_hot_i[4];
  assign data_masked[2538] = data_i[2538] & sel_one_hot_i[4];
  assign data_masked[2537] = data_i[2537] & sel_one_hot_i[4];
  assign data_masked[2536] = data_i[2536] & sel_one_hot_i[4];
  assign data_masked[2535] = data_i[2535] & sel_one_hot_i[4];
  assign data_masked[2534] = data_i[2534] & sel_one_hot_i[4];
  assign data_masked[2533] = data_i[2533] & sel_one_hot_i[4];
  assign data_masked[2532] = data_i[2532] & sel_one_hot_i[4];
  assign data_masked[2531] = data_i[2531] & sel_one_hot_i[4];
  assign data_masked[2530] = data_i[2530] & sel_one_hot_i[4];
  assign data_masked[2529] = data_i[2529] & sel_one_hot_i[4];
  assign data_masked[2528] = data_i[2528] & sel_one_hot_i[4];
  assign data_masked[2527] = data_i[2527] & sel_one_hot_i[4];
  assign data_masked[2526] = data_i[2526] & sel_one_hot_i[4];
  assign data_masked[2525] = data_i[2525] & sel_one_hot_i[4];
  assign data_masked[2524] = data_i[2524] & sel_one_hot_i[4];
  assign data_masked[2523] = data_i[2523] & sel_one_hot_i[4];
  assign data_masked[2522] = data_i[2522] & sel_one_hot_i[4];
  assign data_masked[2521] = data_i[2521] & sel_one_hot_i[4];
  assign data_masked[2520] = data_i[2520] & sel_one_hot_i[4];
  assign data_masked[2519] = data_i[2519] & sel_one_hot_i[4];
  assign data_masked[2518] = data_i[2518] & sel_one_hot_i[4];
  assign data_masked[2517] = data_i[2517] & sel_one_hot_i[4];
  assign data_masked[2516] = data_i[2516] & sel_one_hot_i[4];
  assign data_masked[2515] = data_i[2515] & sel_one_hot_i[4];
  assign data_masked[2514] = data_i[2514] & sel_one_hot_i[4];
  assign data_masked[2513] = data_i[2513] & sel_one_hot_i[4];
  assign data_masked[2512] = data_i[2512] & sel_one_hot_i[4];
  assign data_masked[2511] = data_i[2511] & sel_one_hot_i[4];
  assign data_masked[2510] = data_i[2510] & sel_one_hot_i[4];
  assign data_masked[2509] = data_i[2509] & sel_one_hot_i[4];
  assign data_masked[2508] = data_i[2508] & sel_one_hot_i[4];
  assign data_masked[2507] = data_i[2507] & sel_one_hot_i[4];
  assign data_masked[2506] = data_i[2506] & sel_one_hot_i[4];
  assign data_masked[2505] = data_i[2505] & sel_one_hot_i[4];
  assign data_masked[2504] = data_i[2504] & sel_one_hot_i[4];
  assign data_masked[2503] = data_i[2503] & sel_one_hot_i[4];
  assign data_masked[2502] = data_i[2502] & sel_one_hot_i[4];
  assign data_masked[2501] = data_i[2501] & sel_one_hot_i[4];
  assign data_masked[2500] = data_i[2500] & sel_one_hot_i[4];
  assign data_masked[2499] = data_i[2499] & sel_one_hot_i[4];
  assign data_masked[2498] = data_i[2498] & sel_one_hot_i[4];
  assign data_masked[2497] = data_i[2497] & sel_one_hot_i[4];
  assign data_masked[2496] = data_i[2496] & sel_one_hot_i[4];
  assign data_masked[2495] = data_i[2495] & sel_one_hot_i[4];
  assign data_masked[2494] = data_i[2494] & sel_one_hot_i[4];
  assign data_masked[2493] = data_i[2493] & sel_one_hot_i[4];
  assign data_masked[2492] = data_i[2492] & sel_one_hot_i[4];
  assign data_masked[2491] = data_i[2491] & sel_one_hot_i[4];
  assign data_masked[2490] = data_i[2490] & sel_one_hot_i[4];
  assign data_masked[2489] = data_i[2489] & sel_one_hot_i[4];
  assign data_masked[2488] = data_i[2488] & sel_one_hot_i[4];
  assign data_masked[2487] = data_i[2487] & sel_one_hot_i[4];
  assign data_masked[2486] = data_i[2486] & sel_one_hot_i[4];
  assign data_masked[2485] = data_i[2485] & sel_one_hot_i[4];
  assign data_masked[2484] = data_i[2484] & sel_one_hot_i[4];
  assign data_masked[2483] = data_i[2483] & sel_one_hot_i[4];
  assign data_masked[2482] = data_i[2482] & sel_one_hot_i[4];
  assign data_masked[2481] = data_i[2481] & sel_one_hot_i[4];
  assign data_masked[2480] = data_i[2480] & sel_one_hot_i[4];
  assign data_masked[2479] = data_i[2479] & sel_one_hot_i[4];
  assign data_masked[2478] = data_i[2478] & sel_one_hot_i[4];
  assign data_masked[2477] = data_i[2477] & sel_one_hot_i[4];
  assign data_masked[2476] = data_i[2476] & sel_one_hot_i[4];
  assign data_masked[2475] = data_i[2475] & sel_one_hot_i[4];
  assign data_masked[2474] = data_i[2474] & sel_one_hot_i[4];
  assign data_masked[2473] = data_i[2473] & sel_one_hot_i[4];
  assign data_masked[2472] = data_i[2472] & sel_one_hot_i[4];
  assign data_masked[2471] = data_i[2471] & sel_one_hot_i[4];
  assign data_masked[2470] = data_i[2470] & sel_one_hot_i[4];
  assign data_masked[2469] = data_i[2469] & sel_one_hot_i[4];
  assign data_masked[2468] = data_i[2468] & sel_one_hot_i[4];
  assign data_masked[2467] = data_i[2467] & sel_one_hot_i[4];
  assign data_masked[2466] = data_i[2466] & sel_one_hot_i[4];
  assign data_masked[2465] = data_i[2465] & sel_one_hot_i[4];
  assign data_masked[2464] = data_i[2464] & sel_one_hot_i[4];
  assign data_masked[2463] = data_i[2463] & sel_one_hot_i[4];
  assign data_masked[2462] = data_i[2462] & sel_one_hot_i[4];
  assign data_masked[2461] = data_i[2461] & sel_one_hot_i[4];
  assign data_masked[2460] = data_i[2460] & sel_one_hot_i[4];
  assign data_masked[2459] = data_i[2459] & sel_one_hot_i[4];
  assign data_masked[2458] = data_i[2458] & sel_one_hot_i[4];
  assign data_masked[2457] = data_i[2457] & sel_one_hot_i[4];
  assign data_masked[2456] = data_i[2456] & sel_one_hot_i[4];
  assign data_masked[2455] = data_i[2455] & sel_one_hot_i[4];
  assign data_masked[2454] = data_i[2454] & sel_one_hot_i[4];
  assign data_masked[2453] = data_i[2453] & sel_one_hot_i[4];
  assign data_masked[2452] = data_i[2452] & sel_one_hot_i[4];
  assign data_masked[2451] = data_i[2451] & sel_one_hot_i[4];
  assign data_masked[2450] = data_i[2450] & sel_one_hot_i[4];
  assign data_masked[2449] = data_i[2449] & sel_one_hot_i[4];
  assign data_masked[2448] = data_i[2448] & sel_one_hot_i[4];
  assign data_masked[2447] = data_i[2447] & sel_one_hot_i[4];
  assign data_masked[2446] = data_i[2446] & sel_one_hot_i[4];
  assign data_masked[2445] = data_i[2445] & sel_one_hot_i[4];
  assign data_masked[2444] = data_i[2444] & sel_one_hot_i[4];
  assign data_masked[2443] = data_i[2443] & sel_one_hot_i[4];
  assign data_masked[2442] = data_i[2442] & sel_one_hot_i[4];
  assign data_masked[2441] = data_i[2441] & sel_one_hot_i[4];
  assign data_masked[2440] = data_i[2440] & sel_one_hot_i[4];
  assign data_masked[2439] = data_i[2439] & sel_one_hot_i[4];
  assign data_masked[2438] = data_i[2438] & sel_one_hot_i[4];
  assign data_masked[2437] = data_i[2437] & sel_one_hot_i[4];
  assign data_masked[2436] = data_i[2436] & sel_one_hot_i[4];
  assign data_masked[2435] = data_i[2435] & sel_one_hot_i[4];
  assign data_masked[2434] = data_i[2434] & sel_one_hot_i[4];
  assign data_masked[2433] = data_i[2433] & sel_one_hot_i[4];
  assign data_masked[2432] = data_i[2432] & sel_one_hot_i[4];
  assign data_masked[2431] = data_i[2431] & sel_one_hot_i[4];
  assign data_masked[2430] = data_i[2430] & sel_one_hot_i[4];
  assign data_masked[2429] = data_i[2429] & sel_one_hot_i[4];
  assign data_masked[2428] = data_i[2428] & sel_one_hot_i[4];
  assign data_masked[2427] = data_i[2427] & sel_one_hot_i[4];
  assign data_masked[2426] = data_i[2426] & sel_one_hot_i[4];
  assign data_masked[2425] = data_i[2425] & sel_one_hot_i[4];
  assign data_masked[2424] = data_i[2424] & sel_one_hot_i[4];
  assign data_masked[2423] = data_i[2423] & sel_one_hot_i[4];
  assign data_masked[2422] = data_i[2422] & sel_one_hot_i[4];
  assign data_masked[2421] = data_i[2421] & sel_one_hot_i[4];
  assign data_masked[2420] = data_i[2420] & sel_one_hot_i[4];
  assign data_masked[2419] = data_i[2419] & sel_one_hot_i[4];
  assign data_masked[2418] = data_i[2418] & sel_one_hot_i[4];
  assign data_masked[2417] = data_i[2417] & sel_one_hot_i[4];
  assign data_masked[2416] = data_i[2416] & sel_one_hot_i[4];
  assign data_masked[2415] = data_i[2415] & sel_one_hot_i[4];
  assign data_masked[2414] = data_i[2414] & sel_one_hot_i[4];
  assign data_masked[2413] = data_i[2413] & sel_one_hot_i[4];
  assign data_masked[2412] = data_i[2412] & sel_one_hot_i[4];
  assign data_masked[2411] = data_i[2411] & sel_one_hot_i[4];
  assign data_masked[2410] = data_i[2410] & sel_one_hot_i[4];
  assign data_masked[2409] = data_i[2409] & sel_one_hot_i[4];
  assign data_masked[2408] = data_i[2408] & sel_one_hot_i[4];
  assign data_masked[2407] = data_i[2407] & sel_one_hot_i[4];
  assign data_masked[2406] = data_i[2406] & sel_one_hot_i[4];
  assign data_masked[2405] = data_i[2405] & sel_one_hot_i[4];
  assign data_masked[2404] = data_i[2404] & sel_one_hot_i[4];
  assign data_masked[2403] = data_i[2403] & sel_one_hot_i[4];
  assign data_masked[2402] = data_i[2402] & sel_one_hot_i[4];
  assign data_masked[2401] = data_i[2401] & sel_one_hot_i[4];
  assign data_masked[2400] = data_i[2400] & sel_one_hot_i[4];
  assign data_masked[2399] = data_i[2399] & sel_one_hot_i[4];
  assign data_masked[2398] = data_i[2398] & sel_one_hot_i[4];
  assign data_masked[2397] = data_i[2397] & sel_one_hot_i[4];
  assign data_masked[2396] = data_i[2396] & sel_one_hot_i[4];
  assign data_masked[2395] = data_i[2395] & sel_one_hot_i[4];
  assign data_masked[2394] = data_i[2394] & sel_one_hot_i[4];
  assign data_masked[2393] = data_i[2393] & sel_one_hot_i[4];
  assign data_masked[2392] = data_i[2392] & sel_one_hot_i[4];
  assign data_masked[2391] = data_i[2391] & sel_one_hot_i[4];
  assign data_masked[2390] = data_i[2390] & sel_one_hot_i[4];
  assign data_masked[2389] = data_i[2389] & sel_one_hot_i[4];
  assign data_masked[2388] = data_i[2388] & sel_one_hot_i[4];
  assign data_masked[2387] = data_i[2387] & sel_one_hot_i[4];
  assign data_masked[2386] = data_i[2386] & sel_one_hot_i[4];
  assign data_masked[2385] = data_i[2385] & sel_one_hot_i[4];
  assign data_masked[2384] = data_i[2384] & sel_one_hot_i[4];
  assign data_masked[2383] = data_i[2383] & sel_one_hot_i[4];
  assign data_masked[2382] = data_i[2382] & sel_one_hot_i[4];
  assign data_masked[2381] = data_i[2381] & sel_one_hot_i[4];
  assign data_masked[2380] = data_i[2380] & sel_one_hot_i[4];
  assign data_masked[2379] = data_i[2379] & sel_one_hot_i[4];
  assign data_masked[2378] = data_i[2378] & sel_one_hot_i[4];
  assign data_masked[2377] = data_i[2377] & sel_one_hot_i[4];
  assign data_masked[2376] = data_i[2376] & sel_one_hot_i[4];
  assign data_masked[2375] = data_i[2375] & sel_one_hot_i[4];
  assign data_masked[2374] = data_i[2374] & sel_one_hot_i[4];
  assign data_masked[2373] = data_i[2373] & sel_one_hot_i[4];
  assign data_masked[2372] = data_i[2372] & sel_one_hot_i[4];
  assign data_masked[2371] = data_i[2371] & sel_one_hot_i[4];
  assign data_masked[2370] = data_i[2370] & sel_one_hot_i[4];
  assign data_masked[2369] = data_i[2369] & sel_one_hot_i[4];
  assign data_masked[2368] = data_i[2368] & sel_one_hot_i[4];
  assign data_masked[2367] = data_i[2367] & sel_one_hot_i[4];
  assign data_masked[2366] = data_i[2366] & sel_one_hot_i[4];
  assign data_masked[2365] = data_i[2365] & sel_one_hot_i[4];
  assign data_masked[2364] = data_i[2364] & sel_one_hot_i[4];
  assign data_masked[2363] = data_i[2363] & sel_one_hot_i[4];
  assign data_masked[2362] = data_i[2362] & sel_one_hot_i[4];
  assign data_masked[2361] = data_i[2361] & sel_one_hot_i[4];
  assign data_masked[2360] = data_i[2360] & sel_one_hot_i[4];
  assign data_masked[2359] = data_i[2359] & sel_one_hot_i[4];
  assign data_masked[2358] = data_i[2358] & sel_one_hot_i[4];
  assign data_masked[2357] = data_i[2357] & sel_one_hot_i[4];
  assign data_masked[2356] = data_i[2356] & sel_one_hot_i[4];
  assign data_masked[2355] = data_i[2355] & sel_one_hot_i[4];
  assign data_masked[2354] = data_i[2354] & sel_one_hot_i[4];
  assign data_masked[2353] = data_i[2353] & sel_one_hot_i[4];
  assign data_masked[2352] = data_i[2352] & sel_one_hot_i[4];
  assign data_masked[2351] = data_i[2351] & sel_one_hot_i[4];
  assign data_masked[2350] = data_i[2350] & sel_one_hot_i[4];
  assign data_masked[2349] = data_i[2349] & sel_one_hot_i[4];
  assign data_masked[2348] = data_i[2348] & sel_one_hot_i[4];
  assign data_masked[2347] = data_i[2347] & sel_one_hot_i[4];
  assign data_masked[2346] = data_i[2346] & sel_one_hot_i[4];
  assign data_masked[2345] = data_i[2345] & sel_one_hot_i[4];
  assign data_masked[2344] = data_i[2344] & sel_one_hot_i[4];
  assign data_masked[2343] = data_i[2343] & sel_one_hot_i[4];
  assign data_masked[2342] = data_i[2342] & sel_one_hot_i[4];
  assign data_masked[2341] = data_i[2341] & sel_one_hot_i[4];
  assign data_masked[2340] = data_i[2340] & sel_one_hot_i[4];
  assign data_masked[2339] = data_i[2339] & sel_one_hot_i[4];
  assign data_masked[2338] = data_i[2338] & sel_one_hot_i[4];
  assign data_masked[2337] = data_i[2337] & sel_one_hot_i[4];
  assign data_masked[2336] = data_i[2336] & sel_one_hot_i[4];
  assign data_masked[2335] = data_i[2335] & sel_one_hot_i[4];
  assign data_masked[2334] = data_i[2334] & sel_one_hot_i[4];
  assign data_masked[2333] = data_i[2333] & sel_one_hot_i[4];
  assign data_masked[2332] = data_i[2332] & sel_one_hot_i[4];
  assign data_masked[2331] = data_i[2331] & sel_one_hot_i[4];
  assign data_masked[2330] = data_i[2330] & sel_one_hot_i[4];
  assign data_masked[2329] = data_i[2329] & sel_one_hot_i[4];
  assign data_masked[2328] = data_i[2328] & sel_one_hot_i[4];
  assign data_masked[2327] = data_i[2327] & sel_one_hot_i[4];
  assign data_masked[2326] = data_i[2326] & sel_one_hot_i[4];
  assign data_masked[2325] = data_i[2325] & sel_one_hot_i[4];
  assign data_masked[2324] = data_i[2324] & sel_one_hot_i[4];
  assign data_masked[2323] = data_i[2323] & sel_one_hot_i[4];
  assign data_masked[2322] = data_i[2322] & sel_one_hot_i[4];
  assign data_masked[2321] = data_i[2321] & sel_one_hot_i[4];
  assign data_masked[2320] = data_i[2320] & sel_one_hot_i[4];
  assign data_masked[2319] = data_i[2319] & sel_one_hot_i[4];
  assign data_masked[2318] = data_i[2318] & sel_one_hot_i[4];
  assign data_masked[2317] = data_i[2317] & sel_one_hot_i[4];
  assign data_masked[2316] = data_i[2316] & sel_one_hot_i[4];
  assign data_masked[2315] = data_i[2315] & sel_one_hot_i[4];
  assign data_masked[2314] = data_i[2314] & sel_one_hot_i[4];
  assign data_masked[2313] = data_i[2313] & sel_one_hot_i[4];
  assign data_masked[2312] = data_i[2312] & sel_one_hot_i[4];
  assign data_masked[2311] = data_i[2311] & sel_one_hot_i[4];
  assign data_masked[2310] = data_i[2310] & sel_one_hot_i[4];
  assign data_masked[2309] = data_i[2309] & sel_one_hot_i[4];
  assign data_masked[2308] = data_i[2308] & sel_one_hot_i[4];
  assign data_masked[2307] = data_i[2307] & sel_one_hot_i[4];
  assign data_masked[2306] = data_i[2306] & sel_one_hot_i[4];
  assign data_masked[2305] = data_i[2305] & sel_one_hot_i[4];
  assign data_masked[2304] = data_i[2304] & sel_one_hot_i[4];
  assign data_masked[2303] = data_i[2303] & sel_one_hot_i[4];
  assign data_masked[2302] = data_i[2302] & sel_one_hot_i[4];
  assign data_masked[2301] = data_i[2301] & sel_one_hot_i[4];
  assign data_masked[2300] = data_i[2300] & sel_one_hot_i[4];
  assign data_masked[2299] = data_i[2299] & sel_one_hot_i[4];
  assign data_masked[2298] = data_i[2298] & sel_one_hot_i[4];
  assign data_masked[2297] = data_i[2297] & sel_one_hot_i[4];
  assign data_masked[2296] = data_i[2296] & sel_one_hot_i[4];
  assign data_masked[2295] = data_i[2295] & sel_one_hot_i[4];
  assign data_masked[2294] = data_i[2294] & sel_one_hot_i[4];
  assign data_masked[2293] = data_i[2293] & sel_one_hot_i[4];
  assign data_masked[2292] = data_i[2292] & sel_one_hot_i[4];
  assign data_masked[2291] = data_i[2291] & sel_one_hot_i[4];
  assign data_masked[2290] = data_i[2290] & sel_one_hot_i[4];
  assign data_masked[2289] = data_i[2289] & sel_one_hot_i[4];
  assign data_masked[2288] = data_i[2288] & sel_one_hot_i[4];
  assign data_masked[2287] = data_i[2287] & sel_one_hot_i[4];
  assign data_masked[2286] = data_i[2286] & sel_one_hot_i[4];
  assign data_masked[2285] = data_i[2285] & sel_one_hot_i[4];
  assign data_masked[2284] = data_i[2284] & sel_one_hot_i[4];
  assign data_masked[2283] = data_i[2283] & sel_one_hot_i[4];
  assign data_masked[2282] = data_i[2282] & sel_one_hot_i[4];
  assign data_masked[2281] = data_i[2281] & sel_one_hot_i[4];
  assign data_masked[2280] = data_i[2280] & sel_one_hot_i[4];
  assign data_masked[2279] = data_i[2279] & sel_one_hot_i[4];
  assign data_masked[2278] = data_i[2278] & sel_one_hot_i[4];
  assign data_masked[2277] = data_i[2277] & sel_one_hot_i[4];
  assign data_masked[2276] = data_i[2276] & sel_one_hot_i[4];
  assign data_masked[2275] = data_i[2275] & sel_one_hot_i[4];
  assign data_masked[2274] = data_i[2274] & sel_one_hot_i[4];
  assign data_masked[2273] = data_i[2273] & sel_one_hot_i[4];
  assign data_masked[2272] = data_i[2272] & sel_one_hot_i[4];
  assign data_masked[2271] = data_i[2271] & sel_one_hot_i[4];
  assign data_masked[2270] = data_i[2270] & sel_one_hot_i[4];
  assign data_masked[2269] = data_i[2269] & sel_one_hot_i[4];
  assign data_masked[2268] = data_i[2268] & sel_one_hot_i[4];
  assign data_masked[2267] = data_i[2267] & sel_one_hot_i[4];
  assign data_masked[2266] = data_i[2266] & sel_one_hot_i[4];
  assign data_masked[2265] = data_i[2265] & sel_one_hot_i[4];
  assign data_masked[2264] = data_i[2264] & sel_one_hot_i[4];
  assign data_masked[2263] = data_i[2263] & sel_one_hot_i[4];
  assign data_masked[2262] = data_i[2262] & sel_one_hot_i[4];
  assign data_masked[2261] = data_i[2261] & sel_one_hot_i[4];
  assign data_masked[2260] = data_i[2260] & sel_one_hot_i[4];
  assign data_masked[2259] = data_i[2259] & sel_one_hot_i[4];
  assign data_masked[2258] = data_i[2258] & sel_one_hot_i[4];
  assign data_masked[2257] = data_i[2257] & sel_one_hot_i[4];
  assign data_masked[2256] = data_i[2256] & sel_one_hot_i[4];
  assign data_masked[2255] = data_i[2255] & sel_one_hot_i[4];
  assign data_masked[2254] = data_i[2254] & sel_one_hot_i[4];
  assign data_masked[2253] = data_i[2253] & sel_one_hot_i[4];
  assign data_masked[2252] = data_i[2252] & sel_one_hot_i[4];
  assign data_masked[2251] = data_i[2251] & sel_one_hot_i[4];
  assign data_masked[2250] = data_i[2250] & sel_one_hot_i[4];
  assign data_masked[2249] = data_i[2249] & sel_one_hot_i[4];
  assign data_masked[2248] = data_i[2248] & sel_one_hot_i[4];
  assign data_masked[2247] = data_i[2247] & sel_one_hot_i[4];
  assign data_masked[2246] = data_i[2246] & sel_one_hot_i[4];
  assign data_masked[2245] = data_i[2245] & sel_one_hot_i[4];
  assign data_masked[2244] = data_i[2244] & sel_one_hot_i[4];
  assign data_masked[2243] = data_i[2243] & sel_one_hot_i[4];
  assign data_masked[2242] = data_i[2242] & sel_one_hot_i[4];
  assign data_masked[2241] = data_i[2241] & sel_one_hot_i[4];
  assign data_masked[2240] = data_i[2240] & sel_one_hot_i[4];
  assign data_masked[2239] = data_i[2239] & sel_one_hot_i[4];
  assign data_masked[2238] = data_i[2238] & sel_one_hot_i[4];
  assign data_masked[2237] = data_i[2237] & sel_one_hot_i[4];
  assign data_masked[2236] = data_i[2236] & sel_one_hot_i[4];
  assign data_masked[2235] = data_i[2235] & sel_one_hot_i[4];
  assign data_masked[2234] = data_i[2234] & sel_one_hot_i[4];
  assign data_masked[2233] = data_i[2233] & sel_one_hot_i[4];
  assign data_masked[2232] = data_i[2232] & sel_one_hot_i[4];
  assign data_masked[2231] = data_i[2231] & sel_one_hot_i[4];
  assign data_masked[2230] = data_i[2230] & sel_one_hot_i[4];
  assign data_masked[2229] = data_i[2229] & sel_one_hot_i[4];
  assign data_masked[2228] = data_i[2228] & sel_one_hot_i[4];
  assign data_masked[2227] = data_i[2227] & sel_one_hot_i[4];
  assign data_masked[2226] = data_i[2226] & sel_one_hot_i[4];
  assign data_masked[2225] = data_i[2225] & sel_one_hot_i[4];
  assign data_masked[2224] = data_i[2224] & sel_one_hot_i[4];
  assign data_masked[2223] = data_i[2223] & sel_one_hot_i[4];
  assign data_masked[2222] = data_i[2222] & sel_one_hot_i[4];
  assign data_masked[2221] = data_i[2221] & sel_one_hot_i[4];
  assign data_masked[2220] = data_i[2220] & sel_one_hot_i[4];
  assign data_masked[2219] = data_i[2219] & sel_one_hot_i[4];
  assign data_masked[2218] = data_i[2218] & sel_one_hot_i[4];
  assign data_masked[2217] = data_i[2217] & sel_one_hot_i[4];
  assign data_masked[2216] = data_i[2216] & sel_one_hot_i[4];
  assign data_masked[2215] = data_i[2215] & sel_one_hot_i[4];
  assign data_masked[2214] = data_i[2214] & sel_one_hot_i[4];
  assign data_masked[2213] = data_i[2213] & sel_one_hot_i[4];
  assign data_masked[2212] = data_i[2212] & sel_one_hot_i[4];
  assign data_masked[2211] = data_i[2211] & sel_one_hot_i[4];
  assign data_masked[2210] = data_i[2210] & sel_one_hot_i[4];
  assign data_masked[2209] = data_i[2209] & sel_one_hot_i[4];
  assign data_masked[2208] = data_i[2208] & sel_one_hot_i[4];
  assign data_masked[2207] = data_i[2207] & sel_one_hot_i[4];
  assign data_masked[2206] = data_i[2206] & sel_one_hot_i[4];
  assign data_masked[2205] = data_i[2205] & sel_one_hot_i[4];
  assign data_masked[2204] = data_i[2204] & sel_one_hot_i[4];
  assign data_masked[2203] = data_i[2203] & sel_one_hot_i[4];
  assign data_masked[2202] = data_i[2202] & sel_one_hot_i[4];
  assign data_masked[2201] = data_i[2201] & sel_one_hot_i[4];
  assign data_masked[2200] = data_i[2200] & sel_one_hot_i[4];
  assign data_masked[2199] = data_i[2199] & sel_one_hot_i[4];
  assign data_masked[2198] = data_i[2198] & sel_one_hot_i[4];
  assign data_masked[2197] = data_i[2197] & sel_one_hot_i[4];
  assign data_masked[2196] = data_i[2196] & sel_one_hot_i[4];
  assign data_masked[2195] = data_i[2195] & sel_one_hot_i[4];
  assign data_masked[2194] = data_i[2194] & sel_one_hot_i[4];
  assign data_masked[2193] = data_i[2193] & sel_one_hot_i[4];
  assign data_masked[2192] = data_i[2192] & sel_one_hot_i[4];
  assign data_masked[2191] = data_i[2191] & sel_one_hot_i[4];
  assign data_masked[2190] = data_i[2190] & sel_one_hot_i[4];
  assign data_masked[2189] = data_i[2189] & sel_one_hot_i[4];
  assign data_masked[2188] = data_i[2188] & sel_one_hot_i[4];
  assign data_masked[2187] = data_i[2187] & sel_one_hot_i[4];
  assign data_masked[2186] = data_i[2186] & sel_one_hot_i[4];
  assign data_masked[2185] = data_i[2185] & sel_one_hot_i[4];
  assign data_masked[2184] = data_i[2184] & sel_one_hot_i[4];
  assign data_masked[2183] = data_i[2183] & sel_one_hot_i[4];
  assign data_masked[2182] = data_i[2182] & sel_one_hot_i[4];
  assign data_masked[2181] = data_i[2181] & sel_one_hot_i[4];
  assign data_masked[2180] = data_i[2180] & sel_one_hot_i[4];
  assign data_masked[2179] = data_i[2179] & sel_one_hot_i[4];
  assign data_masked[2178] = data_i[2178] & sel_one_hot_i[4];
  assign data_masked[2177] = data_i[2177] & sel_one_hot_i[4];
  assign data_masked[2176] = data_i[2176] & sel_one_hot_i[4];
  assign data_masked[2175] = data_i[2175] & sel_one_hot_i[4];
  assign data_masked[2174] = data_i[2174] & sel_one_hot_i[4];
  assign data_masked[2173] = data_i[2173] & sel_one_hot_i[4];
  assign data_masked[2172] = data_i[2172] & sel_one_hot_i[4];
  assign data_masked[2171] = data_i[2171] & sel_one_hot_i[4];
  assign data_masked[2170] = data_i[2170] & sel_one_hot_i[4];
  assign data_masked[2169] = data_i[2169] & sel_one_hot_i[4];
  assign data_masked[2168] = data_i[2168] & sel_one_hot_i[4];
  assign data_masked[2167] = data_i[2167] & sel_one_hot_i[4];
  assign data_masked[2166] = data_i[2166] & sel_one_hot_i[4];
  assign data_masked[2165] = data_i[2165] & sel_one_hot_i[4];
  assign data_masked[2164] = data_i[2164] & sel_one_hot_i[4];
  assign data_masked[2163] = data_i[2163] & sel_one_hot_i[4];
  assign data_masked[2162] = data_i[2162] & sel_one_hot_i[4];
  assign data_masked[2161] = data_i[2161] & sel_one_hot_i[4];
  assign data_masked[2160] = data_i[2160] & sel_one_hot_i[4];
  assign data_masked[2159] = data_i[2159] & sel_one_hot_i[4];
  assign data_masked[2158] = data_i[2158] & sel_one_hot_i[4];
  assign data_masked[2157] = data_i[2157] & sel_one_hot_i[4];
  assign data_masked[2156] = data_i[2156] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[539];
  assign N1 = N0 | data_masked[1078];
  assign N0 = data_masked[2156] | data_masked[1617];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[540];
  assign N4 = N3 | data_masked[1079];
  assign N3 = data_masked[2157] | data_masked[1618];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[541];
  assign N7 = N6 | data_masked[1080];
  assign N6 = data_masked[2158] | data_masked[1619];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[542];
  assign N10 = N9 | data_masked[1081];
  assign N9 = data_masked[2159] | data_masked[1620];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[543];
  assign N13 = N12 | data_masked[1082];
  assign N12 = data_masked[2160] | data_masked[1621];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[544];
  assign N16 = N15 | data_masked[1083];
  assign N15 = data_masked[2161] | data_masked[1622];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[545];
  assign N19 = N18 | data_masked[1084];
  assign N18 = data_masked[2162] | data_masked[1623];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[546];
  assign N22 = N21 | data_masked[1085];
  assign N21 = data_masked[2163] | data_masked[1624];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[547];
  assign N25 = N24 | data_masked[1086];
  assign N24 = data_masked[2164] | data_masked[1625];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[548];
  assign N28 = N27 | data_masked[1087];
  assign N27 = data_masked[2165] | data_masked[1626];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[549];
  assign N31 = N30 | data_masked[1088];
  assign N30 = data_masked[2166] | data_masked[1627];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[550];
  assign N34 = N33 | data_masked[1089];
  assign N33 = data_masked[2167] | data_masked[1628];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[551];
  assign N37 = N36 | data_masked[1090];
  assign N36 = data_masked[2168] | data_masked[1629];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[552];
  assign N40 = N39 | data_masked[1091];
  assign N39 = data_masked[2169] | data_masked[1630];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[553];
  assign N43 = N42 | data_masked[1092];
  assign N42 = data_masked[2170] | data_masked[1631];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[554];
  assign N46 = N45 | data_masked[1093];
  assign N45 = data_masked[2171] | data_masked[1632];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[555];
  assign N49 = N48 | data_masked[1094];
  assign N48 = data_masked[2172] | data_masked[1633];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[556];
  assign N52 = N51 | data_masked[1095];
  assign N51 = data_masked[2173] | data_masked[1634];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[557];
  assign N55 = N54 | data_masked[1096];
  assign N54 = data_masked[2174] | data_masked[1635];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[558];
  assign N58 = N57 | data_masked[1097];
  assign N57 = data_masked[2175] | data_masked[1636];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[559];
  assign N61 = N60 | data_masked[1098];
  assign N60 = data_masked[2176] | data_masked[1637];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[560];
  assign N64 = N63 | data_masked[1099];
  assign N63 = data_masked[2177] | data_masked[1638];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[561];
  assign N67 = N66 | data_masked[1100];
  assign N66 = data_masked[2178] | data_masked[1639];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[562];
  assign N70 = N69 | data_masked[1101];
  assign N69 = data_masked[2179] | data_masked[1640];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[563];
  assign N73 = N72 | data_masked[1102];
  assign N72 = data_masked[2180] | data_masked[1641];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[564];
  assign N76 = N75 | data_masked[1103];
  assign N75 = data_masked[2181] | data_masked[1642];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[565];
  assign N79 = N78 | data_masked[1104];
  assign N78 = data_masked[2182] | data_masked[1643];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[566];
  assign N82 = N81 | data_masked[1105];
  assign N81 = data_masked[2183] | data_masked[1644];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[567];
  assign N85 = N84 | data_masked[1106];
  assign N84 = data_masked[2184] | data_masked[1645];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[568];
  assign N88 = N87 | data_masked[1107];
  assign N87 = data_masked[2185] | data_masked[1646];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[569];
  assign N91 = N90 | data_masked[1108];
  assign N90 = data_masked[2186] | data_masked[1647];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[570];
  assign N94 = N93 | data_masked[1109];
  assign N93 = data_masked[2187] | data_masked[1648];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[571];
  assign N97 = N96 | data_masked[1110];
  assign N96 = data_masked[2188] | data_masked[1649];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[572];
  assign N100 = N99 | data_masked[1111];
  assign N99 = data_masked[2189] | data_masked[1650];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[573];
  assign N103 = N102 | data_masked[1112];
  assign N102 = data_masked[2190] | data_masked[1651];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[574];
  assign N106 = N105 | data_masked[1113];
  assign N105 = data_masked[2191] | data_masked[1652];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[575];
  assign N109 = N108 | data_masked[1114];
  assign N108 = data_masked[2192] | data_masked[1653];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[576];
  assign N112 = N111 | data_masked[1115];
  assign N111 = data_masked[2193] | data_masked[1654];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[577];
  assign N115 = N114 | data_masked[1116];
  assign N114 = data_masked[2194] | data_masked[1655];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[578];
  assign N118 = N117 | data_masked[1117];
  assign N117 = data_masked[2195] | data_masked[1656];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[579];
  assign N121 = N120 | data_masked[1118];
  assign N120 = data_masked[2196] | data_masked[1657];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[580];
  assign N124 = N123 | data_masked[1119];
  assign N123 = data_masked[2197] | data_masked[1658];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[581];
  assign N127 = N126 | data_masked[1120];
  assign N126 = data_masked[2198] | data_masked[1659];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[582];
  assign N130 = N129 | data_masked[1121];
  assign N129 = data_masked[2199] | data_masked[1660];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[583];
  assign N133 = N132 | data_masked[1122];
  assign N132 = data_masked[2200] | data_masked[1661];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[584];
  assign N136 = N135 | data_masked[1123];
  assign N135 = data_masked[2201] | data_masked[1662];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[585];
  assign N139 = N138 | data_masked[1124];
  assign N138 = data_masked[2202] | data_masked[1663];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[586];
  assign N142 = N141 | data_masked[1125];
  assign N141 = data_masked[2203] | data_masked[1664];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[587];
  assign N145 = N144 | data_masked[1126];
  assign N144 = data_masked[2204] | data_masked[1665];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[588];
  assign N148 = N147 | data_masked[1127];
  assign N147 = data_masked[2205] | data_masked[1666];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[589];
  assign N151 = N150 | data_masked[1128];
  assign N150 = data_masked[2206] | data_masked[1667];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[590];
  assign N154 = N153 | data_masked[1129];
  assign N153 = data_masked[2207] | data_masked[1668];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[591];
  assign N157 = N156 | data_masked[1130];
  assign N156 = data_masked[2208] | data_masked[1669];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[592];
  assign N160 = N159 | data_masked[1131];
  assign N159 = data_masked[2209] | data_masked[1670];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[593];
  assign N163 = N162 | data_masked[1132];
  assign N162 = data_masked[2210] | data_masked[1671];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[594];
  assign N166 = N165 | data_masked[1133];
  assign N165 = data_masked[2211] | data_masked[1672];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[595];
  assign N169 = N168 | data_masked[1134];
  assign N168 = data_masked[2212] | data_masked[1673];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[596];
  assign N172 = N171 | data_masked[1135];
  assign N171 = data_masked[2213] | data_masked[1674];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[597];
  assign N175 = N174 | data_masked[1136];
  assign N174 = data_masked[2214] | data_masked[1675];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[598];
  assign N178 = N177 | data_masked[1137];
  assign N177 = data_masked[2215] | data_masked[1676];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[599];
  assign N181 = N180 | data_masked[1138];
  assign N180 = data_masked[2216] | data_masked[1677];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[600];
  assign N184 = N183 | data_masked[1139];
  assign N183 = data_masked[2217] | data_masked[1678];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[601];
  assign N187 = N186 | data_masked[1140];
  assign N186 = data_masked[2218] | data_masked[1679];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[602];
  assign N190 = N189 | data_masked[1141];
  assign N189 = data_masked[2219] | data_masked[1680];
  assign data_o[64] = N194 | data_masked[64];
  assign N194 = N193 | data_masked[603];
  assign N193 = N192 | data_masked[1142];
  assign N192 = data_masked[2220] | data_masked[1681];
  assign data_o[65] = N197 | data_masked[65];
  assign N197 = N196 | data_masked[604];
  assign N196 = N195 | data_masked[1143];
  assign N195 = data_masked[2221] | data_masked[1682];
  assign data_o[66] = N200 | data_masked[66];
  assign N200 = N199 | data_masked[605];
  assign N199 = N198 | data_masked[1144];
  assign N198 = data_masked[2222] | data_masked[1683];
  assign data_o[67] = N203 | data_masked[67];
  assign N203 = N202 | data_masked[606];
  assign N202 = N201 | data_masked[1145];
  assign N201 = data_masked[2223] | data_masked[1684];
  assign data_o[68] = N206 | data_masked[68];
  assign N206 = N205 | data_masked[607];
  assign N205 = N204 | data_masked[1146];
  assign N204 = data_masked[2224] | data_masked[1685];
  assign data_o[69] = N209 | data_masked[69];
  assign N209 = N208 | data_masked[608];
  assign N208 = N207 | data_masked[1147];
  assign N207 = data_masked[2225] | data_masked[1686];
  assign data_o[70] = N212 | data_masked[70];
  assign N212 = N211 | data_masked[609];
  assign N211 = N210 | data_masked[1148];
  assign N210 = data_masked[2226] | data_masked[1687];
  assign data_o[71] = N215 | data_masked[71];
  assign N215 = N214 | data_masked[610];
  assign N214 = N213 | data_masked[1149];
  assign N213 = data_masked[2227] | data_masked[1688];
  assign data_o[72] = N218 | data_masked[72];
  assign N218 = N217 | data_masked[611];
  assign N217 = N216 | data_masked[1150];
  assign N216 = data_masked[2228] | data_masked[1689];
  assign data_o[73] = N221 | data_masked[73];
  assign N221 = N220 | data_masked[612];
  assign N220 = N219 | data_masked[1151];
  assign N219 = data_masked[2229] | data_masked[1690];
  assign data_o[74] = N224 | data_masked[74];
  assign N224 = N223 | data_masked[613];
  assign N223 = N222 | data_masked[1152];
  assign N222 = data_masked[2230] | data_masked[1691];
  assign data_o[75] = N227 | data_masked[75];
  assign N227 = N226 | data_masked[614];
  assign N226 = N225 | data_masked[1153];
  assign N225 = data_masked[2231] | data_masked[1692];
  assign data_o[76] = N230 | data_masked[76];
  assign N230 = N229 | data_masked[615];
  assign N229 = N228 | data_masked[1154];
  assign N228 = data_masked[2232] | data_masked[1693];
  assign data_o[77] = N233 | data_masked[77];
  assign N233 = N232 | data_masked[616];
  assign N232 = N231 | data_masked[1155];
  assign N231 = data_masked[2233] | data_masked[1694];
  assign data_o[78] = N236 | data_masked[78];
  assign N236 = N235 | data_masked[617];
  assign N235 = N234 | data_masked[1156];
  assign N234 = data_masked[2234] | data_masked[1695];
  assign data_o[79] = N239 | data_masked[79];
  assign N239 = N238 | data_masked[618];
  assign N238 = N237 | data_masked[1157];
  assign N237 = data_masked[2235] | data_masked[1696];
  assign data_o[80] = N242 | data_masked[80];
  assign N242 = N241 | data_masked[619];
  assign N241 = N240 | data_masked[1158];
  assign N240 = data_masked[2236] | data_masked[1697];
  assign data_o[81] = N245 | data_masked[81];
  assign N245 = N244 | data_masked[620];
  assign N244 = N243 | data_masked[1159];
  assign N243 = data_masked[2237] | data_masked[1698];
  assign data_o[82] = N248 | data_masked[82];
  assign N248 = N247 | data_masked[621];
  assign N247 = N246 | data_masked[1160];
  assign N246 = data_masked[2238] | data_masked[1699];
  assign data_o[83] = N251 | data_masked[83];
  assign N251 = N250 | data_masked[622];
  assign N250 = N249 | data_masked[1161];
  assign N249 = data_masked[2239] | data_masked[1700];
  assign data_o[84] = N254 | data_masked[84];
  assign N254 = N253 | data_masked[623];
  assign N253 = N252 | data_masked[1162];
  assign N252 = data_masked[2240] | data_masked[1701];
  assign data_o[85] = N257 | data_masked[85];
  assign N257 = N256 | data_masked[624];
  assign N256 = N255 | data_masked[1163];
  assign N255 = data_masked[2241] | data_masked[1702];
  assign data_o[86] = N260 | data_masked[86];
  assign N260 = N259 | data_masked[625];
  assign N259 = N258 | data_masked[1164];
  assign N258 = data_masked[2242] | data_masked[1703];
  assign data_o[87] = N263 | data_masked[87];
  assign N263 = N262 | data_masked[626];
  assign N262 = N261 | data_masked[1165];
  assign N261 = data_masked[2243] | data_masked[1704];
  assign data_o[88] = N266 | data_masked[88];
  assign N266 = N265 | data_masked[627];
  assign N265 = N264 | data_masked[1166];
  assign N264 = data_masked[2244] | data_masked[1705];
  assign data_o[89] = N269 | data_masked[89];
  assign N269 = N268 | data_masked[628];
  assign N268 = N267 | data_masked[1167];
  assign N267 = data_masked[2245] | data_masked[1706];
  assign data_o[90] = N272 | data_masked[90];
  assign N272 = N271 | data_masked[629];
  assign N271 = N270 | data_masked[1168];
  assign N270 = data_masked[2246] | data_masked[1707];
  assign data_o[91] = N275 | data_masked[91];
  assign N275 = N274 | data_masked[630];
  assign N274 = N273 | data_masked[1169];
  assign N273 = data_masked[2247] | data_masked[1708];
  assign data_o[92] = N278 | data_masked[92];
  assign N278 = N277 | data_masked[631];
  assign N277 = N276 | data_masked[1170];
  assign N276 = data_masked[2248] | data_masked[1709];
  assign data_o[93] = N281 | data_masked[93];
  assign N281 = N280 | data_masked[632];
  assign N280 = N279 | data_masked[1171];
  assign N279 = data_masked[2249] | data_masked[1710];
  assign data_o[94] = N284 | data_masked[94];
  assign N284 = N283 | data_masked[633];
  assign N283 = N282 | data_masked[1172];
  assign N282 = data_masked[2250] | data_masked[1711];
  assign data_o[95] = N287 | data_masked[95];
  assign N287 = N286 | data_masked[634];
  assign N286 = N285 | data_masked[1173];
  assign N285 = data_masked[2251] | data_masked[1712];
  assign data_o[96] = N290 | data_masked[96];
  assign N290 = N289 | data_masked[635];
  assign N289 = N288 | data_masked[1174];
  assign N288 = data_masked[2252] | data_masked[1713];
  assign data_o[97] = N293 | data_masked[97];
  assign N293 = N292 | data_masked[636];
  assign N292 = N291 | data_masked[1175];
  assign N291 = data_masked[2253] | data_masked[1714];
  assign data_o[98] = N296 | data_masked[98];
  assign N296 = N295 | data_masked[637];
  assign N295 = N294 | data_masked[1176];
  assign N294 = data_masked[2254] | data_masked[1715];
  assign data_o[99] = N299 | data_masked[99];
  assign N299 = N298 | data_masked[638];
  assign N298 = N297 | data_masked[1177];
  assign N297 = data_masked[2255] | data_masked[1716];
  assign data_o[100] = N302 | data_masked[100];
  assign N302 = N301 | data_masked[639];
  assign N301 = N300 | data_masked[1178];
  assign N300 = data_masked[2256] | data_masked[1717];
  assign data_o[101] = N305 | data_masked[101];
  assign N305 = N304 | data_masked[640];
  assign N304 = N303 | data_masked[1179];
  assign N303 = data_masked[2257] | data_masked[1718];
  assign data_o[102] = N308 | data_masked[102];
  assign N308 = N307 | data_masked[641];
  assign N307 = N306 | data_masked[1180];
  assign N306 = data_masked[2258] | data_masked[1719];
  assign data_o[103] = N311 | data_masked[103];
  assign N311 = N310 | data_masked[642];
  assign N310 = N309 | data_masked[1181];
  assign N309 = data_masked[2259] | data_masked[1720];
  assign data_o[104] = N314 | data_masked[104];
  assign N314 = N313 | data_masked[643];
  assign N313 = N312 | data_masked[1182];
  assign N312 = data_masked[2260] | data_masked[1721];
  assign data_o[105] = N317 | data_masked[105];
  assign N317 = N316 | data_masked[644];
  assign N316 = N315 | data_masked[1183];
  assign N315 = data_masked[2261] | data_masked[1722];
  assign data_o[106] = N320 | data_masked[106];
  assign N320 = N319 | data_masked[645];
  assign N319 = N318 | data_masked[1184];
  assign N318 = data_masked[2262] | data_masked[1723];
  assign data_o[107] = N323 | data_masked[107];
  assign N323 = N322 | data_masked[646];
  assign N322 = N321 | data_masked[1185];
  assign N321 = data_masked[2263] | data_masked[1724];
  assign data_o[108] = N326 | data_masked[108];
  assign N326 = N325 | data_masked[647];
  assign N325 = N324 | data_masked[1186];
  assign N324 = data_masked[2264] | data_masked[1725];
  assign data_o[109] = N329 | data_masked[109];
  assign N329 = N328 | data_masked[648];
  assign N328 = N327 | data_masked[1187];
  assign N327 = data_masked[2265] | data_masked[1726];
  assign data_o[110] = N332 | data_masked[110];
  assign N332 = N331 | data_masked[649];
  assign N331 = N330 | data_masked[1188];
  assign N330 = data_masked[2266] | data_masked[1727];
  assign data_o[111] = N335 | data_masked[111];
  assign N335 = N334 | data_masked[650];
  assign N334 = N333 | data_masked[1189];
  assign N333 = data_masked[2267] | data_masked[1728];
  assign data_o[112] = N338 | data_masked[112];
  assign N338 = N337 | data_masked[651];
  assign N337 = N336 | data_masked[1190];
  assign N336 = data_masked[2268] | data_masked[1729];
  assign data_o[113] = N341 | data_masked[113];
  assign N341 = N340 | data_masked[652];
  assign N340 = N339 | data_masked[1191];
  assign N339 = data_masked[2269] | data_masked[1730];
  assign data_o[114] = N344 | data_masked[114];
  assign N344 = N343 | data_masked[653];
  assign N343 = N342 | data_masked[1192];
  assign N342 = data_masked[2270] | data_masked[1731];
  assign data_o[115] = N347 | data_masked[115];
  assign N347 = N346 | data_masked[654];
  assign N346 = N345 | data_masked[1193];
  assign N345 = data_masked[2271] | data_masked[1732];
  assign data_o[116] = N350 | data_masked[116];
  assign N350 = N349 | data_masked[655];
  assign N349 = N348 | data_masked[1194];
  assign N348 = data_masked[2272] | data_masked[1733];
  assign data_o[117] = N353 | data_masked[117];
  assign N353 = N352 | data_masked[656];
  assign N352 = N351 | data_masked[1195];
  assign N351 = data_masked[2273] | data_masked[1734];
  assign data_o[118] = N356 | data_masked[118];
  assign N356 = N355 | data_masked[657];
  assign N355 = N354 | data_masked[1196];
  assign N354 = data_masked[2274] | data_masked[1735];
  assign data_o[119] = N359 | data_masked[119];
  assign N359 = N358 | data_masked[658];
  assign N358 = N357 | data_masked[1197];
  assign N357 = data_masked[2275] | data_masked[1736];
  assign data_o[120] = N362 | data_masked[120];
  assign N362 = N361 | data_masked[659];
  assign N361 = N360 | data_masked[1198];
  assign N360 = data_masked[2276] | data_masked[1737];
  assign data_o[121] = N365 | data_masked[121];
  assign N365 = N364 | data_masked[660];
  assign N364 = N363 | data_masked[1199];
  assign N363 = data_masked[2277] | data_masked[1738];
  assign data_o[122] = N368 | data_masked[122];
  assign N368 = N367 | data_masked[661];
  assign N367 = N366 | data_masked[1200];
  assign N366 = data_masked[2278] | data_masked[1739];
  assign data_o[123] = N371 | data_masked[123];
  assign N371 = N370 | data_masked[662];
  assign N370 = N369 | data_masked[1201];
  assign N369 = data_masked[2279] | data_masked[1740];
  assign data_o[124] = N374 | data_masked[124];
  assign N374 = N373 | data_masked[663];
  assign N373 = N372 | data_masked[1202];
  assign N372 = data_masked[2280] | data_masked[1741];
  assign data_o[125] = N377 | data_masked[125];
  assign N377 = N376 | data_masked[664];
  assign N376 = N375 | data_masked[1203];
  assign N375 = data_masked[2281] | data_masked[1742];
  assign data_o[126] = N380 | data_masked[126];
  assign N380 = N379 | data_masked[665];
  assign N379 = N378 | data_masked[1204];
  assign N378 = data_masked[2282] | data_masked[1743];
  assign data_o[127] = N383 | data_masked[127];
  assign N383 = N382 | data_masked[666];
  assign N382 = N381 | data_masked[1205];
  assign N381 = data_masked[2283] | data_masked[1744];
  assign data_o[128] = N386 | data_masked[128];
  assign N386 = N385 | data_masked[667];
  assign N385 = N384 | data_masked[1206];
  assign N384 = data_masked[2284] | data_masked[1745];
  assign data_o[129] = N389 | data_masked[129];
  assign N389 = N388 | data_masked[668];
  assign N388 = N387 | data_masked[1207];
  assign N387 = data_masked[2285] | data_masked[1746];
  assign data_o[130] = N392 | data_masked[130];
  assign N392 = N391 | data_masked[669];
  assign N391 = N390 | data_masked[1208];
  assign N390 = data_masked[2286] | data_masked[1747];
  assign data_o[131] = N395 | data_masked[131];
  assign N395 = N394 | data_masked[670];
  assign N394 = N393 | data_masked[1209];
  assign N393 = data_masked[2287] | data_masked[1748];
  assign data_o[132] = N398 | data_masked[132];
  assign N398 = N397 | data_masked[671];
  assign N397 = N396 | data_masked[1210];
  assign N396 = data_masked[2288] | data_masked[1749];
  assign data_o[133] = N401 | data_masked[133];
  assign N401 = N400 | data_masked[672];
  assign N400 = N399 | data_masked[1211];
  assign N399 = data_masked[2289] | data_masked[1750];
  assign data_o[134] = N404 | data_masked[134];
  assign N404 = N403 | data_masked[673];
  assign N403 = N402 | data_masked[1212];
  assign N402 = data_masked[2290] | data_masked[1751];
  assign data_o[135] = N407 | data_masked[135];
  assign N407 = N406 | data_masked[674];
  assign N406 = N405 | data_masked[1213];
  assign N405 = data_masked[2291] | data_masked[1752];
  assign data_o[136] = N410 | data_masked[136];
  assign N410 = N409 | data_masked[675];
  assign N409 = N408 | data_masked[1214];
  assign N408 = data_masked[2292] | data_masked[1753];
  assign data_o[137] = N413 | data_masked[137];
  assign N413 = N412 | data_masked[676];
  assign N412 = N411 | data_masked[1215];
  assign N411 = data_masked[2293] | data_masked[1754];
  assign data_o[138] = N416 | data_masked[138];
  assign N416 = N415 | data_masked[677];
  assign N415 = N414 | data_masked[1216];
  assign N414 = data_masked[2294] | data_masked[1755];
  assign data_o[139] = N419 | data_masked[139];
  assign N419 = N418 | data_masked[678];
  assign N418 = N417 | data_masked[1217];
  assign N417 = data_masked[2295] | data_masked[1756];
  assign data_o[140] = N422 | data_masked[140];
  assign N422 = N421 | data_masked[679];
  assign N421 = N420 | data_masked[1218];
  assign N420 = data_masked[2296] | data_masked[1757];
  assign data_o[141] = N425 | data_masked[141];
  assign N425 = N424 | data_masked[680];
  assign N424 = N423 | data_masked[1219];
  assign N423 = data_masked[2297] | data_masked[1758];
  assign data_o[142] = N428 | data_masked[142];
  assign N428 = N427 | data_masked[681];
  assign N427 = N426 | data_masked[1220];
  assign N426 = data_masked[2298] | data_masked[1759];
  assign data_o[143] = N431 | data_masked[143];
  assign N431 = N430 | data_masked[682];
  assign N430 = N429 | data_masked[1221];
  assign N429 = data_masked[2299] | data_masked[1760];
  assign data_o[144] = N434 | data_masked[144];
  assign N434 = N433 | data_masked[683];
  assign N433 = N432 | data_masked[1222];
  assign N432 = data_masked[2300] | data_masked[1761];
  assign data_o[145] = N437 | data_masked[145];
  assign N437 = N436 | data_masked[684];
  assign N436 = N435 | data_masked[1223];
  assign N435 = data_masked[2301] | data_masked[1762];
  assign data_o[146] = N440 | data_masked[146];
  assign N440 = N439 | data_masked[685];
  assign N439 = N438 | data_masked[1224];
  assign N438 = data_masked[2302] | data_masked[1763];
  assign data_o[147] = N443 | data_masked[147];
  assign N443 = N442 | data_masked[686];
  assign N442 = N441 | data_masked[1225];
  assign N441 = data_masked[2303] | data_masked[1764];
  assign data_o[148] = N446 | data_masked[148];
  assign N446 = N445 | data_masked[687];
  assign N445 = N444 | data_masked[1226];
  assign N444 = data_masked[2304] | data_masked[1765];
  assign data_o[149] = N449 | data_masked[149];
  assign N449 = N448 | data_masked[688];
  assign N448 = N447 | data_masked[1227];
  assign N447 = data_masked[2305] | data_masked[1766];
  assign data_o[150] = N452 | data_masked[150];
  assign N452 = N451 | data_masked[689];
  assign N451 = N450 | data_masked[1228];
  assign N450 = data_masked[2306] | data_masked[1767];
  assign data_o[151] = N455 | data_masked[151];
  assign N455 = N454 | data_masked[690];
  assign N454 = N453 | data_masked[1229];
  assign N453 = data_masked[2307] | data_masked[1768];
  assign data_o[152] = N458 | data_masked[152];
  assign N458 = N457 | data_masked[691];
  assign N457 = N456 | data_masked[1230];
  assign N456 = data_masked[2308] | data_masked[1769];
  assign data_o[153] = N461 | data_masked[153];
  assign N461 = N460 | data_masked[692];
  assign N460 = N459 | data_masked[1231];
  assign N459 = data_masked[2309] | data_masked[1770];
  assign data_o[154] = N464 | data_masked[154];
  assign N464 = N463 | data_masked[693];
  assign N463 = N462 | data_masked[1232];
  assign N462 = data_masked[2310] | data_masked[1771];
  assign data_o[155] = N467 | data_masked[155];
  assign N467 = N466 | data_masked[694];
  assign N466 = N465 | data_masked[1233];
  assign N465 = data_masked[2311] | data_masked[1772];
  assign data_o[156] = N470 | data_masked[156];
  assign N470 = N469 | data_masked[695];
  assign N469 = N468 | data_masked[1234];
  assign N468 = data_masked[2312] | data_masked[1773];
  assign data_o[157] = N473 | data_masked[157];
  assign N473 = N472 | data_masked[696];
  assign N472 = N471 | data_masked[1235];
  assign N471 = data_masked[2313] | data_masked[1774];
  assign data_o[158] = N476 | data_masked[158];
  assign N476 = N475 | data_masked[697];
  assign N475 = N474 | data_masked[1236];
  assign N474 = data_masked[2314] | data_masked[1775];
  assign data_o[159] = N479 | data_masked[159];
  assign N479 = N478 | data_masked[698];
  assign N478 = N477 | data_masked[1237];
  assign N477 = data_masked[2315] | data_masked[1776];
  assign data_o[160] = N482 | data_masked[160];
  assign N482 = N481 | data_masked[699];
  assign N481 = N480 | data_masked[1238];
  assign N480 = data_masked[2316] | data_masked[1777];
  assign data_o[161] = N485 | data_masked[161];
  assign N485 = N484 | data_masked[700];
  assign N484 = N483 | data_masked[1239];
  assign N483 = data_masked[2317] | data_masked[1778];
  assign data_o[162] = N488 | data_masked[162];
  assign N488 = N487 | data_masked[701];
  assign N487 = N486 | data_masked[1240];
  assign N486 = data_masked[2318] | data_masked[1779];
  assign data_o[163] = N491 | data_masked[163];
  assign N491 = N490 | data_masked[702];
  assign N490 = N489 | data_masked[1241];
  assign N489 = data_masked[2319] | data_masked[1780];
  assign data_o[164] = N494 | data_masked[164];
  assign N494 = N493 | data_masked[703];
  assign N493 = N492 | data_masked[1242];
  assign N492 = data_masked[2320] | data_masked[1781];
  assign data_o[165] = N497 | data_masked[165];
  assign N497 = N496 | data_masked[704];
  assign N496 = N495 | data_masked[1243];
  assign N495 = data_masked[2321] | data_masked[1782];
  assign data_o[166] = N500 | data_masked[166];
  assign N500 = N499 | data_masked[705];
  assign N499 = N498 | data_masked[1244];
  assign N498 = data_masked[2322] | data_masked[1783];
  assign data_o[167] = N503 | data_masked[167];
  assign N503 = N502 | data_masked[706];
  assign N502 = N501 | data_masked[1245];
  assign N501 = data_masked[2323] | data_masked[1784];
  assign data_o[168] = N506 | data_masked[168];
  assign N506 = N505 | data_masked[707];
  assign N505 = N504 | data_masked[1246];
  assign N504 = data_masked[2324] | data_masked[1785];
  assign data_o[169] = N509 | data_masked[169];
  assign N509 = N508 | data_masked[708];
  assign N508 = N507 | data_masked[1247];
  assign N507 = data_masked[2325] | data_masked[1786];
  assign data_o[170] = N512 | data_masked[170];
  assign N512 = N511 | data_masked[709];
  assign N511 = N510 | data_masked[1248];
  assign N510 = data_masked[2326] | data_masked[1787];
  assign data_o[171] = N515 | data_masked[171];
  assign N515 = N514 | data_masked[710];
  assign N514 = N513 | data_masked[1249];
  assign N513 = data_masked[2327] | data_masked[1788];
  assign data_o[172] = N518 | data_masked[172];
  assign N518 = N517 | data_masked[711];
  assign N517 = N516 | data_masked[1250];
  assign N516 = data_masked[2328] | data_masked[1789];
  assign data_o[173] = N521 | data_masked[173];
  assign N521 = N520 | data_masked[712];
  assign N520 = N519 | data_masked[1251];
  assign N519 = data_masked[2329] | data_masked[1790];
  assign data_o[174] = N524 | data_masked[174];
  assign N524 = N523 | data_masked[713];
  assign N523 = N522 | data_masked[1252];
  assign N522 = data_masked[2330] | data_masked[1791];
  assign data_o[175] = N527 | data_masked[175];
  assign N527 = N526 | data_masked[714];
  assign N526 = N525 | data_masked[1253];
  assign N525 = data_masked[2331] | data_masked[1792];
  assign data_o[176] = N530 | data_masked[176];
  assign N530 = N529 | data_masked[715];
  assign N529 = N528 | data_masked[1254];
  assign N528 = data_masked[2332] | data_masked[1793];
  assign data_o[177] = N533 | data_masked[177];
  assign N533 = N532 | data_masked[716];
  assign N532 = N531 | data_masked[1255];
  assign N531 = data_masked[2333] | data_masked[1794];
  assign data_o[178] = N536 | data_masked[178];
  assign N536 = N535 | data_masked[717];
  assign N535 = N534 | data_masked[1256];
  assign N534 = data_masked[2334] | data_masked[1795];
  assign data_o[179] = N539 | data_masked[179];
  assign N539 = N538 | data_masked[718];
  assign N538 = N537 | data_masked[1257];
  assign N537 = data_masked[2335] | data_masked[1796];
  assign data_o[180] = N542 | data_masked[180];
  assign N542 = N541 | data_masked[719];
  assign N541 = N540 | data_masked[1258];
  assign N540 = data_masked[2336] | data_masked[1797];
  assign data_o[181] = N545 | data_masked[181];
  assign N545 = N544 | data_masked[720];
  assign N544 = N543 | data_masked[1259];
  assign N543 = data_masked[2337] | data_masked[1798];
  assign data_o[182] = N548 | data_masked[182];
  assign N548 = N547 | data_masked[721];
  assign N547 = N546 | data_masked[1260];
  assign N546 = data_masked[2338] | data_masked[1799];
  assign data_o[183] = N551 | data_masked[183];
  assign N551 = N550 | data_masked[722];
  assign N550 = N549 | data_masked[1261];
  assign N549 = data_masked[2339] | data_masked[1800];
  assign data_o[184] = N554 | data_masked[184];
  assign N554 = N553 | data_masked[723];
  assign N553 = N552 | data_masked[1262];
  assign N552 = data_masked[2340] | data_masked[1801];
  assign data_o[185] = N557 | data_masked[185];
  assign N557 = N556 | data_masked[724];
  assign N556 = N555 | data_masked[1263];
  assign N555 = data_masked[2341] | data_masked[1802];
  assign data_o[186] = N560 | data_masked[186];
  assign N560 = N559 | data_masked[725];
  assign N559 = N558 | data_masked[1264];
  assign N558 = data_masked[2342] | data_masked[1803];
  assign data_o[187] = N563 | data_masked[187];
  assign N563 = N562 | data_masked[726];
  assign N562 = N561 | data_masked[1265];
  assign N561 = data_masked[2343] | data_masked[1804];
  assign data_o[188] = N566 | data_masked[188];
  assign N566 = N565 | data_masked[727];
  assign N565 = N564 | data_masked[1266];
  assign N564 = data_masked[2344] | data_masked[1805];
  assign data_o[189] = N569 | data_masked[189];
  assign N569 = N568 | data_masked[728];
  assign N568 = N567 | data_masked[1267];
  assign N567 = data_masked[2345] | data_masked[1806];
  assign data_o[190] = N572 | data_masked[190];
  assign N572 = N571 | data_masked[729];
  assign N571 = N570 | data_masked[1268];
  assign N570 = data_masked[2346] | data_masked[1807];
  assign data_o[191] = N575 | data_masked[191];
  assign N575 = N574 | data_masked[730];
  assign N574 = N573 | data_masked[1269];
  assign N573 = data_masked[2347] | data_masked[1808];
  assign data_o[192] = N578 | data_masked[192];
  assign N578 = N577 | data_masked[731];
  assign N577 = N576 | data_masked[1270];
  assign N576 = data_masked[2348] | data_masked[1809];
  assign data_o[193] = N581 | data_masked[193];
  assign N581 = N580 | data_masked[732];
  assign N580 = N579 | data_masked[1271];
  assign N579 = data_masked[2349] | data_masked[1810];
  assign data_o[194] = N584 | data_masked[194];
  assign N584 = N583 | data_masked[733];
  assign N583 = N582 | data_masked[1272];
  assign N582 = data_masked[2350] | data_masked[1811];
  assign data_o[195] = N587 | data_masked[195];
  assign N587 = N586 | data_masked[734];
  assign N586 = N585 | data_masked[1273];
  assign N585 = data_masked[2351] | data_masked[1812];
  assign data_o[196] = N590 | data_masked[196];
  assign N590 = N589 | data_masked[735];
  assign N589 = N588 | data_masked[1274];
  assign N588 = data_masked[2352] | data_masked[1813];
  assign data_o[197] = N593 | data_masked[197];
  assign N593 = N592 | data_masked[736];
  assign N592 = N591 | data_masked[1275];
  assign N591 = data_masked[2353] | data_masked[1814];
  assign data_o[198] = N596 | data_masked[198];
  assign N596 = N595 | data_masked[737];
  assign N595 = N594 | data_masked[1276];
  assign N594 = data_masked[2354] | data_masked[1815];
  assign data_o[199] = N599 | data_masked[199];
  assign N599 = N598 | data_masked[738];
  assign N598 = N597 | data_masked[1277];
  assign N597 = data_masked[2355] | data_masked[1816];
  assign data_o[200] = N602 | data_masked[200];
  assign N602 = N601 | data_masked[739];
  assign N601 = N600 | data_masked[1278];
  assign N600 = data_masked[2356] | data_masked[1817];
  assign data_o[201] = N605 | data_masked[201];
  assign N605 = N604 | data_masked[740];
  assign N604 = N603 | data_masked[1279];
  assign N603 = data_masked[2357] | data_masked[1818];
  assign data_o[202] = N608 | data_masked[202];
  assign N608 = N607 | data_masked[741];
  assign N607 = N606 | data_masked[1280];
  assign N606 = data_masked[2358] | data_masked[1819];
  assign data_o[203] = N611 | data_masked[203];
  assign N611 = N610 | data_masked[742];
  assign N610 = N609 | data_masked[1281];
  assign N609 = data_masked[2359] | data_masked[1820];
  assign data_o[204] = N614 | data_masked[204];
  assign N614 = N613 | data_masked[743];
  assign N613 = N612 | data_masked[1282];
  assign N612 = data_masked[2360] | data_masked[1821];
  assign data_o[205] = N617 | data_masked[205];
  assign N617 = N616 | data_masked[744];
  assign N616 = N615 | data_masked[1283];
  assign N615 = data_masked[2361] | data_masked[1822];
  assign data_o[206] = N620 | data_masked[206];
  assign N620 = N619 | data_masked[745];
  assign N619 = N618 | data_masked[1284];
  assign N618 = data_masked[2362] | data_masked[1823];
  assign data_o[207] = N623 | data_masked[207];
  assign N623 = N622 | data_masked[746];
  assign N622 = N621 | data_masked[1285];
  assign N621 = data_masked[2363] | data_masked[1824];
  assign data_o[208] = N626 | data_masked[208];
  assign N626 = N625 | data_masked[747];
  assign N625 = N624 | data_masked[1286];
  assign N624 = data_masked[2364] | data_masked[1825];
  assign data_o[209] = N629 | data_masked[209];
  assign N629 = N628 | data_masked[748];
  assign N628 = N627 | data_masked[1287];
  assign N627 = data_masked[2365] | data_masked[1826];
  assign data_o[210] = N632 | data_masked[210];
  assign N632 = N631 | data_masked[749];
  assign N631 = N630 | data_masked[1288];
  assign N630 = data_masked[2366] | data_masked[1827];
  assign data_o[211] = N635 | data_masked[211];
  assign N635 = N634 | data_masked[750];
  assign N634 = N633 | data_masked[1289];
  assign N633 = data_masked[2367] | data_masked[1828];
  assign data_o[212] = N638 | data_masked[212];
  assign N638 = N637 | data_masked[751];
  assign N637 = N636 | data_masked[1290];
  assign N636 = data_masked[2368] | data_masked[1829];
  assign data_o[213] = N641 | data_masked[213];
  assign N641 = N640 | data_masked[752];
  assign N640 = N639 | data_masked[1291];
  assign N639 = data_masked[2369] | data_masked[1830];
  assign data_o[214] = N644 | data_masked[214];
  assign N644 = N643 | data_masked[753];
  assign N643 = N642 | data_masked[1292];
  assign N642 = data_masked[2370] | data_masked[1831];
  assign data_o[215] = N647 | data_masked[215];
  assign N647 = N646 | data_masked[754];
  assign N646 = N645 | data_masked[1293];
  assign N645 = data_masked[2371] | data_masked[1832];
  assign data_o[216] = N650 | data_masked[216];
  assign N650 = N649 | data_masked[755];
  assign N649 = N648 | data_masked[1294];
  assign N648 = data_masked[2372] | data_masked[1833];
  assign data_o[217] = N653 | data_masked[217];
  assign N653 = N652 | data_masked[756];
  assign N652 = N651 | data_masked[1295];
  assign N651 = data_masked[2373] | data_masked[1834];
  assign data_o[218] = N656 | data_masked[218];
  assign N656 = N655 | data_masked[757];
  assign N655 = N654 | data_masked[1296];
  assign N654 = data_masked[2374] | data_masked[1835];
  assign data_o[219] = N659 | data_masked[219];
  assign N659 = N658 | data_masked[758];
  assign N658 = N657 | data_masked[1297];
  assign N657 = data_masked[2375] | data_masked[1836];
  assign data_o[220] = N662 | data_masked[220];
  assign N662 = N661 | data_masked[759];
  assign N661 = N660 | data_masked[1298];
  assign N660 = data_masked[2376] | data_masked[1837];
  assign data_o[221] = N665 | data_masked[221];
  assign N665 = N664 | data_masked[760];
  assign N664 = N663 | data_masked[1299];
  assign N663 = data_masked[2377] | data_masked[1838];
  assign data_o[222] = N668 | data_masked[222];
  assign N668 = N667 | data_masked[761];
  assign N667 = N666 | data_masked[1300];
  assign N666 = data_masked[2378] | data_masked[1839];
  assign data_o[223] = N671 | data_masked[223];
  assign N671 = N670 | data_masked[762];
  assign N670 = N669 | data_masked[1301];
  assign N669 = data_masked[2379] | data_masked[1840];
  assign data_o[224] = N674 | data_masked[224];
  assign N674 = N673 | data_masked[763];
  assign N673 = N672 | data_masked[1302];
  assign N672 = data_masked[2380] | data_masked[1841];
  assign data_o[225] = N677 | data_masked[225];
  assign N677 = N676 | data_masked[764];
  assign N676 = N675 | data_masked[1303];
  assign N675 = data_masked[2381] | data_masked[1842];
  assign data_o[226] = N680 | data_masked[226];
  assign N680 = N679 | data_masked[765];
  assign N679 = N678 | data_masked[1304];
  assign N678 = data_masked[2382] | data_masked[1843];
  assign data_o[227] = N683 | data_masked[227];
  assign N683 = N682 | data_masked[766];
  assign N682 = N681 | data_masked[1305];
  assign N681 = data_masked[2383] | data_masked[1844];
  assign data_o[228] = N686 | data_masked[228];
  assign N686 = N685 | data_masked[767];
  assign N685 = N684 | data_masked[1306];
  assign N684 = data_masked[2384] | data_masked[1845];
  assign data_o[229] = N689 | data_masked[229];
  assign N689 = N688 | data_masked[768];
  assign N688 = N687 | data_masked[1307];
  assign N687 = data_masked[2385] | data_masked[1846];
  assign data_o[230] = N692 | data_masked[230];
  assign N692 = N691 | data_masked[769];
  assign N691 = N690 | data_masked[1308];
  assign N690 = data_masked[2386] | data_masked[1847];
  assign data_o[231] = N695 | data_masked[231];
  assign N695 = N694 | data_masked[770];
  assign N694 = N693 | data_masked[1309];
  assign N693 = data_masked[2387] | data_masked[1848];
  assign data_o[232] = N698 | data_masked[232];
  assign N698 = N697 | data_masked[771];
  assign N697 = N696 | data_masked[1310];
  assign N696 = data_masked[2388] | data_masked[1849];
  assign data_o[233] = N701 | data_masked[233];
  assign N701 = N700 | data_masked[772];
  assign N700 = N699 | data_masked[1311];
  assign N699 = data_masked[2389] | data_masked[1850];
  assign data_o[234] = N704 | data_masked[234];
  assign N704 = N703 | data_masked[773];
  assign N703 = N702 | data_masked[1312];
  assign N702 = data_masked[2390] | data_masked[1851];
  assign data_o[235] = N707 | data_masked[235];
  assign N707 = N706 | data_masked[774];
  assign N706 = N705 | data_masked[1313];
  assign N705 = data_masked[2391] | data_masked[1852];
  assign data_o[236] = N710 | data_masked[236];
  assign N710 = N709 | data_masked[775];
  assign N709 = N708 | data_masked[1314];
  assign N708 = data_masked[2392] | data_masked[1853];
  assign data_o[237] = N713 | data_masked[237];
  assign N713 = N712 | data_masked[776];
  assign N712 = N711 | data_masked[1315];
  assign N711 = data_masked[2393] | data_masked[1854];
  assign data_o[238] = N716 | data_masked[238];
  assign N716 = N715 | data_masked[777];
  assign N715 = N714 | data_masked[1316];
  assign N714 = data_masked[2394] | data_masked[1855];
  assign data_o[239] = N719 | data_masked[239];
  assign N719 = N718 | data_masked[778];
  assign N718 = N717 | data_masked[1317];
  assign N717 = data_masked[2395] | data_masked[1856];
  assign data_o[240] = N722 | data_masked[240];
  assign N722 = N721 | data_masked[779];
  assign N721 = N720 | data_masked[1318];
  assign N720 = data_masked[2396] | data_masked[1857];
  assign data_o[241] = N725 | data_masked[241];
  assign N725 = N724 | data_masked[780];
  assign N724 = N723 | data_masked[1319];
  assign N723 = data_masked[2397] | data_masked[1858];
  assign data_o[242] = N728 | data_masked[242];
  assign N728 = N727 | data_masked[781];
  assign N727 = N726 | data_masked[1320];
  assign N726 = data_masked[2398] | data_masked[1859];
  assign data_o[243] = N731 | data_masked[243];
  assign N731 = N730 | data_masked[782];
  assign N730 = N729 | data_masked[1321];
  assign N729 = data_masked[2399] | data_masked[1860];
  assign data_o[244] = N734 | data_masked[244];
  assign N734 = N733 | data_masked[783];
  assign N733 = N732 | data_masked[1322];
  assign N732 = data_masked[2400] | data_masked[1861];
  assign data_o[245] = N737 | data_masked[245];
  assign N737 = N736 | data_masked[784];
  assign N736 = N735 | data_masked[1323];
  assign N735 = data_masked[2401] | data_masked[1862];
  assign data_o[246] = N740 | data_masked[246];
  assign N740 = N739 | data_masked[785];
  assign N739 = N738 | data_masked[1324];
  assign N738 = data_masked[2402] | data_masked[1863];
  assign data_o[247] = N743 | data_masked[247];
  assign N743 = N742 | data_masked[786];
  assign N742 = N741 | data_masked[1325];
  assign N741 = data_masked[2403] | data_masked[1864];
  assign data_o[248] = N746 | data_masked[248];
  assign N746 = N745 | data_masked[787];
  assign N745 = N744 | data_masked[1326];
  assign N744 = data_masked[2404] | data_masked[1865];
  assign data_o[249] = N749 | data_masked[249];
  assign N749 = N748 | data_masked[788];
  assign N748 = N747 | data_masked[1327];
  assign N747 = data_masked[2405] | data_masked[1866];
  assign data_o[250] = N752 | data_masked[250];
  assign N752 = N751 | data_masked[789];
  assign N751 = N750 | data_masked[1328];
  assign N750 = data_masked[2406] | data_masked[1867];
  assign data_o[251] = N755 | data_masked[251];
  assign N755 = N754 | data_masked[790];
  assign N754 = N753 | data_masked[1329];
  assign N753 = data_masked[2407] | data_masked[1868];
  assign data_o[252] = N758 | data_masked[252];
  assign N758 = N757 | data_masked[791];
  assign N757 = N756 | data_masked[1330];
  assign N756 = data_masked[2408] | data_masked[1869];
  assign data_o[253] = N761 | data_masked[253];
  assign N761 = N760 | data_masked[792];
  assign N760 = N759 | data_masked[1331];
  assign N759 = data_masked[2409] | data_masked[1870];
  assign data_o[254] = N764 | data_masked[254];
  assign N764 = N763 | data_masked[793];
  assign N763 = N762 | data_masked[1332];
  assign N762 = data_masked[2410] | data_masked[1871];
  assign data_o[255] = N767 | data_masked[255];
  assign N767 = N766 | data_masked[794];
  assign N766 = N765 | data_masked[1333];
  assign N765 = data_masked[2411] | data_masked[1872];
  assign data_o[256] = N770 | data_masked[256];
  assign N770 = N769 | data_masked[795];
  assign N769 = N768 | data_masked[1334];
  assign N768 = data_masked[2412] | data_masked[1873];
  assign data_o[257] = N773 | data_masked[257];
  assign N773 = N772 | data_masked[796];
  assign N772 = N771 | data_masked[1335];
  assign N771 = data_masked[2413] | data_masked[1874];
  assign data_o[258] = N776 | data_masked[258];
  assign N776 = N775 | data_masked[797];
  assign N775 = N774 | data_masked[1336];
  assign N774 = data_masked[2414] | data_masked[1875];
  assign data_o[259] = N779 | data_masked[259];
  assign N779 = N778 | data_masked[798];
  assign N778 = N777 | data_masked[1337];
  assign N777 = data_masked[2415] | data_masked[1876];
  assign data_o[260] = N782 | data_masked[260];
  assign N782 = N781 | data_masked[799];
  assign N781 = N780 | data_masked[1338];
  assign N780 = data_masked[2416] | data_masked[1877];
  assign data_o[261] = N785 | data_masked[261];
  assign N785 = N784 | data_masked[800];
  assign N784 = N783 | data_masked[1339];
  assign N783 = data_masked[2417] | data_masked[1878];
  assign data_o[262] = N788 | data_masked[262];
  assign N788 = N787 | data_masked[801];
  assign N787 = N786 | data_masked[1340];
  assign N786 = data_masked[2418] | data_masked[1879];
  assign data_o[263] = N791 | data_masked[263];
  assign N791 = N790 | data_masked[802];
  assign N790 = N789 | data_masked[1341];
  assign N789 = data_masked[2419] | data_masked[1880];
  assign data_o[264] = N794 | data_masked[264];
  assign N794 = N793 | data_masked[803];
  assign N793 = N792 | data_masked[1342];
  assign N792 = data_masked[2420] | data_masked[1881];
  assign data_o[265] = N797 | data_masked[265];
  assign N797 = N796 | data_masked[804];
  assign N796 = N795 | data_masked[1343];
  assign N795 = data_masked[2421] | data_masked[1882];
  assign data_o[266] = N800 | data_masked[266];
  assign N800 = N799 | data_masked[805];
  assign N799 = N798 | data_masked[1344];
  assign N798 = data_masked[2422] | data_masked[1883];
  assign data_o[267] = N803 | data_masked[267];
  assign N803 = N802 | data_masked[806];
  assign N802 = N801 | data_masked[1345];
  assign N801 = data_masked[2423] | data_masked[1884];
  assign data_o[268] = N806 | data_masked[268];
  assign N806 = N805 | data_masked[807];
  assign N805 = N804 | data_masked[1346];
  assign N804 = data_masked[2424] | data_masked[1885];
  assign data_o[269] = N809 | data_masked[269];
  assign N809 = N808 | data_masked[808];
  assign N808 = N807 | data_masked[1347];
  assign N807 = data_masked[2425] | data_masked[1886];
  assign data_o[270] = N812 | data_masked[270];
  assign N812 = N811 | data_masked[809];
  assign N811 = N810 | data_masked[1348];
  assign N810 = data_masked[2426] | data_masked[1887];
  assign data_o[271] = N815 | data_masked[271];
  assign N815 = N814 | data_masked[810];
  assign N814 = N813 | data_masked[1349];
  assign N813 = data_masked[2427] | data_masked[1888];
  assign data_o[272] = N818 | data_masked[272];
  assign N818 = N817 | data_masked[811];
  assign N817 = N816 | data_masked[1350];
  assign N816 = data_masked[2428] | data_masked[1889];
  assign data_o[273] = N821 | data_masked[273];
  assign N821 = N820 | data_masked[812];
  assign N820 = N819 | data_masked[1351];
  assign N819 = data_masked[2429] | data_masked[1890];
  assign data_o[274] = N824 | data_masked[274];
  assign N824 = N823 | data_masked[813];
  assign N823 = N822 | data_masked[1352];
  assign N822 = data_masked[2430] | data_masked[1891];
  assign data_o[275] = N827 | data_masked[275];
  assign N827 = N826 | data_masked[814];
  assign N826 = N825 | data_masked[1353];
  assign N825 = data_masked[2431] | data_masked[1892];
  assign data_o[276] = N830 | data_masked[276];
  assign N830 = N829 | data_masked[815];
  assign N829 = N828 | data_masked[1354];
  assign N828 = data_masked[2432] | data_masked[1893];
  assign data_o[277] = N833 | data_masked[277];
  assign N833 = N832 | data_masked[816];
  assign N832 = N831 | data_masked[1355];
  assign N831 = data_masked[2433] | data_masked[1894];
  assign data_o[278] = N836 | data_masked[278];
  assign N836 = N835 | data_masked[817];
  assign N835 = N834 | data_masked[1356];
  assign N834 = data_masked[2434] | data_masked[1895];
  assign data_o[279] = N839 | data_masked[279];
  assign N839 = N838 | data_masked[818];
  assign N838 = N837 | data_masked[1357];
  assign N837 = data_masked[2435] | data_masked[1896];
  assign data_o[280] = N842 | data_masked[280];
  assign N842 = N841 | data_masked[819];
  assign N841 = N840 | data_masked[1358];
  assign N840 = data_masked[2436] | data_masked[1897];
  assign data_o[281] = N845 | data_masked[281];
  assign N845 = N844 | data_masked[820];
  assign N844 = N843 | data_masked[1359];
  assign N843 = data_masked[2437] | data_masked[1898];
  assign data_o[282] = N848 | data_masked[282];
  assign N848 = N847 | data_masked[821];
  assign N847 = N846 | data_masked[1360];
  assign N846 = data_masked[2438] | data_masked[1899];
  assign data_o[283] = N851 | data_masked[283];
  assign N851 = N850 | data_masked[822];
  assign N850 = N849 | data_masked[1361];
  assign N849 = data_masked[2439] | data_masked[1900];
  assign data_o[284] = N854 | data_masked[284];
  assign N854 = N853 | data_masked[823];
  assign N853 = N852 | data_masked[1362];
  assign N852 = data_masked[2440] | data_masked[1901];
  assign data_o[285] = N857 | data_masked[285];
  assign N857 = N856 | data_masked[824];
  assign N856 = N855 | data_masked[1363];
  assign N855 = data_masked[2441] | data_masked[1902];
  assign data_o[286] = N860 | data_masked[286];
  assign N860 = N859 | data_masked[825];
  assign N859 = N858 | data_masked[1364];
  assign N858 = data_masked[2442] | data_masked[1903];
  assign data_o[287] = N863 | data_masked[287];
  assign N863 = N862 | data_masked[826];
  assign N862 = N861 | data_masked[1365];
  assign N861 = data_masked[2443] | data_masked[1904];
  assign data_o[288] = N866 | data_masked[288];
  assign N866 = N865 | data_masked[827];
  assign N865 = N864 | data_masked[1366];
  assign N864 = data_masked[2444] | data_masked[1905];
  assign data_o[289] = N869 | data_masked[289];
  assign N869 = N868 | data_masked[828];
  assign N868 = N867 | data_masked[1367];
  assign N867 = data_masked[2445] | data_masked[1906];
  assign data_o[290] = N872 | data_masked[290];
  assign N872 = N871 | data_masked[829];
  assign N871 = N870 | data_masked[1368];
  assign N870 = data_masked[2446] | data_masked[1907];
  assign data_o[291] = N875 | data_masked[291];
  assign N875 = N874 | data_masked[830];
  assign N874 = N873 | data_masked[1369];
  assign N873 = data_masked[2447] | data_masked[1908];
  assign data_o[292] = N878 | data_masked[292];
  assign N878 = N877 | data_masked[831];
  assign N877 = N876 | data_masked[1370];
  assign N876 = data_masked[2448] | data_masked[1909];
  assign data_o[293] = N881 | data_masked[293];
  assign N881 = N880 | data_masked[832];
  assign N880 = N879 | data_masked[1371];
  assign N879 = data_masked[2449] | data_masked[1910];
  assign data_o[294] = N884 | data_masked[294];
  assign N884 = N883 | data_masked[833];
  assign N883 = N882 | data_masked[1372];
  assign N882 = data_masked[2450] | data_masked[1911];
  assign data_o[295] = N887 | data_masked[295];
  assign N887 = N886 | data_masked[834];
  assign N886 = N885 | data_masked[1373];
  assign N885 = data_masked[2451] | data_masked[1912];
  assign data_o[296] = N890 | data_masked[296];
  assign N890 = N889 | data_masked[835];
  assign N889 = N888 | data_masked[1374];
  assign N888 = data_masked[2452] | data_masked[1913];
  assign data_o[297] = N893 | data_masked[297];
  assign N893 = N892 | data_masked[836];
  assign N892 = N891 | data_masked[1375];
  assign N891 = data_masked[2453] | data_masked[1914];
  assign data_o[298] = N896 | data_masked[298];
  assign N896 = N895 | data_masked[837];
  assign N895 = N894 | data_masked[1376];
  assign N894 = data_masked[2454] | data_masked[1915];
  assign data_o[299] = N899 | data_masked[299];
  assign N899 = N898 | data_masked[838];
  assign N898 = N897 | data_masked[1377];
  assign N897 = data_masked[2455] | data_masked[1916];
  assign data_o[300] = N902 | data_masked[300];
  assign N902 = N901 | data_masked[839];
  assign N901 = N900 | data_masked[1378];
  assign N900 = data_masked[2456] | data_masked[1917];
  assign data_o[301] = N905 | data_masked[301];
  assign N905 = N904 | data_masked[840];
  assign N904 = N903 | data_masked[1379];
  assign N903 = data_masked[2457] | data_masked[1918];
  assign data_o[302] = N908 | data_masked[302];
  assign N908 = N907 | data_masked[841];
  assign N907 = N906 | data_masked[1380];
  assign N906 = data_masked[2458] | data_masked[1919];
  assign data_o[303] = N911 | data_masked[303];
  assign N911 = N910 | data_masked[842];
  assign N910 = N909 | data_masked[1381];
  assign N909 = data_masked[2459] | data_masked[1920];
  assign data_o[304] = N914 | data_masked[304];
  assign N914 = N913 | data_masked[843];
  assign N913 = N912 | data_masked[1382];
  assign N912 = data_masked[2460] | data_masked[1921];
  assign data_o[305] = N917 | data_masked[305];
  assign N917 = N916 | data_masked[844];
  assign N916 = N915 | data_masked[1383];
  assign N915 = data_masked[2461] | data_masked[1922];
  assign data_o[306] = N920 | data_masked[306];
  assign N920 = N919 | data_masked[845];
  assign N919 = N918 | data_masked[1384];
  assign N918 = data_masked[2462] | data_masked[1923];
  assign data_o[307] = N923 | data_masked[307];
  assign N923 = N922 | data_masked[846];
  assign N922 = N921 | data_masked[1385];
  assign N921 = data_masked[2463] | data_masked[1924];
  assign data_o[308] = N926 | data_masked[308];
  assign N926 = N925 | data_masked[847];
  assign N925 = N924 | data_masked[1386];
  assign N924 = data_masked[2464] | data_masked[1925];
  assign data_o[309] = N929 | data_masked[309];
  assign N929 = N928 | data_masked[848];
  assign N928 = N927 | data_masked[1387];
  assign N927 = data_masked[2465] | data_masked[1926];
  assign data_o[310] = N932 | data_masked[310];
  assign N932 = N931 | data_masked[849];
  assign N931 = N930 | data_masked[1388];
  assign N930 = data_masked[2466] | data_masked[1927];
  assign data_o[311] = N935 | data_masked[311];
  assign N935 = N934 | data_masked[850];
  assign N934 = N933 | data_masked[1389];
  assign N933 = data_masked[2467] | data_masked[1928];
  assign data_o[312] = N938 | data_masked[312];
  assign N938 = N937 | data_masked[851];
  assign N937 = N936 | data_masked[1390];
  assign N936 = data_masked[2468] | data_masked[1929];
  assign data_o[313] = N941 | data_masked[313];
  assign N941 = N940 | data_masked[852];
  assign N940 = N939 | data_masked[1391];
  assign N939 = data_masked[2469] | data_masked[1930];
  assign data_o[314] = N944 | data_masked[314];
  assign N944 = N943 | data_masked[853];
  assign N943 = N942 | data_masked[1392];
  assign N942 = data_masked[2470] | data_masked[1931];
  assign data_o[315] = N947 | data_masked[315];
  assign N947 = N946 | data_masked[854];
  assign N946 = N945 | data_masked[1393];
  assign N945 = data_masked[2471] | data_masked[1932];
  assign data_o[316] = N950 | data_masked[316];
  assign N950 = N949 | data_masked[855];
  assign N949 = N948 | data_masked[1394];
  assign N948 = data_masked[2472] | data_masked[1933];
  assign data_o[317] = N953 | data_masked[317];
  assign N953 = N952 | data_masked[856];
  assign N952 = N951 | data_masked[1395];
  assign N951 = data_masked[2473] | data_masked[1934];
  assign data_o[318] = N956 | data_masked[318];
  assign N956 = N955 | data_masked[857];
  assign N955 = N954 | data_masked[1396];
  assign N954 = data_masked[2474] | data_masked[1935];
  assign data_o[319] = N959 | data_masked[319];
  assign N959 = N958 | data_masked[858];
  assign N958 = N957 | data_masked[1397];
  assign N957 = data_masked[2475] | data_masked[1936];
  assign data_o[320] = N962 | data_masked[320];
  assign N962 = N961 | data_masked[859];
  assign N961 = N960 | data_masked[1398];
  assign N960 = data_masked[2476] | data_masked[1937];
  assign data_o[321] = N965 | data_masked[321];
  assign N965 = N964 | data_masked[860];
  assign N964 = N963 | data_masked[1399];
  assign N963 = data_masked[2477] | data_masked[1938];
  assign data_o[322] = N968 | data_masked[322];
  assign N968 = N967 | data_masked[861];
  assign N967 = N966 | data_masked[1400];
  assign N966 = data_masked[2478] | data_masked[1939];
  assign data_o[323] = N971 | data_masked[323];
  assign N971 = N970 | data_masked[862];
  assign N970 = N969 | data_masked[1401];
  assign N969 = data_masked[2479] | data_masked[1940];
  assign data_o[324] = N974 | data_masked[324];
  assign N974 = N973 | data_masked[863];
  assign N973 = N972 | data_masked[1402];
  assign N972 = data_masked[2480] | data_masked[1941];
  assign data_o[325] = N977 | data_masked[325];
  assign N977 = N976 | data_masked[864];
  assign N976 = N975 | data_masked[1403];
  assign N975 = data_masked[2481] | data_masked[1942];
  assign data_o[326] = N980 | data_masked[326];
  assign N980 = N979 | data_masked[865];
  assign N979 = N978 | data_masked[1404];
  assign N978 = data_masked[2482] | data_masked[1943];
  assign data_o[327] = N983 | data_masked[327];
  assign N983 = N982 | data_masked[866];
  assign N982 = N981 | data_masked[1405];
  assign N981 = data_masked[2483] | data_masked[1944];
  assign data_o[328] = N986 | data_masked[328];
  assign N986 = N985 | data_masked[867];
  assign N985 = N984 | data_masked[1406];
  assign N984 = data_masked[2484] | data_masked[1945];
  assign data_o[329] = N989 | data_masked[329];
  assign N989 = N988 | data_masked[868];
  assign N988 = N987 | data_masked[1407];
  assign N987 = data_masked[2485] | data_masked[1946];
  assign data_o[330] = N992 | data_masked[330];
  assign N992 = N991 | data_masked[869];
  assign N991 = N990 | data_masked[1408];
  assign N990 = data_masked[2486] | data_masked[1947];
  assign data_o[331] = N995 | data_masked[331];
  assign N995 = N994 | data_masked[870];
  assign N994 = N993 | data_masked[1409];
  assign N993 = data_masked[2487] | data_masked[1948];
  assign data_o[332] = N998 | data_masked[332];
  assign N998 = N997 | data_masked[871];
  assign N997 = N996 | data_masked[1410];
  assign N996 = data_masked[2488] | data_masked[1949];
  assign data_o[333] = N1001 | data_masked[333];
  assign N1001 = N1000 | data_masked[872];
  assign N1000 = N999 | data_masked[1411];
  assign N999 = data_masked[2489] | data_masked[1950];
  assign data_o[334] = N1004 | data_masked[334];
  assign N1004 = N1003 | data_masked[873];
  assign N1003 = N1002 | data_masked[1412];
  assign N1002 = data_masked[2490] | data_masked[1951];
  assign data_o[335] = N1007 | data_masked[335];
  assign N1007 = N1006 | data_masked[874];
  assign N1006 = N1005 | data_masked[1413];
  assign N1005 = data_masked[2491] | data_masked[1952];
  assign data_o[336] = N1010 | data_masked[336];
  assign N1010 = N1009 | data_masked[875];
  assign N1009 = N1008 | data_masked[1414];
  assign N1008 = data_masked[2492] | data_masked[1953];
  assign data_o[337] = N1013 | data_masked[337];
  assign N1013 = N1012 | data_masked[876];
  assign N1012 = N1011 | data_masked[1415];
  assign N1011 = data_masked[2493] | data_masked[1954];
  assign data_o[338] = N1016 | data_masked[338];
  assign N1016 = N1015 | data_masked[877];
  assign N1015 = N1014 | data_masked[1416];
  assign N1014 = data_masked[2494] | data_masked[1955];
  assign data_o[339] = N1019 | data_masked[339];
  assign N1019 = N1018 | data_masked[878];
  assign N1018 = N1017 | data_masked[1417];
  assign N1017 = data_masked[2495] | data_masked[1956];
  assign data_o[340] = N1022 | data_masked[340];
  assign N1022 = N1021 | data_masked[879];
  assign N1021 = N1020 | data_masked[1418];
  assign N1020 = data_masked[2496] | data_masked[1957];
  assign data_o[341] = N1025 | data_masked[341];
  assign N1025 = N1024 | data_masked[880];
  assign N1024 = N1023 | data_masked[1419];
  assign N1023 = data_masked[2497] | data_masked[1958];
  assign data_o[342] = N1028 | data_masked[342];
  assign N1028 = N1027 | data_masked[881];
  assign N1027 = N1026 | data_masked[1420];
  assign N1026 = data_masked[2498] | data_masked[1959];
  assign data_o[343] = N1031 | data_masked[343];
  assign N1031 = N1030 | data_masked[882];
  assign N1030 = N1029 | data_masked[1421];
  assign N1029 = data_masked[2499] | data_masked[1960];
  assign data_o[344] = N1034 | data_masked[344];
  assign N1034 = N1033 | data_masked[883];
  assign N1033 = N1032 | data_masked[1422];
  assign N1032 = data_masked[2500] | data_masked[1961];
  assign data_o[345] = N1037 | data_masked[345];
  assign N1037 = N1036 | data_masked[884];
  assign N1036 = N1035 | data_masked[1423];
  assign N1035 = data_masked[2501] | data_masked[1962];
  assign data_o[346] = N1040 | data_masked[346];
  assign N1040 = N1039 | data_masked[885];
  assign N1039 = N1038 | data_masked[1424];
  assign N1038 = data_masked[2502] | data_masked[1963];
  assign data_o[347] = N1043 | data_masked[347];
  assign N1043 = N1042 | data_masked[886];
  assign N1042 = N1041 | data_masked[1425];
  assign N1041 = data_masked[2503] | data_masked[1964];
  assign data_o[348] = N1046 | data_masked[348];
  assign N1046 = N1045 | data_masked[887];
  assign N1045 = N1044 | data_masked[1426];
  assign N1044 = data_masked[2504] | data_masked[1965];
  assign data_o[349] = N1049 | data_masked[349];
  assign N1049 = N1048 | data_masked[888];
  assign N1048 = N1047 | data_masked[1427];
  assign N1047 = data_masked[2505] | data_masked[1966];
  assign data_o[350] = N1052 | data_masked[350];
  assign N1052 = N1051 | data_masked[889];
  assign N1051 = N1050 | data_masked[1428];
  assign N1050 = data_masked[2506] | data_masked[1967];
  assign data_o[351] = N1055 | data_masked[351];
  assign N1055 = N1054 | data_masked[890];
  assign N1054 = N1053 | data_masked[1429];
  assign N1053 = data_masked[2507] | data_masked[1968];
  assign data_o[352] = N1058 | data_masked[352];
  assign N1058 = N1057 | data_masked[891];
  assign N1057 = N1056 | data_masked[1430];
  assign N1056 = data_masked[2508] | data_masked[1969];
  assign data_o[353] = N1061 | data_masked[353];
  assign N1061 = N1060 | data_masked[892];
  assign N1060 = N1059 | data_masked[1431];
  assign N1059 = data_masked[2509] | data_masked[1970];
  assign data_o[354] = N1064 | data_masked[354];
  assign N1064 = N1063 | data_masked[893];
  assign N1063 = N1062 | data_masked[1432];
  assign N1062 = data_masked[2510] | data_masked[1971];
  assign data_o[355] = N1067 | data_masked[355];
  assign N1067 = N1066 | data_masked[894];
  assign N1066 = N1065 | data_masked[1433];
  assign N1065 = data_masked[2511] | data_masked[1972];
  assign data_o[356] = N1070 | data_masked[356];
  assign N1070 = N1069 | data_masked[895];
  assign N1069 = N1068 | data_masked[1434];
  assign N1068 = data_masked[2512] | data_masked[1973];
  assign data_o[357] = N1073 | data_masked[357];
  assign N1073 = N1072 | data_masked[896];
  assign N1072 = N1071 | data_masked[1435];
  assign N1071 = data_masked[2513] | data_masked[1974];
  assign data_o[358] = N1076 | data_masked[358];
  assign N1076 = N1075 | data_masked[897];
  assign N1075 = N1074 | data_masked[1436];
  assign N1074 = data_masked[2514] | data_masked[1975];
  assign data_o[359] = N1079 | data_masked[359];
  assign N1079 = N1078 | data_masked[898];
  assign N1078 = N1077 | data_masked[1437];
  assign N1077 = data_masked[2515] | data_masked[1976];
  assign data_o[360] = N1082 | data_masked[360];
  assign N1082 = N1081 | data_masked[899];
  assign N1081 = N1080 | data_masked[1438];
  assign N1080 = data_masked[2516] | data_masked[1977];
  assign data_o[361] = N1085 | data_masked[361];
  assign N1085 = N1084 | data_masked[900];
  assign N1084 = N1083 | data_masked[1439];
  assign N1083 = data_masked[2517] | data_masked[1978];
  assign data_o[362] = N1088 | data_masked[362];
  assign N1088 = N1087 | data_masked[901];
  assign N1087 = N1086 | data_masked[1440];
  assign N1086 = data_masked[2518] | data_masked[1979];
  assign data_o[363] = N1091 | data_masked[363];
  assign N1091 = N1090 | data_masked[902];
  assign N1090 = N1089 | data_masked[1441];
  assign N1089 = data_masked[2519] | data_masked[1980];
  assign data_o[364] = N1094 | data_masked[364];
  assign N1094 = N1093 | data_masked[903];
  assign N1093 = N1092 | data_masked[1442];
  assign N1092 = data_masked[2520] | data_masked[1981];
  assign data_o[365] = N1097 | data_masked[365];
  assign N1097 = N1096 | data_masked[904];
  assign N1096 = N1095 | data_masked[1443];
  assign N1095 = data_masked[2521] | data_masked[1982];
  assign data_o[366] = N1100 | data_masked[366];
  assign N1100 = N1099 | data_masked[905];
  assign N1099 = N1098 | data_masked[1444];
  assign N1098 = data_masked[2522] | data_masked[1983];
  assign data_o[367] = N1103 | data_masked[367];
  assign N1103 = N1102 | data_masked[906];
  assign N1102 = N1101 | data_masked[1445];
  assign N1101 = data_masked[2523] | data_masked[1984];
  assign data_o[368] = N1106 | data_masked[368];
  assign N1106 = N1105 | data_masked[907];
  assign N1105 = N1104 | data_masked[1446];
  assign N1104 = data_masked[2524] | data_masked[1985];
  assign data_o[369] = N1109 | data_masked[369];
  assign N1109 = N1108 | data_masked[908];
  assign N1108 = N1107 | data_masked[1447];
  assign N1107 = data_masked[2525] | data_masked[1986];
  assign data_o[370] = N1112 | data_masked[370];
  assign N1112 = N1111 | data_masked[909];
  assign N1111 = N1110 | data_masked[1448];
  assign N1110 = data_masked[2526] | data_masked[1987];
  assign data_o[371] = N1115 | data_masked[371];
  assign N1115 = N1114 | data_masked[910];
  assign N1114 = N1113 | data_masked[1449];
  assign N1113 = data_masked[2527] | data_masked[1988];
  assign data_o[372] = N1118 | data_masked[372];
  assign N1118 = N1117 | data_masked[911];
  assign N1117 = N1116 | data_masked[1450];
  assign N1116 = data_masked[2528] | data_masked[1989];
  assign data_o[373] = N1121 | data_masked[373];
  assign N1121 = N1120 | data_masked[912];
  assign N1120 = N1119 | data_masked[1451];
  assign N1119 = data_masked[2529] | data_masked[1990];
  assign data_o[374] = N1124 | data_masked[374];
  assign N1124 = N1123 | data_masked[913];
  assign N1123 = N1122 | data_masked[1452];
  assign N1122 = data_masked[2530] | data_masked[1991];
  assign data_o[375] = N1127 | data_masked[375];
  assign N1127 = N1126 | data_masked[914];
  assign N1126 = N1125 | data_masked[1453];
  assign N1125 = data_masked[2531] | data_masked[1992];
  assign data_o[376] = N1130 | data_masked[376];
  assign N1130 = N1129 | data_masked[915];
  assign N1129 = N1128 | data_masked[1454];
  assign N1128 = data_masked[2532] | data_masked[1993];
  assign data_o[377] = N1133 | data_masked[377];
  assign N1133 = N1132 | data_masked[916];
  assign N1132 = N1131 | data_masked[1455];
  assign N1131 = data_masked[2533] | data_masked[1994];
  assign data_o[378] = N1136 | data_masked[378];
  assign N1136 = N1135 | data_masked[917];
  assign N1135 = N1134 | data_masked[1456];
  assign N1134 = data_masked[2534] | data_masked[1995];
  assign data_o[379] = N1139 | data_masked[379];
  assign N1139 = N1138 | data_masked[918];
  assign N1138 = N1137 | data_masked[1457];
  assign N1137 = data_masked[2535] | data_masked[1996];
  assign data_o[380] = N1142 | data_masked[380];
  assign N1142 = N1141 | data_masked[919];
  assign N1141 = N1140 | data_masked[1458];
  assign N1140 = data_masked[2536] | data_masked[1997];
  assign data_o[381] = N1145 | data_masked[381];
  assign N1145 = N1144 | data_masked[920];
  assign N1144 = N1143 | data_masked[1459];
  assign N1143 = data_masked[2537] | data_masked[1998];
  assign data_o[382] = N1148 | data_masked[382];
  assign N1148 = N1147 | data_masked[921];
  assign N1147 = N1146 | data_masked[1460];
  assign N1146 = data_masked[2538] | data_masked[1999];
  assign data_o[383] = N1151 | data_masked[383];
  assign N1151 = N1150 | data_masked[922];
  assign N1150 = N1149 | data_masked[1461];
  assign N1149 = data_masked[2539] | data_masked[2000];
  assign data_o[384] = N1154 | data_masked[384];
  assign N1154 = N1153 | data_masked[923];
  assign N1153 = N1152 | data_masked[1462];
  assign N1152 = data_masked[2540] | data_masked[2001];
  assign data_o[385] = N1157 | data_masked[385];
  assign N1157 = N1156 | data_masked[924];
  assign N1156 = N1155 | data_masked[1463];
  assign N1155 = data_masked[2541] | data_masked[2002];
  assign data_o[386] = N1160 | data_masked[386];
  assign N1160 = N1159 | data_masked[925];
  assign N1159 = N1158 | data_masked[1464];
  assign N1158 = data_masked[2542] | data_masked[2003];
  assign data_o[387] = N1163 | data_masked[387];
  assign N1163 = N1162 | data_masked[926];
  assign N1162 = N1161 | data_masked[1465];
  assign N1161 = data_masked[2543] | data_masked[2004];
  assign data_o[388] = N1166 | data_masked[388];
  assign N1166 = N1165 | data_masked[927];
  assign N1165 = N1164 | data_masked[1466];
  assign N1164 = data_masked[2544] | data_masked[2005];
  assign data_o[389] = N1169 | data_masked[389];
  assign N1169 = N1168 | data_masked[928];
  assign N1168 = N1167 | data_masked[1467];
  assign N1167 = data_masked[2545] | data_masked[2006];
  assign data_o[390] = N1172 | data_masked[390];
  assign N1172 = N1171 | data_masked[929];
  assign N1171 = N1170 | data_masked[1468];
  assign N1170 = data_masked[2546] | data_masked[2007];
  assign data_o[391] = N1175 | data_masked[391];
  assign N1175 = N1174 | data_masked[930];
  assign N1174 = N1173 | data_masked[1469];
  assign N1173 = data_masked[2547] | data_masked[2008];
  assign data_o[392] = N1178 | data_masked[392];
  assign N1178 = N1177 | data_masked[931];
  assign N1177 = N1176 | data_masked[1470];
  assign N1176 = data_masked[2548] | data_masked[2009];
  assign data_o[393] = N1181 | data_masked[393];
  assign N1181 = N1180 | data_masked[932];
  assign N1180 = N1179 | data_masked[1471];
  assign N1179 = data_masked[2549] | data_masked[2010];
  assign data_o[394] = N1184 | data_masked[394];
  assign N1184 = N1183 | data_masked[933];
  assign N1183 = N1182 | data_masked[1472];
  assign N1182 = data_masked[2550] | data_masked[2011];
  assign data_o[395] = N1187 | data_masked[395];
  assign N1187 = N1186 | data_masked[934];
  assign N1186 = N1185 | data_masked[1473];
  assign N1185 = data_masked[2551] | data_masked[2012];
  assign data_o[396] = N1190 | data_masked[396];
  assign N1190 = N1189 | data_masked[935];
  assign N1189 = N1188 | data_masked[1474];
  assign N1188 = data_masked[2552] | data_masked[2013];
  assign data_o[397] = N1193 | data_masked[397];
  assign N1193 = N1192 | data_masked[936];
  assign N1192 = N1191 | data_masked[1475];
  assign N1191 = data_masked[2553] | data_masked[2014];
  assign data_o[398] = N1196 | data_masked[398];
  assign N1196 = N1195 | data_masked[937];
  assign N1195 = N1194 | data_masked[1476];
  assign N1194 = data_masked[2554] | data_masked[2015];
  assign data_o[399] = N1199 | data_masked[399];
  assign N1199 = N1198 | data_masked[938];
  assign N1198 = N1197 | data_masked[1477];
  assign N1197 = data_masked[2555] | data_masked[2016];
  assign data_o[400] = N1202 | data_masked[400];
  assign N1202 = N1201 | data_masked[939];
  assign N1201 = N1200 | data_masked[1478];
  assign N1200 = data_masked[2556] | data_masked[2017];
  assign data_o[401] = N1205 | data_masked[401];
  assign N1205 = N1204 | data_masked[940];
  assign N1204 = N1203 | data_masked[1479];
  assign N1203 = data_masked[2557] | data_masked[2018];
  assign data_o[402] = N1208 | data_masked[402];
  assign N1208 = N1207 | data_masked[941];
  assign N1207 = N1206 | data_masked[1480];
  assign N1206 = data_masked[2558] | data_masked[2019];
  assign data_o[403] = N1211 | data_masked[403];
  assign N1211 = N1210 | data_masked[942];
  assign N1210 = N1209 | data_masked[1481];
  assign N1209 = data_masked[2559] | data_masked[2020];
  assign data_o[404] = N1214 | data_masked[404];
  assign N1214 = N1213 | data_masked[943];
  assign N1213 = N1212 | data_masked[1482];
  assign N1212 = data_masked[2560] | data_masked[2021];
  assign data_o[405] = N1217 | data_masked[405];
  assign N1217 = N1216 | data_masked[944];
  assign N1216 = N1215 | data_masked[1483];
  assign N1215 = data_masked[2561] | data_masked[2022];
  assign data_o[406] = N1220 | data_masked[406];
  assign N1220 = N1219 | data_masked[945];
  assign N1219 = N1218 | data_masked[1484];
  assign N1218 = data_masked[2562] | data_masked[2023];
  assign data_o[407] = N1223 | data_masked[407];
  assign N1223 = N1222 | data_masked[946];
  assign N1222 = N1221 | data_masked[1485];
  assign N1221 = data_masked[2563] | data_masked[2024];
  assign data_o[408] = N1226 | data_masked[408];
  assign N1226 = N1225 | data_masked[947];
  assign N1225 = N1224 | data_masked[1486];
  assign N1224 = data_masked[2564] | data_masked[2025];
  assign data_o[409] = N1229 | data_masked[409];
  assign N1229 = N1228 | data_masked[948];
  assign N1228 = N1227 | data_masked[1487];
  assign N1227 = data_masked[2565] | data_masked[2026];
  assign data_o[410] = N1232 | data_masked[410];
  assign N1232 = N1231 | data_masked[949];
  assign N1231 = N1230 | data_masked[1488];
  assign N1230 = data_masked[2566] | data_masked[2027];
  assign data_o[411] = N1235 | data_masked[411];
  assign N1235 = N1234 | data_masked[950];
  assign N1234 = N1233 | data_masked[1489];
  assign N1233 = data_masked[2567] | data_masked[2028];
  assign data_o[412] = N1238 | data_masked[412];
  assign N1238 = N1237 | data_masked[951];
  assign N1237 = N1236 | data_masked[1490];
  assign N1236 = data_masked[2568] | data_masked[2029];
  assign data_o[413] = N1241 | data_masked[413];
  assign N1241 = N1240 | data_masked[952];
  assign N1240 = N1239 | data_masked[1491];
  assign N1239 = data_masked[2569] | data_masked[2030];
  assign data_o[414] = N1244 | data_masked[414];
  assign N1244 = N1243 | data_masked[953];
  assign N1243 = N1242 | data_masked[1492];
  assign N1242 = data_masked[2570] | data_masked[2031];
  assign data_o[415] = N1247 | data_masked[415];
  assign N1247 = N1246 | data_masked[954];
  assign N1246 = N1245 | data_masked[1493];
  assign N1245 = data_masked[2571] | data_masked[2032];
  assign data_o[416] = N1250 | data_masked[416];
  assign N1250 = N1249 | data_masked[955];
  assign N1249 = N1248 | data_masked[1494];
  assign N1248 = data_masked[2572] | data_masked[2033];
  assign data_o[417] = N1253 | data_masked[417];
  assign N1253 = N1252 | data_masked[956];
  assign N1252 = N1251 | data_masked[1495];
  assign N1251 = data_masked[2573] | data_masked[2034];
  assign data_o[418] = N1256 | data_masked[418];
  assign N1256 = N1255 | data_masked[957];
  assign N1255 = N1254 | data_masked[1496];
  assign N1254 = data_masked[2574] | data_masked[2035];
  assign data_o[419] = N1259 | data_masked[419];
  assign N1259 = N1258 | data_masked[958];
  assign N1258 = N1257 | data_masked[1497];
  assign N1257 = data_masked[2575] | data_masked[2036];
  assign data_o[420] = N1262 | data_masked[420];
  assign N1262 = N1261 | data_masked[959];
  assign N1261 = N1260 | data_masked[1498];
  assign N1260 = data_masked[2576] | data_masked[2037];
  assign data_o[421] = N1265 | data_masked[421];
  assign N1265 = N1264 | data_masked[960];
  assign N1264 = N1263 | data_masked[1499];
  assign N1263 = data_masked[2577] | data_masked[2038];
  assign data_o[422] = N1268 | data_masked[422];
  assign N1268 = N1267 | data_masked[961];
  assign N1267 = N1266 | data_masked[1500];
  assign N1266 = data_masked[2578] | data_masked[2039];
  assign data_o[423] = N1271 | data_masked[423];
  assign N1271 = N1270 | data_masked[962];
  assign N1270 = N1269 | data_masked[1501];
  assign N1269 = data_masked[2579] | data_masked[2040];
  assign data_o[424] = N1274 | data_masked[424];
  assign N1274 = N1273 | data_masked[963];
  assign N1273 = N1272 | data_masked[1502];
  assign N1272 = data_masked[2580] | data_masked[2041];
  assign data_o[425] = N1277 | data_masked[425];
  assign N1277 = N1276 | data_masked[964];
  assign N1276 = N1275 | data_masked[1503];
  assign N1275 = data_masked[2581] | data_masked[2042];
  assign data_o[426] = N1280 | data_masked[426];
  assign N1280 = N1279 | data_masked[965];
  assign N1279 = N1278 | data_masked[1504];
  assign N1278 = data_masked[2582] | data_masked[2043];
  assign data_o[427] = N1283 | data_masked[427];
  assign N1283 = N1282 | data_masked[966];
  assign N1282 = N1281 | data_masked[1505];
  assign N1281 = data_masked[2583] | data_masked[2044];
  assign data_o[428] = N1286 | data_masked[428];
  assign N1286 = N1285 | data_masked[967];
  assign N1285 = N1284 | data_masked[1506];
  assign N1284 = data_masked[2584] | data_masked[2045];
  assign data_o[429] = N1289 | data_masked[429];
  assign N1289 = N1288 | data_masked[968];
  assign N1288 = N1287 | data_masked[1507];
  assign N1287 = data_masked[2585] | data_masked[2046];
  assign data_o[430] = N1292 | data_masked[430];
  assign N1292 = N1291 | data_masked[969];
  assign N1291 = N1290 | data_masked[1508];
  assign N1290 = data_masked[2586] | data_masked[2047];
  assign data_o[431] = N1295 | data_masked[431];
  assign N1295 = N1294 | data_masked[970];
  assign N1294 = N1293 | data_masked[1509];
  assign N1293 = data_masked[2587] | data_masked[2048];
  assign data_o[432] = N1298 | data_masked[432];
  assign N1298 = N1297 | data_masked[971];
  assign N1297 = N1296 | data_masked[1510];
  assign N1296 = data_masked[2588] | data_masked[2049];
  assign data_o[433] = N1301 | data_masked[433];
  assign N1301 = N1300 | data_masked[972];
  assign N1300 = N1299 | data_masked[1511];
  assign N1299 = data_masked[2589] | data_masked[2050];
  assign data_o[434] = N1304 | data_masked[434];
  assign N1304 = N1303 | data_masked[973];
  assign N1303 = N1302 | data_masked[1512];
  assign N1302 = data_masked[2590] | data_masked[2051];
  assign data_o[435] = N1307 | data_masked[435];
  assign N1307 = N1306 | data_masked[974];
  assign N1306 = N1305 | data_masked[1513];
  assign N1305 = data_masked[2591] | data_masked[2052];
  assign data_o[436] = N1310 | data_masked[436];
  assign N1310 = N1309 | data_masked[975];
  assign N1309 = N1308 | data_masked[1514];
  assign N1308 = data_masked[2592] | data_masked[2053];
  assign data_o[437] = N1313 | data_masked[437];
  assign N1313 = N1312 | data_masked[976];
  assign N1312 = N1311 | data_masked[1515];
  assign N1311 = data_masked[2593] | data_masked[2054];
  assign data_o[438] = N1316 | data_masked[438];
  assign N1316 = N1315 | data_masked[977];
  assign N1315 = N1314 | data_masked[1516];
  assign N1314 = data_masked[2594] | data_masked[2055];
  assign data_o[439] = N1319 | data_masked[439];
  assign N1319 = N1318 | data_masked[978];
  assign N1318 = N1317 | data_masked[1517];
  assign N1317 = data_masked[2595] | data_masked[2056];
  assign data_o[440] = N1322 | data_masked[440];
  assign N1322 = N1321 | data_masked[979];
  assign N1321 = N1320 | data_masked[1518];
  assign N1320 = data_masked[2596] | data_masked[2057];
  assign data_o[441] = N1325 | data_masked[441];
  assign N1325 = N1324 | data_masked[980];
  assign N1324 = N1323 | data_masked[1519];
  assign N1323 = data_masked[2597] | data_masked[2058];
  assign data_o[442] = N1328 | data_masked[442];
  assign N1328 = N1327 | data_masked[981];
  assign N1327 = N1326 | data_masked[1520];
  assign N1326 = data_masked[2598] | data_masked[2059];
  assign data_o[443] = N1331 | data_masked[443];
  assign N1331 = N1330 | data_masked[982];
  assign N1330 = N1329 | data_masked[1521];
  assign N1329 = data_masked[2599] | data_masked[2060];
  assign data_o[444] = N1334 | data_masked[444];
  assign N1334 = N1333 | data_masked[983];
  assign N1333 = N1332 | data_masked[1522];
  assign N1332 = data_masked[2600] | data_masked[2061];
  assign data_o[445] = N1337 | data_masked[445];
  assign N1337 = N1336 | data_masked[984];
  assign N1336 = N1335 | data_masked[1523];
  assign N1335 = data_masked[2601] | data_masked[2062];
  assign data_o[446] = N1340 | data_masked[446];
  assign N1340 = N1339 | data_masked[985];
  assign N1339 = N1338 | data_masked[1524];
  assign N1338 = data_masked[2602] | data_masked[2063];
  assign data_o[447] = N1343 | data_masked[447];
  assign N1343 = N1342 | data_masked[986];
  assign N1342 = N1341 | data_masked[1525];
  assign N1341 = data_masked[2603] | data_masked[2064];
  assign data_o[448] = N1346 | data_masked[448];
  assign N1346 = N1345 | data_masked[987];
  assign N1345 = N1344 | data_masked[1526];
  assign N1344 = data_masked[2604] | data_masked[2065];
  assign data_o[449] = N1349 | data_masked[449];
  assign N1349 = N1348 | data_masked[988];
  assign N1348 = N1347 | data_masked[1527];
  assign N1347 = data_masked[2605] | data_masked[2066];
  assign data_o[450] = N1352 | data_masked[450];
  assign N1352 = N1351 | data_masked[989];
  assign N1351 = N1350 | data_masked[1528];
  assign N1350 = data_masked[2606] | data_masked[2067];
  assign data_o[451] = N1355 | data_masked[451];
  assign N1355 = N1354 | data_masked[990];
  assign N1354 = N1353 | data_masked[1529];
  assign N1353 = data_masked[2607] | data_masked[2068];
  assign data_o[452] = N1358 | data_masked[452];
  assign N1358 = N1357 | data_masked[991];
  assign N1357 = N1356 | data_masked[1530];
  assign N1356 = data_masked[2608] | data_masked[2069];
  assign data_o[453] = N1361 | data_masked[453];
  assign N1361 = N1360 | data_masked[992];
  assign N1360 = N1359 | data_masked[1531];
  assign N1359 = data_masked[2609] | data_masked[2070];
  assign data_o[454] = N1364 | data_masked[454];
  assign N1364 = N1363 | data_masked[993];
  assign N1363 = N1362 | data_masked[1532];
  assign N1362 = data_masked[2610] | data_masked[2071];
  assign data_o[455] = N1367 | data_masked[455];
  assign N1367 = N1366 | data_masked[994];
  assign N1366 = N1365 | data_masked[1533];
  assign N1365 = data_masked[2611] | data_masked[2072];
  assign data_o[456] = N1370 | data_masked[456];
  assign N1370 = N1369 | data_masked[995];
  assign N1369 = N1368 | data_masked[1534];
  assign N1368 = data_masked[2612] | data_masked[2073];
  assign data_o[457] = N1373 | data_masked[457];
  assign N1373 = N1372 | data_masked[996];
  assign N1372 = N1371 | data_masked[1535];
  assign N1371 = data_masked[2613] | data_masked[2074];
  assign data_o[458] = N1376 | data_masked[458];
  assign N1376 = N1375 | data_masked[997];
  assign N1375 = N1374 | data_masked[1536];
  assign N1374 = data_masked[2614] | data_masked[2075];
  assign data_o[459] = N1379 | data_masked[459];
  assign N1379 = N1378 | data_masked[998];
  assign N1378 = N1377 | data_masked[1537];
  assign N1377 = data_masked[2615] | data_masked[2076];
  assign data_o[460] = N1382 | data_masked[460];
  assign N1382 = N1381 | data_masked[999];
  assign N1381 = N1380 | data_masked[1538];
  assign N1380 = data_masked[2616] | data_masked[2077];
  assign data_o[461] = N1385 | data_masked[461];
  assign N1385 = N1384 | data_masked[1000];
  assign N1384 = N1383 | data_masked[1539];
  assign N1383 = data_masked[2617] | data_masked[2078];
  assign data_o[462] = N1388 | data_masked[462];
  assign N1388 = N1387 | data_masked[1001];
  assign N1387 = N1386 | data_masked[1540];
  assign N1386 = data_masked[2618] | data_masked[2079];
  assign data_o[463] = N1391 | data_masked[463];
  assign N1391 = N1390 | data_masked[1002];
  assign N1390 = N1389 | data_masked[1541];
  assign N1389 = data_masked[2619] | data_masked[2080];
  assign data_o[464] = N1394 | data_masked[464];
  assign N1394 = N1393 | data_masked[1003];
  assign N1393 = N1392 | data_masked[1542];
  assign N1392 = data_masked[2620] | data_masked[2081];
  assign data_o[465] = N1397 | data_masked[465];
  assign N1397 = N1396 | data_masked[1004];
  assign N1396 = N1395 | data_masked[1543];
  assign N1395 = data_masked[2621] | data_masked[2082];
  assign data_o[466] = N1400 | data_masked[466];
  assign N1400 = N1399 | data_masked[1005];
  assign N1399 = N1398 | data_masked[1544];
  assign N1398 = data_masked[2622] | data_masked[2083];
  assign data_o[467] = N1403 | data_masked[467];
  assign N1403 = N1402 | data_masked[1006];
  assign N1402 = N1401 | data_masked[1545];
  assign N1401 = data_masked[2623] | data_masked[2084];
  assign data_o[468] = N1406 | data_masked[468];
  assign N1406 = N1405 | data_masked[1007];
  assign N1405 = N1404 | data_masked[1546];
  assign N1404 = data_masked[2624] | data_masked[2085];
  assign data_o[469] = N1409 | data_masked[469];
  assign N1409 = N1408 | data_masked[1008];
  assign N1408 = N1407 | data_masked[1547];
  assign N1407 = data_masked[2625] | data_masked[2086];
  assign data_o[470] = N1412 | data_masked[470];
  assign N1412 = N1411 | data_masked[1009];
  assign N1411 = N1410 | data_masked[1548];
  assign N1410 = data_masked[2626] | data_masked[2087];
  assign data_o[471] = N1415 | data_masked[471];
  assign N1415 = N1414 | data_masked[1010];
  assign N1414 = N1413 | data_masked[1549];
  assign N1413 = data_masked[2627] | data_masked[2088];
  assign data_o[472] = N1418 | data_masked[472];
  assign N1418 = N1417 | data_masked[1011];
  assign N1417 = N1416 | data_masked[1550];
  assign N1416 = data_masked[2628] | data_masked[2089];
  assign data_o[473] = N1421 | data_masked[473];
  assign N1421 = N1420 | data_masked[1012];
  assign N1420 = N1419 | data_masked[1551];
  assign N1419 = data_masked[2629] | data_masked[2090];
  assign data_o[474] = N1424 | data_masked[474];
  assign N1424 = N1423 | data_masked[1013];
  assign N1423 = N1422 | data_masked[1552];
  assign N1422 = data_masked[2630] | data_masked[2091];
  assign data_o[475] = N1427 | data_masked[475];
  assign N1427 = N1426 | data_masked[1014];
  assign N1426 = N1425 | data_masked[1553];
  assign N1425 = data_masked[2631] | data_masked[2092];
  assign data_o[476] = N1430 | data_masked[476];
  assign N1430 = N1429 | data_masked[1015];
  assign N1429 = N1428 | data_masked[1554];
  assign N1428 = data_masked[2632] | data_masked[2093];
  assign data_o[477] = N1433 | data_masked[477];
  assign N1433 = N1432 | data_masked[1016];
  assign N1432 = N1431 | data_masked[1555];
  assign N1431 = data_masked[2633] | data_masked[2094];
  assign data_o[478] = N1436 | data_masked[478];
  assign N1436 = N1435 | data_masked[1017];
  assign N1435 = N1434 | data_masked[1556];
  assign N1434 = data_masked[2634] | data_masked[2095];
  assign data_o[479] = N1439 | data_masked[479];
  assign N1439 = N1438 | data_masked[1018];
  assign N1438 = N1437 | data_masked[1557];
  assign N1437 = data_masked[2635] | data_masked[2096];
  assign data_o[480] = N1442 | data_masked[480];
  assign N1442 = N1441 | data_masked[1019];
  assign N1441 = N1440 | data_masked[1558];
  assign N1440 = data_masked[2636] | data_masked[2097];
  assign data_o[481] = N1445 | data_masked[481];
  assign N1445 = N1444 | data_masked[1020];
  assign N1444 = N1443 | data_masked[1559];
  assign N1443 = data_masked[2637] | data_masked[2098];
  assign data_o[482] = N1448 | data_masked[482];
  assign N1448 = N1447 | data_masked[1021];
  assign N1447 = N1446 | data_masked[1560];
  assign N1446 = data_masked[2638] | data_masked[2099];
  assign data_o[483] = N1451 | data_masked[483];
  assign N1451 = N1450 | data_masked[1022];
  assign N1450 = N1449 | data_masked[1561];
  assign N1449 = data_masked[2639] | data_masked[2100];
  assign data_o[484] = N1454 | data_masked[484];
  assign N1454 = N1453 | data_masked[1023];
  assign N1453 = N1452 | data_masked[1562];
  assign N1452 = data_masked[2640] | data_masked[2101];
  assign data_o[485] = N1457 | data_masked[485];
  assign N1457 = N1456 | data_masked[1024];
  assign N1456 = N1455 | data_masked[1563];
  assign N1455 = data_masked[2641] | data_masked[2102];
  assign data_o[486] = N1460 | data_masked[486];
  assign N1460 = N1459 | data_masked[1025];
  assign N1459 = N1458 | data_masked[1564];
  assign N1458 = data_masked[2642] | data_masked[2103];
  assign data_o[487] = N1463 | data_masked[487];
  assign N1463 = N1462 | data_masked[1026];
  assign N1462 = N1461 | data_masked[1565];
  assign N1461 = data_masked[2643] | data_masked[2104];
  assign data_o[488] = N1466 | data_masked[488];
  assign N1466 = N1465 | data_masked[1027];
  assign N1465 = N1464 | data_masked[1566];
  assign N1464 = data_masked[2644] | data_masked[2105];
  assign data_o[489] = N1469 | data_masked[489];
  assign N1469 = N1468 | data_masked[1028];
  assign N1468 = N1467 | data_masked[1567];
  assign N1467 = data_masked[2645] | data_masked[2106];
  assign data_o[490] = N1472 | data_masked[490];
  assign N1472 = N1471 | data_masked[1029];
  assign N1471 = N1470 | data_masked[1568];
  assign N1470 = data_masked[2646] | data_masked[2107];
  assign data_o[491] = N1475 | data_masked[491];
  assign N1475 = N1474 | data_masked[1030];
  assign N1474 = N1473 | data_masked[1569];
  assign N1473 = data_masked[2647] | data_masked[2108];
  assign data_o[492] = N1478 | data_masked[492];
  assign N1478 = N1477 | data_masked[1031];
  assign N1477 = N1476 | data_masked[1570];
  assign N1476 = data_masked[2648] | data_masked[2109];
  assign data_o[493] = N1481 | data_masked[493];
  assign N1481 = N1480 | data_masked[1032];
  assign N1480 = N1479 | data_masked[1571];
  assign N1479 = data_masked[2649] | data_masked[2110];
  assign data_o[494] = N1484 | data_masked[494];
  assign N1484 = N1483 | data_masked[1033];
  assign N1483 = N1482 | data_masked[1572];
  assign N1482 = data_masked[2650] | data_masked[2111];
  assign data_o[495] = N1487 | data_masked[495];
  assign N1487 = N1486 | data_masked[1034];
  assign N1486 = N1485 | data_masked[1573];
  assign N1485 = data_masked[2651] | data_masked[2112];
  assign data_o[496] = N1490 | data_masked[496];
  assign N1490 = N1489 | data_masked[1035];
  assign N1489 = N1488 | data_masked[1574];
  assign N1488 = data_masked[2652] | data_masked[2113];
  assign data_o[497] = N1493 | data_masked[497];
  assign N1493 = N1492 | data_masked[1036];
  assign N1492 = N1491 | data_masked[1575];
  assign N1491 = data_masked[2653] | data_masked[2114];
  assign data_o[498] = N1496 | data_masked[498];
  assign N1496 = N1495 | data_masked[1037];
  assign N1495 = N1494 | data_masked[1576];
  assign N1494 = data_masked[2654] | data_masked[2115];
  assign data_o[499] = N1499 | data_masked[499];
  assign N1499 = N1498 | data_masked[1038];
  assign N1498 = N1497 | data_masked[1577];
  assign N1497 = data_masked[2655] | data_masked[2116];
  assign data_o[500] = N1502 | data_masked[500];
  assign N1502 = N1501 | data_masked[1039];
  assign N1501 = N1500 | data_masked[1578];
  assign N1500 = data_masked[2656] | data_masked[2117];
  assign data_o[501] = N1505 | data_masked[501];
  assign N1505 = N1504 | data_masked[1040];
  assign N1504 = N1503 | data_masked[1579];
  assign N1503 = data_masked[2657] | data_masked[2118];
  assign data_o[502] = N1508 | data_masked[502];
  assign N1508 = N1507 | data_masked[1041];
  assign N1507 = N1506 | data_masked[1580];
  assign N1506 = data_masked[2658] | data_masked[2119];
  assign data_o[503] = N1511 | data_masked[503];
  assign N1511 = N1510 | data_masked[1042];
  assign N1510 = N1509 | data_masked[1581];
  assign N1509 = data_masked[2659] | data_masked[2120];
  assign data_o[504] = N1514 | data_masked[504];
  assign N1514 = N1513 | data_masked[1043];
  assign N1513 = N1512 | data_masked[1582];
  assign N1512 = data_masked[2660] | data_masked[2121];
  assign data_o[505] = N1517 | data_masked[505];
  assign N1517 = N1516 | data_masked[1044];
  assign N1516 = N1515 | data_masked[1583];
  assign N1515 = data_masked[2661] | data_masked[2122];
  assign data_o[506] = N1520 | data_masked[506];
  assign N1520 = N1519 | data_masked[1045];
  assign N1519 = N1518 | data_masked[1584];
  assign N1518 = data_masked[2662] | data_masked[2123];
  assign data_o[507] = N1523 | data_masked[507];
  assign N1523 = N1522 | data_masked[1046];
  assign N1522 = N1521 | data_masked[1585];
  assign N1521 = data_masked[2663] | data_masked[2124];
  assign data_o[508] = N1526 | data_masked[508];
  assign N1526 = N1525 | data_masked[1047];
  assign N1525 = N1524 | data_masked[1586];
  assign N1524 = data_masked[2664] | data_masked[2125];
  assign data_o[509] = N1529 | data_masked[509];
  assign N1529 = N1528 | data_masked[1048];
  assign N1528 = N1527 | data_masked[1587];
  assign N1527 = data_masked[2665] | data_masked[2126];
  assign data_o[510] = N1532 | data_masked[510];
  assign N1532 = N1531 | data_masked[1049];
  assign N1531 = N1530 | data_masked[1588];
  assign N1530 = data_masked[2666] | data_masked[2127];
  assign data_o[511] = N1535 | data_masked[511];
  assign N1535 = N1534 | data_masked[1050];
  assign N1534 = N1533 | data_masked[1589];
  assign N1533 = data_masked[2667] | data_masked[2128];
  assign data_o[512] = N1538 | data_masked[512];
  assign N1538 = N1537 | data_masked[1051];
  assign N1537 = N1536 | data_masked[1590];
  assign N1536 = data_masked[2668] | data_masked[2129];
  assign data_o[513] = N1541 | data_masked[513];
  assign N1541 = N1540 | data_masked[1052];
  assign N1540 = N1539 | data_masked[1591];
  assign N1539 = data_masked[2669] | data_masked[2130];
  assign data_o[514] = N1544 | data_masked[514];
  assign N1544 = N1543 | data_masked[1053];
  assign N1543 = N1542 | data_masked[1592];
  assign N1542 = data_masked[2670] | data_masked[2131];
  assign data_o[515] = N1547 | data_masked[515];
  assign N1547 = N1546 | data_masked[1054];
  assign N1546 = N1545 | data_masked[1593];
  assign N1545 = data_masked[2671] | data_masked[2132];
  assign data_o[516] = N1550 | data_masked[516];
  assign N1550 = N1549 | data_masked[1055];
  assign N1549 = N1548 | data_masked[1594];
  assign N1548 = data_masked[2672] | data_masked[2133];
  assign data_o[517] = N1553 | data_masked[517];
  assign N1553 = N1552 | data_masked[1056];
  assign N1552 = N1551 | data_masked[1595];
  assign N1551 = data_masked[2673] | data_masked[2134];
  assign data_o[518] = N1556 | data_masked[518];
  assign N1556 = N1555 | data_masked[1057];
  assign N1555 = N1554 | data_masked[1596];
  assign N1554 = data_masked[2674] | data_masked[2135];
  assign data_o[519] = N1559 | data_masked[519];
  assign N1559 = N1558 | data_masked[1058];
  assign N1558 = N1557 | data_masked[1597];
  assign N1557 = data_masked[2675] | data_masked[2136];
  assign data_o[520] = N1562 | data_masked[520];
  assign N1562 = N1561 | data_masked[1059];
  assign N1561 = N1560 | data_masked[1598];
  assign N1560 = data_masked[2676] | data_masked[2137];
  assign data_o[521] = N1565 | data_masked[521];
  assign N1565 = N1564 | data_masked[1060];
  assign N1564 = N1563 | data_masked[1599];
  assign N1563 = data_masked[2677] | data_masked[2138];
  assign data_o[522] = N1568 | data_masked[522];
  assign N1568 = N1567 | data_masked[1061];
  assign N1567 = N1566 | data_masked[1600];
  assign N1566 = data_masked[2678] | data_masked[2139];
  assign data_o[523] = N1571 | data_masked[523];
  assign N1571 = N1570 | data_masked[1062];
  assign N1570 = N1569 | data_masked[1601];
  assign N1569 = data_masked[2679] | data_masked[2140];
  assign data_o[524] = N1574 | data_masked[524];
  assign N1574 = N1573 | data_masked[1063];
  assign N1573 = N1572 | data_masked[1602];
  assign N1572 = data_masked[2680] | data_masked[2141];
  assign data_o[525] = N1577 | data_masked[525];
  assign N1577 = N1576 | data_masked[1064];
  assign N1576 = N1575 | data_masked[1603];
  assign N1575 = data_masked[2681] | data_masked[2142];
  assign data_o[526] = N1580 | data_masked[526];
  assign N1580 = N1579 | data_masked[1065];
  assign N1579 = N1578 | data_masked[1604];
  assign N1578 = data_masked[2682] | data_masked[2143];
  assign data_o[527] = N1583 | data_masked[527];
  assign N1583 = N1582 | data_masked[1066];
  assign N1582 = N1581 | data_masked[1605];
  assign N1581 = data_masked[2683] | data_masked[2144];
  assign data_o[528] = N1586 | data_masked[528];
  assign N1586 = N1585 | data_masked[1067];
  assign N1585 = N1584 | data_masked[1606];
  assign N1584 = data_masked[2684] | data_masked[2145];
  assign data_o[529] = N1589 | data_masked[529];
  assign N1589 = N1588 | data_masked[1068];
  assign N1588 = N1587 | data_masked[1607];
  assign N1587 = data_masked[2685] | data_masked[2146];
  assign data_o[530] = N1592 | data_masked[530];
  assign N1592 = N1591 | data_masked[1069];
  assign N1591 = N1590 | data_masked[1608];
  assign N1590 = data_masked[2686] | data_masked[2147];
  assign data_o[531] = N1595 | data_masked[531];
  assign N1595 = N1594 | data_masked[1070];
  assign N1594 = N1593 | data_masked[1609];
  assign N1593 = data_masked[2687] | data_masked[2148];
  assign data_o[532] = N1598 | data_masked[532];
  assign N1598 = N1597 | data_masked[1071];
  assign N1597 = N1596 | data_masked[1610];
  assign N1596 = data_masked[2688] | data_masked[2149];
  assign data_o[533] = N1601 | data_masked[533];
  assign N1601 = N1600 | data_masked[1072];
  assign N1600 = N1599 | data_masked[1611];
  assign N1599 = data_masked[2689] | data_masked[2150];
  assign data_o[534] = N1604 | data_masked[534];
  assign N1604 = N1603 | data_masked[1073];
  assign N1603 = N1602 | data_masked[1612];
  assign N1602 = data_masked[2690] | data_masked[2151];
  assign data_o[535] = N1607 | data_masked[535];
  assign N1607 = N1606 | data_masked[1074];
  assign N1606 = N1605 | data_masked[1613];
  assign N1605 = data_masked[2691] | data_masked[2152];
  assign data_o[536] = N1610 | data_masked[536];
  assign N1610 = N1609 | data_masked[1075];
  assign N1609 = N1608 | data_masked[1614];
  assign N1608 = data_masked[2692] | data_masked[2153];
  assign data_o[537] = N1613 | data_masked[537];
  assign N1613 = N1612 | data_masked[1076];
  assign N1612 = N1611 | data_masked[1615];
  assign N1611 = data_masked[2693] | data_masked[2154];
  assign data_o[538] = N1616 | data_masked[538];
  assign N1616 = N1615 | data_masked[1077];
  assign N1615 = N1614 | data_masked[1616];
  assign N1614 = data_masked[2694] | data_masked[2155];

endmodule