module bsg_mem_1rw_sync_mask_write_bit_synth_width_p15_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [14:0] data_i;
  input [5:0] addr_i;
  input [14:0] w_mask_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [14:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290;
  wire [5:0] addr_r;
  wire [959:0] mem;
  reg addr_r_5_sv2v_reg,addr_r_4_sv2v_reg,addr_r_3_sv2v_reg,addr_r_2_sv2v_reg,
  addr_r_1_sv2v_reg,addr_r_0_sv2v_reg,mem_959_sv2v_reg,mem_958_sv2v_reg,mem_957_sv2v_reg,
  mem_956_sv2v_reg,mem_955_sv2v_reg,mem_954_sv2v_reg,mem_953_sv2v_reg,
  mem_952_sv2v_reg,mem_951_sv2v_reg,mem_950_sv2v_reg,mem_949_sv2v_reg,mem_948_sv2v_reg,
  mem_947_sv2v_reg,mem_946_sv2v_reg,mem_945_sv2v_reg,mem_944_sv2v_reg,mem_943_sv2v_reg,
  mem_942_sv2v_reg,mem_941_sv2v_reg,mem_940_sv2v_reg,mem_939_sv2v_reg,
  mem_938_sv2v_reg,mem_937_sv2v_reg,mem_936_sv2v_reg,mem_935_sv2v_reg,mem_934_sv2v_reg,
  mem_933_sv2v_reg,mem_932_sv2v_reg,mem_931_sv2v_reg,mem_930_sv2v_reg,mem_929_sv2v_reg,
  mem_928_sv2v_reg,mem_927_sv2v_reg,mem_926_sv2v_reg,mem_925_sv2v_reg,mem_924_sv2v_reg,
  mem_923_sv2v_reg,mem_922_sv2v_reg,mem_921_sv2v_reg,mem_920_sv2v_reg,
  mem_919_sv2v_reg,mem_918_sv2v_reg,mem_917_sv2v_reg,mem_916_sv2v_reg,mem_915_sv2v_reg,
  mem_914_sv2v_reg,mem_913_sv2v_reg,mem_912_sv2v_reg,mem_911_sv2v_reg,mem_910_sv2v_reg,
  mem_909_sv2v_reg,mem_908_sv2v_reg,mem_907_sv2v_reg,mem_906_sv2v_reg,
  mem_905_sv2v_reg,mem_904_sv2v_reg,mem_903_sv2v_reg,mem_902_sv2v_reg,mem_901_sv2v_reg,
  mem_900_sv2v_reg,mem_899_sv2v_reg,mem_898_sv2v_reg,mem_897_sv2v_reg,mem_896_sv2v_reg,
  mem_895_sv2v_reg,mem_894_sv2v_reg,mem_893_sv2v_reg,mem_892_sv2v_reg,
  mem_891_sv2v_reg,mem_890_sv2v_reg,mem_889_sv2v_reg,mem_888_sv2v_reg,mem_887_sv2v_reg,
  mem_886_sv2v_reg,mem_885_sv2v_reg,mem_884_sv2v_reg,mem_883_sv2v_reg,mem_882_sv2v_reg,
  mem_881_sv2v_reg,mem_880_sv2v_reg,mem_879_sv2v_reg,mem_878_sv2v_reg,mem_877_sv2v_reg,
  mem_876_sv2v_reg,mem_875_sv2v_reg,mem_874_sv2v_reg,mem_873_sv2v_reg,
  mem_872_sv2v_reg,mem_871_sv2v_reg,mem_870_sv2v_reg,mem_869_sv2v_reg,mem_868_sv2v_reg,
  mem_867_sv2v_reg,mem_866_sv2v_reg,mem_865_sv2v_reg,mem_864_sv2v_reg,mem_863_sv2v_reg,
  mem_862_sv2v_reg,mem_861_sv2v_reg,mem_860_sv2v_reg,mem_859_sv2v_reg,
  mem_858_sv2v_reg,mem_857_sv2v_reg,mem_856_sv2v_reg,mem_855_sv2v_reg,mem_854_sv2v_reg,
  mem_853_sv2v_reg,mem_852_sv2v_reg,mem_851_sv2v_reg,mem_850_sv2v_reg,mem_849_sv2v_reg,
  mem_848_sv2v_reg,mem_847_sv2v_reg,mem_846_sv2v_reg,mem_845_sv2v_reg,mem_844_sv2v_reg,
  mem_843_sv2v_reg,mem_842_sv2v_reg,mem_841_sv2v_reg,mem_840_sv2v_reg,
  mem_839_sv2v_reg,mem_838_sv2v_reg,mem_837_sv2v_reg,mem_836_sv2v_reg,mem_835_sv2v_reg,
  mem_834_sv2v_reg,mem_833_sv2v_reg,mem_832_sv2v_reg,mem_831_sv2v_reg,mem_830_sv2v_reg,
  mem_829_sv2v_reg,mem_828_sv2v_reg,mem_827_sv2v_reg,mem_826_sv2v_reg,
  mem_825_sv2v_reg,mem_824_sv2v_reg,mem_823_sv2v_reg,mem_822_sv2v_reg,mem_821_sv2v_reg,
  mem_820_sv2v_reg,mem_819_sv2v_reg,mem_818_sv2v_reg,mem_817_sv2v_reg,mem_816_sv2v_reg,
  mem_815_sv2v_reg,mem_814_sv2v_reg,mem_813_sv2v_reg,mem_812_sv2v_reg,
  mem_811_sv2v_reg,mem_810_sv2v_reg,mem_809_sv2v_reg,mem_808_sv2v_reg,mem_807_sv2v_reg,
  mem_806_sv2v_reg,mem_805_sv2v_reg,mem_804_sv2v_reg,mem_803_sv2v_reg,mem_802_sv2v_reg,
  mem_801_sv2v_reg,mem_800_sv2v_reg,mem_799_sv2v_reg,mem_798_sv2v_reg,mem_797_sv2v_reg,
  mem_796_sv2v_reg,mem_795_sv2v_reg,mem_794_sv2v_reg,mem_793_sv2v_reg,
  mem_792_sv2v_reg,mem_791_sv2v_reg,mem_790_sv2v_reg,mem_789_sv2v_reg,mem_788_sv2v_reg,
  mem_787_sv2v_reg,mem_786_sv2v_reg,mem_785_sv2v_reg,mem_784_sv2v_reg,mem_783_sv2v_reg,
  mem_782_sv2v_reg,mem_781_sv2v_reg,mem_780_sv2v_reg,mem_779_sv2v_reg,
  mem_778_sv2v_reg,mem_777_sv2v_reg,mem_776_sv2v_reg,mem_775_sv2v_reg,mem_774_sv2v_reg,
  mem_773_sv2v_reg,mem_772_sv2v_reg,mem_771_sv2v_reg,mem_770_sv2v_reg,mem_769_sv2v_reg,
  mem_768_sv2v_reg,mem_767_sv2v_reg,mem_766_sv2v_reg,mem_765_sv2v_reg,mem_764_sv2v_reg,
  mem_763_sv2v_reg,mem_762_sv2v_reg,mem_761_sv2v_reg,mem_760_sv2v_reg,
  mem_759_sv2v_reg,mem_758_sv2v_reg,mem_757_sv2v_reg,mem_756_sv2v_reg,mem_755_sv2v_reg,
  mem_754_sv2v_reg,mem_753_sv2v_reg,mem_752_sv2v_reg,mem_751_sv2v_reg,mem_750_sv2v_reg,
  mem_749_sv2v_reg,mem_748_sv2v_reg,mem_747_sv2v_reg,mem_746_sv2v_reg,
  mem_745_sv2v_reg,mem_744_sv2v_reg,mem_743_sv2v_reg,mem_742_sv2v_reg,mem_741_sv2v_reg,
  mem_740_sv2v_reg,mem_739_sv2v_reg,mem_738_sv2v_reg,mem_737_sv2v_reg,mem_736_sv2v_reg,
  mem_735_sv2v_reg,mem_734_sv2v_reg,mem_733_sv2v_reg,mem_732_sv2v_reg,
  mem_731_sv2v_reg,mem_730_sv2v_reg,mem_729_sv2v_reg,mem_728_sv2v_reg,mem_727_sv2v_reg,
  mem_726_sv2v_reg,mem_725_sv2v_reg,mem_724_sv2v_reg,mem_723_sv2v_reg,mem_722_sv2v_reg,
  mem_721_sv2v_reg,mem_720_sv2v_reg,mem_719_sv2v_reg,mem_718_sv2v_reg,mem_717_sv2v_reg,
  mem_716_sv2v_reg,mem_715_sv2v_reg,mem_714_sv2v_reg,mem_713_sv2v_reg,
  mem_712_sv2v_reg,mem_711_sv2v_reg,mem_710_sv2v_reg,mem_709_sv2v_reg,mem_708_sv2v_reg,
  mem_707_sv2v_reg,mem_706_sv2v_reg,mem_705_sv2v_reg,mem_704_sv2v_reg,mem_703_sv2v_reg,
  mem_702_sv2v_reg,mem_701_sv2v_reg,mem_700_sv2v_reg,mem_699_sv2v_reg,
  mem_698_sv2v_reg,mem_697_sv2v_reg,mem_696_sv2v_reg,mem_695_sv2v_reg,mem_694_sv2v_reg,
  mem_693_sv2v_reg,mem_692_sv2v_reg,mem_691_sv2v_reg,mem_690_sv2v_reg,mem_689_sv2v_reg,
  mem_688_sv2v_reg,mem_687_sv2v_reg,mem_686_sv2v_reg,mem_685_sv2v_reg,mem_684_sv2v_reg,
  mem_683_sv2v_reg,mem_682_sv2v_reg,mem_681_sv2v_reg,mem_680_sv2v_reg,
  mem_679_sv2v_reg,mem_678_sv2v_reg,mem_677_sv2v_reg,mem_676_sv2v_reg,mem_675_sv2v_reg,
  mem_674_sv2v_reg,mem_673_sv2v_reg,mem_672_sv2v_reg,mem_671_sv2v_reg,mem_670_sv2v_reg,
  mem_669_sv2v_reg,mem_668_sv2v_reg,mem_667_sv2v_reg,mem_666_sv2v_reg,
  mem_665_sv2v_reg,mem_664_sv2v_reg,mem_663_sv2v_reg,mem_662_sv2v_reg,mem_661_sv2v_reg,
  mem_660_sv2v_reg,mem_659_sv2v_reg,mem_658_sv2v_reg,mem_657_sv2v_reg,mem_656_sv2v_reg,
  mem_655_sv2v_reg,mem_654_sv2v_reg,mem_653_sv2v_reg,mem_652_sv2v_reg,
  mem_651_sv2v_reg,mem_650_sv2v_reg,mem_649_sv2v_reg,mem_648_sv2v_reg,mem_647_sv2v_reg,
  mem_646_sv2v_reg,mem_645_sv2v_reg,mem_644_sv2v_reg,mem_643_sv2v_reg,mem_642_sv2v_reg,
  mem_641_sv2v_reg,mem_640_sv2v_reg,mem_639_sv2v_reg,mem_638_sv2v_reg,mem_637_sv2v_reg,
  mem_636_sv2v_reg,mem_635_sv2v_reg,mem_634_sv2v_reg,mem_633_sv2v_reg,
  mem_632_sv2v_reg,mem_631_sv2v_reg,mem_630_sv2v_reg,mem_629_sv2v_reg,mem_628_sv2v_reg,
  mem_627_sv2v_reg,mem_626_sv2v_reg,mem_625_sv2v_reg,mem_624_sv2v_reg,mem_623_sv2v_reg,
  mem_622_sv2v_reg,mem_621_sv2v_reg,mem_620_sv2v_reg,mem_619_sv2v_reg,
  mem_618_sv2v_reg,mem_617_sv2v_reg,mem_616_sv2v_reg,mem_615_sv2v_reg,mem_614_sv2v_reg,
  mem_613_sv2v_reg,mem_612_sv2v_reg,mem_611_sv2v_reg,mem_610_sv2v_reg,mem_609_sv2v_reg,
  mem_608_sv2v_reg,mem_607_sv2v_reg,mem_606_sv2v_reg,mem_605_sv2v_reg,mem_604_sv2v_reg,
  mem_603_sv2v_reg,mem_602_sv2v_reg,mem_601_sv2v_reg,mem_600_sv2v_reg,
  mem_599_sv2v_reg,mem_598_sv2v_reg,mem_597_sv2v_reg,mem_596_sv2v_reg,mem_595_sv2v_reg,
  mem_594_sv2v_reg,mem_593_sv2v_reg,mem_592_sv2v_reg,mem_591_sv2v_reg,mem_590_sv2v_reg,
  mem_589_sv2v_reg,mem_588_sv2v_reg,mem_587_sv2v_reg,mem_586_sv2v_reg,
  mem_585_sv2v_reg,mem_584_sv2v_reg,mem_583_sv2v_reg,mem_582_sv2v_reg,mem_581_sv2v_reg,
  mem_580_sv2v_reg,mem_579_sv2v_reg,mem_578_sv2v_reg,mem_577_sv2v_reg,mem_576_sv2v_reg,
  mem_575_sv2v_reg,mem_574_sv2v_reg,mem_573_sv2v_reg,mem_572_sv2v_reg,
  mem_571_sv2v_reg,mem_570_sv2v_reg,mem_569_sv2v_reg,mem_568_sv2v_reg,mem_567_sv2v_reg,
  mem_566_sv2v_reg,mem_565_sv2v_reg,mem_564_sv2v_reg,mem_563_sv2v_reg,mem_562_sv2v_reg,
  mem_561_sv2v_reg,mem_560_sv2v_reg,mem_559_sv2v_reg,mem_558_sv2v_reg,mem_557_sv2v_reg,
  mem_556_sv2v_reg,mem_555_sv2v_reg,mem_554_sv2v_reg,mem_553_sv2v_reg,
  mem_552_sv2v_reg,mem_551_sv2v_reg,mem_550_sv2v_reg,mem_549_sv2v_reg,mem_548_sv2v_reg,
  mem_547_sv2v_reg,mem_546_sv2v_reg,mem_545_sv2v_reg,mem_544_sv2v_reg,mem_543_sv2v_reg,
  mem_542_sv2v_reg,mem_541_sv2v_reg,mem_540_sv2v_reg,mem_539_sv2v_reg,
  mem_538_sv2v_reg,mem_537_sv2v_reg,mem_536_sv2v_reg,mem_535_sv2v_reg,mem_534_sv2v_reg,
  mem_533_sv2v_reg,mem_532_sv2v_reg,mem_531_sv2v_reg,mem_530_sv2v_reg,mem_529_sv2v_reg,
  mem_528_sv2v_reg,mem_527_sv2v_reg,mem_526_sv2v_reg,mem_525_sv2v_reg,mem_524_sv2v_reg,
  mem_523_sv2v_reg,mem_522_sv2v_reg,mem_521_sv2v_reg,mem_520_sv2v_reg,
  mem_519_sv2v_reg,mem_518_sv2v_reg,mem_517_sv2v_reg,mem_516_sv2v_reg,mem_515_sv2v_reg,
  mem_514_sv2v_reg,mem_513_sv2v_reg,mem_512_sv2v_reg,mem_511_sv2v_reg,mem_510_sv2v_reg,
  mem_509_sv2v_reg,mem_508_sv2v_reg,mem_507_sv2v_reg,mem_506_sv2v_reg,
  mem_505_sv2v_reg,mem_504_sv2v_reg,mem_503_sv2v_reg,mem_502_sv2v_reg,mem_501_sv2v_reg,
  mem_500_sv2v_reg,mem_499_sv2v_reg,mem_498_sv2v_reg,mem_497_sv2v_reg,mem_496_sv2v_reg,
  mem_495_sv2v_reg,mem_494_sv2v_reg,mem_493_sv2v_reg,mem_492_sv2v_reg,
  mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,mem_488_sv2v_reg,mem_487_sv2v_reg,
  mem_486_sv2v_reg,mem_485_sv2v_reg,mem_484_sv2v_reg,mem_483_sv2v_reg,mem_482_sv2v_reg,
  mem_481_sv2v_reg,mem_480_sv2v_reg,mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,
  mem_476_sv2v_reg,mem_475_sv2v_reg,mem_474_sv2v_reg,mem_473_sv2v_reg,
  mem_472_sv2v_reg,mem_471_sv2v_reg,mem_470_sv2v_reg,mem_469_sv2v_reg,mem_468_sv2v_reg,
  mem_467_sv2v_reg,mem_466_sv2v_reg,mem_465_sv2v_reg,mem_464_sv2v_reg,mem_463_sv2v_reg,
  mem_462_sv2v_reg,mem_461_sv2v_reg,mem_460_sv2v_reg,mem_459_sv2v_reg,
  mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,mem_455_sv2v_reg,mem_454_sv2v_reg,
  mem_453_sv2v_reg,mem_452_sv2v_reg,mem_451_sv2v_reg,mem_450_sv2v_reg,mem_449_sv2v_reg,
  mem_448_sv2v_reg,mem_447_sv2v_reg,mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,
  mem_443_sv2v_reg,mem_442_sv2v_reg,mem_441_sv2v_reg,mem_440_sv2v_reg,
  mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,mem_436_sv2v_reg,mem_435_sv2v_reg,
  mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,mem_431_sv2v_reg,mem_430_sv2v_reg,
  mem_429_sv2v_reg,mem_428_sv2v_reg,mem_427_sv2v_reg,mem_426_sv2v_reg,
  mem_425_sv2v_reg,mem_424_sv2v_reg,mem_423_sv2v_reg,mem_422_sv2v_reg,mem_421_sv2v_reg,
  mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,mem_417_sv2v_reg,mem_416_sv2v_reg,
  mem_415_sv2v_reg,mem_414_sv2v_reg,mem_413_sv2v_reg,mem_412_sv2v_reg,
  mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,mem_408_sv2v_reg,mem_407_sv2v_reg,
  mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,mem_403_sv2v_reg,mem_402_sv2v_reg,
  mem_401_sv2v_reg,mem_400_sv2v_reg,mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,
  mem_396_sv2v_reg,mem_395_sv2v_reg,mem_394_sv2v_reg,mem_393_sv2v_reg,
  mem_392_sv2v_reg,mem_391_sv2v_reg,mem_390_sv2v_reg,mem_389_sv2v_reg,mem_388_sv2v_reg,
  mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,mem_384_sv2v_reg,mem_383_sv2v_reg,
  mem_382_sv2v_reg,mem_381_sv2v_reg,mem_380_sv2v_reg,mem_379_sv2v_reg,
  mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,mem_375_sv2v_reg,mem_374_sv2v_reg,
  mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,mem_370_sv2v_reg,mem_369_sv2v_reg,
  mem_368_sv2v_reg,mem_367_sv2v_reg,mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,
  mem_363_sv2v_reg,mem_362_sv2v_reg,mem_361_sv2v_reg,mem_360_sv2v_reg,
  mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,mem_356_sv2v_reg,mem_355_sv2v_reg,
  mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,mem_351_sv2v_reg,mem_350_sv2v_reg,
  mem_349_sv2v_reg,mem_348_sv2v_reg,mem_347_sv2v_reg,mem_346_sv2v_reg,
  mem_345_sv2v_reg,mem_344_sv2v_reg,mem_343_sv2v_reg,mem_342_sv2v_reg,mem_341_sv2v_reg,
  mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,mem_337_sv2v_reg,mem_336_sv2v_reg,
  mem_335_sv2v_reg,mem_334_sv2v_reg,mem_333_sv2v_reg,mem_332_sv2v_reg,
  mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,mem_328_sv2v_reg,mem_327_sv2v_reg,
  mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,mem_323_sv2v_reg,mem_322_sv2v_reg,
  mem_321_sv2v_reg,mem_320_sv2v_reg,mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,
  mem_316_sv2v_reg,mem_315_sv2v_reg,mem_314_sv2v_reg,mem_313_sv2v_reg,
  mem_312_sv2v_reg,mem_311_sv2v_reg,mem_310_sv2v_reg,mem_309_sv2v_reg,mem_308_sv2v_reg,
  mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,mem_304_sv2v_reg,mem_303_sv2v_reg,
  mem_302_sv2v_reg,mem_301_sv2v_reg,mem_300_sv2v_reg,mem_299_sv2v_reg,
  mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,mem_295_sv2v_reg,mem_294_sv2v_reg,
  mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,mem_290_sv2v_reg,mem_289_sv2v_reg,
  mem_288_sv2v_reg,mem_287_sv2v_reg,mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,
  mem_283_sv2v_reg,mem_282_sv2v_reg,mem_281_sv2v_reg,mem_280_sv2v_reg,
  mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,mem_276_sv2v_reg,mem_275_sv2v_reg,
  mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,mem_271_sv2v_reg,mem_270_sv2v_reg,
  mem_269_sv2v_reg,mem_268_sv2v_reg,mem_267_sv2v_reg,mem_266_sv2v_reg,
  mem_265_sv2v_reg,mem_264_sv2v_reg,mem_263_sv2v_reg,mem_262_sv2v_reg,mem_261_sv2v_reg,
  mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,mem_257_sv2v_reg,mem_256_sv2v_reg,
  mem_255_sv2v_reg,mem_254_sv2v_reg,mem_253_sv2v_reg,mem_252_sv2v_reg,
  mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,mem_248_sv2v_reg,mem_247_sv2v_reg,
  mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,mem_243_sv2v_reg,mem_242_sv2v_reg,
  mem_241_sv2v_reg,mem_240_sv2v_reg,mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,
  mem_236_sv2v_reg,mem_235_sv2v_reg,mem_234_sv2v_reg,mem_233_sv2v_reg,
  mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,mem_229_sv2v_reg,mem_228_sv2v_reg,
  mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,mem_224_sv2v_reg,mem_223_sv2v_reg,
  mem_222_sv2v_reg,mem_221_sv2v_reg,mem_220_sv2v_reg,mem_219_sv2v_reg,
  mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,mem_215_sv2v_reg,mem_214_sv2v_reg,
  mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,mem_210_sv2v_reg,mem_209_sv2v_reg,
  mem_208_sv2v_reg,mem_207_sv2v_reg,mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,
  mem_203_sv2v_reg,mem_202_sv2v_reg,mem_201_sv2v_reg,mem_200_sv2v_reg,
  mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,mem_196_sv2v_reg,mem_195_sv2v_reg,
  mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,mem_191_sv2v_reg,mem_190_sv2v_reg,
  mem_189_sv2v_reg,mem_188_sv2v_reg,mem_187_sv2v_reg,mem_186_sv2v_reg,
  mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,mem_182_sv2v_reg,mem_181_sv2v_reg,
  mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,mem_177_sv2v_reg,mem_176_sv2v_reg,
  mem_175_sv2v_reg,mem_174_sv2v_reg,mem_173_sv2v_reg,mem_172_sv2v_reg,
  mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,mem_168_sv2v_reg,mem_167_sv2v_reg,
  mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,mem_163_sv2v_reg,mem_162_sv2v_reg,
  mem_161_sv2v_reg,mem_160_sv2v_reg,mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,
  mem_156_sv2v_reg,mem_155_sv2v_reg,mem_154_sv2v_reg,mem_153_sv2v_reg,
  mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,mem_149_sv2v_reg,mem_148_sv2v_reg,
  mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,mem_144_sv2v_reg,mem_143_sv2v_reg,
  mem_142_sv2v_reg,mem_141_sv2v_reg,mem_140_sv2v_reg,mem_139_sv2v_reg,
  mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,mem_135_sv2v_reg,mem_134_sv2v_reg,
  mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,mem_130_sv2v_reg,mem_129_sv2v_reg,
  mem_128_sv2v_reg,mem_127_sv2v_reg,mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,
  mem_123_sv2v_reg,mem_122_sv2v_reg,mem_121_sv2v_reg,mem_120_sv2v_reg,
  mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,mem_116_sv2v_reg,mem_115_sv2v_reg,
  mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,mem_111_sv2v_reg,mem_110_sv2v_reg,
  mem_109_sv2v_reg,mem_108_sv2v_reg,mem_107_sv2v_reg,mem_106_sv2v_reg,
  mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,mem_102_sv2v_reg,mem_101_sv2v_reg,
  mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,mem_97_sv2v_reg,mem_96_sv2v_reg,
  mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,mem_92_sv2v_reg,mem_91_sv2v_reg,
  mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,mem_87_sv2v_reg,mem_86_sv2v_reg,
  mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,mem_82_sv2v_reg,mem_81_sv2v_reg,
  mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,mem_77_sv2v_reg,mem_76_sv2v_reg,
  mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,mem_72_sv2v_reg,mem_71_sv2v_reg,
  mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,mem_67_sv2v_reg,mem_66_sv2v_reg,
  mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,
  mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,
  mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,
  mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,
  mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,
  mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,
  mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,
  mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,
  mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,
  mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,
  mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,
  mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,
  mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign addr_r[5] = addr_r_5_sv2v_reg;
  assign addr_r[4] = addr_r_4_sv2v_reg;
  assign addr_r[3] = addr_r_3_sv2v_reg;
  assign addr_r[2] = addr_r_2_sv2v_reg;
  assign addr_r[1] = addr_r_1_sv2v_reg;
  assign addr_r[0] = addr_r_0_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_5_sv2v_reg <= addr_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_4_sv2v_reg <= addr_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_3_sv2v_reg <= addr_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_2_sv2v_reg <= addr_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_1_sv2v_reg <= addr_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_0_sv2v_reg <= addr_i[0];
    end 
  end

  assign data_o[14] = (N90)? mem[14] : 
                      (N92)? mem[29] : 
                      (N94)? mem[44] : 
                      (N96)? mem[59] : 
                      (N98)? mem[74] : 
                      (N100)? mem[89] : 
                      (N102)? mem[104] : 
                      (N104)? mem[119] : 
                      (N106)? mem[134] : 
                      (N108)? mem[149] : 
                      (N110)? mem[164] : 
                      (N112)? mem[179] : 
                      (N114)? mem[194] : 
                      (N116)? mem[209] : 
                      (N118)? mem[224] : 
                      (N120)? mem[239] : 
                      (N122)? mem[254] : 
                      (N124)? mem[269] : 
                      (N126)? mem[284] : 
                      (N128)? mem[299] : 
                      (N130)? mem[314] : 
                      (N132)? mem[329] : 
                      (N134)? mem[344] : 
                      (N136)? mem[359] : 
                      (N138)? mem[374] : 
                      (N140)? mem[389] : 
                      (N142)? mem[404] : 
                      (N144)? mem[419] : 
                      (N146)? mem[434] : 
                      (N148)? mem[449] : 
                      (N150)? mem[464] : 
                      (N152)? mem[479] : 
                      (N91)? mem[494] : 
                      (N93)? mem[509] : 
                      (N95)? mem[524] : 
                      (N97)? mem[539] : 
                      (N99)? mem[554] : 
                      (N101)? mem[569] : 
                      (N103)? mem[584] : 
                      (N105)? mem[599] : 
                      (N107)? mem[614] : 
                      (N109)? mem[629] : 
                      (N111)? mem[644] : 
                      (N113)? mem[659] : 
                      (N115)? mem[674] : 
                      (N117)? mem[689] : 
                      (N119)? mem[704] : 
                      (N121)? mem[719] : 
                      (N123)? mem[734] : 
                      (N125)? mem[749] : 
                      (N127)? mem[764] : 
                      (N129)? mem[779] : 
                      (N131)? mem[794] : 
                      (N133)? mem[809] : 
                      (N135)? mem[824] : 
                      (N137)? mem[839] : 
                      (N139)? mem[854] : 
                      (N141)? mem[869] : 
                      (N143)? mem[884] : 
                      (N145)? mem[899] : 
                      (N147)? mem[914] : 
                      (N149)? mem[929] : 
                      (N151)? mem[944] : 
                      (N153)? mem[959] : 1'b0;
  assign data_o[13] = (N90)? mem[13] : 
                      (N92)? mem[28] : 
                      (N94)? mem[43] : 
                      (N96)? mem[58] : 
                      (N98)? mem[73] : 
                      (N100)? mem[88] : 
                      (N102)? mem[103] : 
                      (N104)? mem[118] : 
                      (N106)? mem[133] : 
                      (N108)? mem[148] : 
                      (N110)? mem[163] : 
                      (N112)? mem[178] : 
                      (N114)? mem[193] : 
                      (N116)? mem[208] : 
                      (N118)? mem[223] : 
                      (N120)? mem[238] : 
                      (N122)? mem[253] : 
                      (N124)? mem[268] : 
                      (N126)? mem[283] : 
                      (N128)? mem[298] : 
                      (N130)? mem[313] : 
                      (N132)? mem[328] : 
                      (N134)? mem[343] : 
                      (N136)? mem[358] : 
                      (N138)? mem[373] : 
                      (N140)? mem[388] : 
                      (N142)? mem[403] : 
                      (N144)? mem[418] : 
                      (N146)? mem[433] : 
                      (N148)? mem[448] : 
                      (N150)? mem[463] : 
                      (N152)? mem[478] : 
                      (N91)? mem[493] : 
                      (N93)? mem[508] : 
                      (N95)? mem[523] : 
                      (N97)? mem[538] : 
                      (N99)? mem[553] : 
                      (N101)? mem[568] : 
                      (N103)? mem[583] : 
                      (N105)? mem[598] : 
                      (N107)? mem[613] : 
                      (N109)? mem[628] : 
                      (N111)? mem[643] : 
                      (N113)? mem[658] : 
                      (N115)? mem[673] : 
                      (N117)? mem[688] : 
                      (N119)? mem[703] : 
                      (N121)? mem[718] : 
                      (N123)? mem[733] : 
                      (N125)? mem[748] : 
                      (N127)? mem[763] : 
                      (N129)? mem[778] : 
                      (N131)? mem[793] : 
                      (N133)? mem[808] : 
                      (N135)? mem[823] : 
                      (N137)? mem[838] : 
                      (N139)? mem[853] : 
                      (N141)? mem[868] : 
                      (N143)? mem[883] : 
                      (N145)? mem[898] : 
                      (N147)? mem[913] : 
                      (N149)? mem[928] : 
                      (N151)? mem[943] : 
                      (N153)? mem[958] : 1'b0;
  assign data_o[12] = (N90)? mem[12] : 
                      (N92)? mem[27] : 
                      (N94)? mem[42] : 
                      (N96)? mem[57] : 
                      (N98)? mem[72] : 
                      (N100)? mem[87] : 
                      (N102)? mem[102] : 
                      (N104)? mem[117] : 
                      (N106)? mem[132] : 
                      (N108)? mem[147] : 
                      (N110)? mem[162] : 
                      (N112)? mem[177] : 
                      (N114)? mem[192] : 
                      (N116)? mem[207] : 
                      (N118)? mem[222] : 
                      (N120)? mem[237] : 
                      (N122)? mem[252] : 
                      (N124)? mem[267] : 
                      (N126)? mem[282] : 
                      (N128)? mem[297] : 
                      (N130)? mem[312] : 
                      (N132)? mem[327] : 
                      (N134)? mem[342] : 
                      (N136)? mem[357] : 
                      (N138)? mem[372] : 
                      (N140)? mem[387] : 
                      (N142)? mem[402] : 
                      (N144)? mem[417] : 
                      (N146)? mem[432] : 
                      (N148)? mem[447] : 
                      (N150)? mem[462] : 
                      (N152)? mem[477] : 
                      (N91)? mem[492] : 
                      (N93)? mem[507] : 
                      (N95)? mem[522] : 
                      (N97)? mem[537] : 
                      (N99)? mem[552] : 
                      (N101)? mem[567] : 
                      (N103)? mem[582] : 
                      (N105)? mem[597] : 
                      (N107)? mem[612] : 
                      (N109)? mem[627] : 
                      (N111)? mem[642] : 
                      (N113)? mem[657] : 
                      (N115)? mem[672] : 
                      (N117)? mem[687] : 
                      (N119)? mem[702] : 
                      (N121)? mem[717] : 
                      (N123)? mem[732] : 
                      (N125)? mem[747] : 
                      (N127)? mem[762] : 
                      (N129)? mem[777] : 
                      (N131)? mem[792] : 
                      (N133)? mem[807] : 
                      (N135)? mem[822] : 
                      (N137)? mem[837] : 
                      (N139)? mem[852] : 
                      (N141)? mem[867] : 
                      (N143)? mem[882] : 
                      (N145)? mem[897] : 
                      (N147)? mem[912] : 
                      (N149)? mem[927] : 
                      (N151)? mem[942] : 
                      (N153)? mem[957] : 1'b0;
  assign data_o[11] = (N90)? mem[11] : 
                      (N92)? mem[26] : 
                      (N94)? mem[41] : 
                      (N96)? mem[56] : 
                      (N98)? mem[71] : 
                      (N100)? mem[86] : 
                      (N102)? mem[101] : 
                      (N104)? mem[116] : 
                      (N106)? mem[131] : 
                      (N108)? mem[146] : 
                      (N110)? mem[161] : 
                      (N112)? mem[176] : 
                      (N114)? mem[191] : 
                      (N116)? mem[206] : 
                      (N118)? mem[221] : 
                      (N120)? mem[236] : 
                      (N122)? mem[251] : 
                      (N124)? mem[266] : 
                      (N126)? mem[281] : 
                      (N128)? mem[296] : 
                      (N130)? mem[311] : 
                      (N132)? mem[326] : 
                      (N134)? mem[341] : 
                      (N136)? mem[356] : 
                      (N138)? mem[371] : 
                      (N140)? mem[386] : 
                      (N142)? mem[401] : 
                      (N144)? mem[416] : 
                      (N146)? mem[431] : 
                      (N148)? mem[446] : 
                      (N150)? mem[461] : 
                      (N152)? mem[476] : 
                      (N91)? mem[491] : 
                      (N93)? mem[506] : 
                      (N95)? mem[521] : 
                      (N97)? mem[536] : 
                      (N99)? mem[551] : 
                      (N101)? mem[566] : 
                      (N103)? mem[581] : 
                      (N105)? mem[596] : 
                      (N107)? mem[611] : 
                      (N109)? mem[626] : 
                      (N111)? mem[641] : 
                      (N113)? mem[656] : 
                      (N115)? mem[671] : 
                      (N117)? mem[686] : 
                      (N119)? mem[701] : 
                      (N121)? mem[716] : 
                      (N123)? mem[731] : 
                      (N125)? mem[746] : 
                      (N127)? mem[761] : 
                      (N129)? mem[776] : 
                      (N131)? mem[791] : 
                      (N133)? mem[806] : 
                      (N135)? mem[821] : 
                      (N137)? mem[836] : 
                      (N139)? mem[851] : 
                      (N141)? mem[866] : 
                      (N143)? mem[881] : 
                      (N145)? mem[896] : 
                      (N147)? mem[911] : 
                      (N149)? mem[926] : 
                      (N151)? mem[941] : 
                      (N153)? mem[956] : 1'b0;
  assign data_o[10] = (N90)? mem[10] : 
                      (N92)? mem[25] : 
                      (N94)? mem[40] : 
                      (N96)? mem[55] : 
                      (N98)? mem[70] : 
                      (N100)? mem[85] : 
                      (N102)? mem[100] : 
                      (N104)? mem[115] : 
                      (N106)? mem[130] : 
                      (N108)? mem[145] : 
                      (N110)? mem[160] : 
                      (N112)? mem[175] : 
                      (N114)? mem[190] : 
                      (N116)? mem[205] : 
                      (N118)? mem[220] : 
                      (N120)? mem[235] : 
                      (N122)? mem[250] : 
                      (N124)? mem[265] : 
                      (N126)? mem[280] : 
                      (N128)? mem[295] : 
                      (N130)? mem[310] : 
                      (N132)? mem[325] : 
                      (N134)? mem[340] : 
                      (N136)? mem[355] : 
                      (N138)? mem[370] : 
                      (N140)? mem[385] : 
                      (N142)? mem[400] : 
                      (N144)? mem[415] : 
                      (N146)? mem[430] : 
                      (N148)? mem[445] : 
                      (N150)? mem[460] : 
                      (N152)? mem[475] : 
                      (N91)? mem[490] : 
                      (N93)? mem[505] : 
                      (N95)? mem[520] : 
                      (N97)? mem[535] : 
                      (N99)? mem[550] : 
                      (N101)? mem[565] : 
                      (N103)? mem[580] : 
                      (N105)? mem[595] : 
                      (N107)? mem[610] : 
                      (N109)? mem[625] : 
                      (N111)? mem[640] : 
                      (N113)? mem[655] : 
                      (N115)? mem[670] : 
                      (N117)? mem[685] : 
                      (N119)? mem[700] : 
                      (N121)? mem[715] : 
                      (N123)? mem[730] : 
                      (N125)? mem[745] : 
                      (N127)? mem[760] : 
                      (N129)? mem[775] : 
                      (N131)? mem[790] : 
                      (N133)? mem[805] : 
                      (N135)? mem[820] : 
                      (N137)? mem[835] : 
                      (N139)? mem[850] : 
                      (N141)? mem[865] : 
                      (N143)? mem[880] : 
                      (N145)? mem[895] : 
                      (N147)? mem[910] : 
                      (N149)? mem[925] : 
                      (N151)? mem[940] : 
                      (N153)? mem[955] : 1'b0;
  assign data_o[9] = (N90)? mem[9] : 
                     (N92)? mem[24] : 
                     (N94)? mem[39] : 
                     (N96)? mem[54] : 
                     (N98)? mem[69] : 
                     (N100)? mem[84] : 
                     (N102)? mem[99] : 
                     (N104)? mem[114] : 
                     (N106)? mem[129] : 
                     (N108)? mem[144] : 
                     (N110)? mem[159] : 
                     (N112)? mem[174] : 
                     (N114)? mem[189] : 
                     (N116)? mem[204] : 
                     (N118)? mem[219] : 
                     (N120)? mem[234] : 
                     (N122)? mem[249] : 
                     (N124)? mem[264] : 
                     (N126)? mem[279] : 
                     (N128)? mem[294] : 
                     (N130)? mem[309] : 
                     (N132)? mem[324] : 
                     (N134)? mem[339] : 
                     (N136)? mem[354] : 
                     (N138)? mem[369] : 
                     (N140)? mem[384] : 
                     (N142)? mem[399] : 
                     (N144)? mem[414] : 
                     (N146)? mem[429] : 
                     (N148)? mem[444] : 
                     (N150)? mem[459] : 
                     (N152)? mem[474] : 
                     (N91)? mem[489] : 
                     (N93)? mem[504] : 
                     (N95)? mem[519] : 
                     (N97)? mem[534] : 
                     (N99)? mem[549] : 
                     (N101)? mem[564] : 
                     (N103)? mem[579] : 
                     (N105)? mem[594] : 
                     (N107)? mem[609] : 
                     (N109)? mem[624] : 
                     (N111)? mem[639] : 
                     (N113)? mem[654] : 
                     (N115)? mem[669] : 
                     (N117)? mem[684] : 
                     (N119)? mem[699] : 
                     (N121)? mem[714] : 
                     (N123)? mem[729] : 
                     (N125)? mem[744] : 
                     (N127)? mem[759] : 
                     (N129)? mem[774] : 
                     (N131)? mem[789] : 
                     (N133)? mem[804] : 
                     (N135)? mem[819] : 
                     (N137)? mem[834] : 
                     (N139)? mem[849] : 
                     (N141)? mem[864] : 
                     (N143)? mem[879] : 
                     (N145)? mem[894] : 
                     (N147)? mem[909] : 
                     (N149)? mem[924] : 
                     (N151)? mem[939] : 
                     (N153)? mem[954] : 1'b0;
  assign data_o[8] = (N90)? mem[8] : 
                     (N92)? mem[23] : 
                     (N94)? mem[38] : 
                     (N96)? mem[53] : 
                     (N98)? mem[68] : 
                     (N100)? mem[83] : 
                     (N102)? mem[98] : 
                     (N104)? mem[113] : 
                     (N106)? mem[128] : 
                     (N108)? mem[143] : 
                     (N110)? mem[158] : 
                     (N112)? mem[173] : 
                     (N114)? mem[188] : 
                     (N116)? mem[203] : 
                     (N118)? mem[218] : 
                     (N120)? mem[233] : 
                     (N122)? mem[248] : 
                     (N124)? mem[263] : 
                     (N126)? mem[278] : 
                     (N128)? mem[293] : 
                     (N130)? mem[308] : 
                     (N132)? mem[323] : 
                     (N134)? mem[338] : 
                     (N136)? mem[353] : 
                     (N138)? mem[368] : 
                     (N140)? mem[383] : 
                     (N142)? mem[398] : 
                     (N144)? mem[413] : 
                     (N146)? mem[428] : 
                     (N148)? mem[443] : 
                     (N150)? mem[458] : 
                     (N152)? mem[473] : 
                     (N91)? mem[488] : 
                     (N93)? mem[503] : 
                     (N95)? mem[518] : 
                     (N97)? mem[533] : 
                     (N99)? mem[548] : 
                     (N101)? mem[563] : 
                     (N103)? mem[578] : 
                     (N105)? mem[593] : 
                     (N107)? mem[608] : 
                     (N109)? mem[623] : 
                     (N111)? mem[638] : 
                     (N113)? mem[653] : 
                     (N115)? mem[668] : 
                     (N117)? mem[683] : 
                     (N119)? mem[698] : 
                     (N121)? mem[713] : 
                     (N123)? mem[728] : 
                     (N125)? mem[743] : 
                     (N127)? mem[758] : 
                     (N129)? mem[773] : 
                     (N131)? mem[788] : 
                     (N133)? mem[803] : 
                     (N135)? mem[818] : 
                     (N137)? mem[833] : 
                     (N139)? mem[848] : 
                     (N141)? mem[863] : 
                     (N143)? mem[878] : 
                     (N145)? mem[893] : 
                     (N147)? mem[908] : 
                     (N149)? mem[923] : 
                     (N151)? mem[938] : 
                     (N153)? mem[953] : 1'b0;
  assign data_o[7] = (N90)? mem[7] : 
                     (N92)? mem[22] : 
                     (N94)? mem[37] : 
                     (N96)? mem[52] : 
                     (N98)? mem[67] : 
                     (N100)? mem[82] : 
                     (N102)? mem[97] : 
                     (N104)? mem[112] : 
                     (N106)? mem[127] : 
                     (N108)? mem[142] : 
                     (N110)? mem[157] : 
                     (N112)? mem[172] : 
                     (N114)? mem[187] : 
                     (N116)? mem[202] : 
                     (N118)? mem[217] : 
                     (N120)? mem[232] : 
                     (N122)? mem[247] : 
                     (N124)? mem[262] : 
                     (N126)? mem[277] : 
                     (N128)? mem[292] : 
                     (N130)? mem[307] : 
                     (N132)? mem[322] : 
                     (N134)? mem[337] : 
                     (N136)? mem[352] : 
                     (N138)? mem[367] : 
                     (N140)? mem[382] : 
                     (N142)? mem[397] : 
                     (N144)? mem[412] : 
                     (N146)? mem[427] : 
                     (N148)? mem[442] : 
                     (N150)? mem[457] : 
                     (N152)? mem[472] : 
                     (N91)? mem[487] : 
                     (N93)? mem[502] : 
                     (N95)? mem[517] : 
                     (N97)? mem[532] : 
                     (N99)? mem[547] : 
                     (N101)? mem[562] : 
                     (N103)? mem[577] : 
                     (N105)? mem[592] : 
                     (N107)? mem[607] : 
                     (N109)? mem[622] : 
                     (N111)? mem[637] : 
                     (N113)? mem[652] : 
                     (N115)? mem[667] : 
                     (N117)? mem[682] : 
                     (N119)? mem[697] : 
                     (N121)? mem[712] : 
                     (N123)? mem[727] : 
                     (N125)? mem[742] : 
                     (N127)? mem[757] : 
                     (N129)? mem[772] : 
                     (N131)? mem[787] : 
                     (N133)? mem[802] : 
                     (N135)? mem[817] : 
                     (N137)? mem[832] : 
                     (N139)? mem[847] : 
                     (N141)? mem[862] : 
                     (N143)? mem[877] : 
                     (N145)? mem[892] : 
                     (N147)? mem[907] : 
                     (N149)? mem[922] : 
                     (N151)? mem[937] : 
                     (N153)? mem[952] : 1'b0;
  assign data_o[6] = (N90)? mem[6] : 
                     (N92)? mem[21] : 
                     (N94)? mem[36] : 
                     (N96)? mem[51] : 
                     (N98)? mem[66] : 
                     (N100)? mem[81] : 
                     (N102)? mem[96] : 
                     (N104)? mem[111] : 
                     (N106)? mem[126] : 
                     (N108)? mem[141] : 
                     (N110)? mem[156] : 
                     (N112)? mem[171] : 
                     (N114)? mem[186] : 
                     (N116)? mem[201] : 
                     (N118)? mem[216] : 
                     (N120)? mem[231] : 
                     (N122)? mem[246] : 
                     (N124)? mem[261] : 
                     (N126)? mem[276] : 
                     (N128)? mem[291] : 
                     (N130)? mem[306] : 
                     (N132)? mem[321] : 
                     (N134)? mem[336] : 
                     (N136)? mem[351] : 
                     (N138)? mem[366] : 
                     (N140)? mem[381] : 
                     (N142)? mem[396] : 
                     (N144)? mem[411] : 
                     (N146)? mem[426] : 
                     (N148)? mem[441] : 
                     (N150)? mem[456] : 
                     (N152)? mem[471] : 
                     (N91)? mem[486] : 
                     (N93)? mem[501] : 
                     (N95)? mem[516] : 
                     (N97)? mem[531] : 
                     (N99)? mem[546] : 
                     (N101)? mem[561] : 
                     (N103)? mem[576] : 
                     (N105)? mem[591] : 
                     (N107)? mem[606] : 
                     (N109)? mem[621] : 
                     (N111)? mem[636] : 
                     (N113)? mem[651] : 
                     (N115)? mem[666] : 
                     (N117)? mem[681] : 
                     (N119)? mem[696] : 
                     (N121)? mem[711] : 
                     (N123)? mem[726] : 
                     (N125)? mem[741] : 
                     (N127)? mem[756] : 
                     (N129)? mem[771] : 
                     (N131)? mem[786] : 
                     (N133)? mem[801] : 
                     (N135)? mem[816] : 
                     (N137)? mem[831] : 
                     (N139)? mem[846] : 
                     (N141)? mem[861] : 
                     (N143)? mem[876] : 
                     (N145)? mem[891] : 
                     (N147)? mem[906] : 
                     (N149)? mem[921] : 
                     (N151)? mem[936] : 
                     (N153)? mem[951] : 1'b0;
  assign data_o[5] = (N90)? mem[5] : 
                     (N92)? mem[20] : 
                     (N94)? mem[35] : 
                     (N96)? mem[50] : 
                     (N98)? mem[65] : 
                     (N100)? mem[80] : 
                     (N102)? mem[95] : 
                     (N104)? mem[110] : 
                     (N106)? mem[125] : 
                     (N108)? mem[140] : 
                     (N110)? mem[155] : 
                     (N112)? mem[170] : 
                     (N114)? mem[185] : 
                     (N116)? mem[200] : 
                     (N118)? mem[215] : 
                     (N120)? mem[230] : 
                     (N122)? mem[245] : 
                     (N124)? mem[260] : 
                     (N126)? mem[275] : 
                     (N128)? mem[290] : 
                     (N130)? mem[305] : 
                     (N132)? mem[320] : 
                     (N134)? mem[335] : 
                     (N136)? mem[350] : 
                     (N138)? mem[365] : 
                     (N140)? mem[380] : 
                     (N142)? mem[395] : 
                     (N144)? mem[410] : 
                     (N146)? mem[425] : 
                     (N148)? mem[440] : 
                     (N150)? mem[455] : 
                     (N152)? mem[470] : 
                     (N91)? mem[485] : 
                     (N93)? mem[500] : 
                     (N95)? mem[515] : 
                     (N97)? mem[530] : 
                     (N99)? mem[545] : 
                     (N101)? mem[560] : 
                     (N103)? mem[575] : 
                     (N105)? mem[590] : 
                     (N107)? mem[605] : 
                     (N109)? mem[620] : 
                     (N111)? mem[635] : 
                     (N113)? mem[650] : 
                     (N115)? mem[665] : 
                     (N117)? mem[680] : 
                     (N119)? mem[695] : 
                     (N121)? mem[710] : 
                     (N123)? mem[725] : 
                     (N125)? mem[740] : 
                     (N127)? mem[755] : 
                     (N129)? mem[770] : 
                     (N131)? mem[785] : 
                     (N133)? mem[800] : 
                     (N135)? mem[815] : 
                     (N137)? mem[830] : 
                     (N139)? mem[845] : 
                     (N141)? mem[860] : 
                     (N143)? mem[875] : 
                     (N145)? mem[890] : 
                     (N147)? mem[905] : 
                     (N149)? mem[920] : 
                     (N151)? mem[935] : 
                     (N153)? mem[950] : 1'b0;
  assign data_o[4] = (N90)? mem[4] : 
                     (N92)? mem[19] : 
                     (N94)? mem[34] : 
                     (N96)? mem[49] : 
                     (N98)? mem[64] : 
                     (N100)? mem[79] : 
                     (N102)? mem[94] : 
                     (N104)? mem[109] : 
                     (N106)? mem[124] : 
                     (N108)? mem[139] : 
                     (N110)? mem[154] : 
                     (N112)? mem[169] : 
                     (N114)? mem[184] : 
                     (N116)? mem[199] : 
                     (N118)? mem[214] : 
                     (N120)? mem[229] : 
                     (N122)? mem[244] : 
                     (N124)? mem[259] : 
                     (N126)? mem[274] : 
                     (N128)? mem[289] : 
                     (N130)? mem[304] : 
                     (N132)? mem[319] : 
                     (N134)? mem[334] : 
                     (N136)? mem[349] : 
                     (N138)? mem[364] : 
                     (N140)? mem[379] : 
                     (N142)? mem[394] : 
                     (N144)? mem[409] : 
                     (N146)? mem[424] : 
                     (N148)? mem[439] : 
                     (N150)? mem[454] : 
                     (N152)? mem[469] : 
                     (N91)? mem[484] : 
                     (N93)? mem[499] : 
                     (N95)? mem[514] : 
                     (N97)? mem[529] : 
                     (N99)? mem[544] : 
                     (N101)? mem[559] : 
                     (N103)? mem[574] : 
                     (N105)? mem[589] : 
                     (N107)? mem[604] : 
                     (N109)? mem[619] : 
                     (N111)? mem[634] : 
                     (N113)? mem[649] : 
                     (N115)? mem[664] : 
                     (N117)? mem[679] : 
                     (N119)? mem[694] : 
                     (N121)? mem[709] : 
                     (N123)? mem[724] : 
                     (N125)? mem[739] : 
                     (N127)? mem[754] : 
                     (N129)? mem[769] : 
                     (N131)? mem[784] : 
                     (N133)? mem[799] : 
                     (N135)? mem[814] : 
                     (N137)? mem[829] : 
                     (N139)? mem[844] : 
                     (N141)? mem[859] : 
                     (N143)? mem[874] : 
                     (N145)? mem[889] : 
                     (N147)? mem[904] : 
                     (N149)? mem[919] : 
                     (N151)? mem[934] : 
                     (N153)? mem[949] : 1'b0;
  assign data_o[3] = (N90)? mem[3] : 
                     (N92)? mem[18] : 
                     (N94)? mem[33] : 
                     (N96)? mem[48] : 
                     (N98)? mem[63] : 
                     (N100)? mem[78] : 
                     (N102)? mem[93] : 
                     (N104)? mem[108] : 
                     (N106)? mem[123] : 
                     (N108)? mem[138] : 
                     (N110)? mem[153] : 
                     (N112)? mem[168] : 
                     (N114)? mem[183] : 
                     (N116)? mem[198] : 
                     (N118)? mem[213] : 
                     (N120)? mem[228] : 
                     (N122)? mem[243] : 
                     (N124)? mem[258] : 
                     (N126)? mem[273] : 
                     (N128)? mem[288] : 
                     (N130)? mem[303] : 
                     (N132)? mem[318] : 
                     (N134)? mem[333] : 
                     (N136)? mem[348] : 
                     (N138)? mem[363] : 
                     (N140)? mem[378] : 
                     (N142)? mem[393] : 
                     (N144)? mem[408] : 
                     (N146)? mem[423] : 
                     (N148)? mem[438] : 
                     (N150)? mem[453] : 
                     (N152)? mem[468] : 
                     (N91)? mem[483] : 
                     (N93)? mem[498] : 
                     (N95)? mem[513] : 
                     (N97)? mem[528] : 
                     (N99)? mem[543] : 
                     (N101)? mem[558] : 
                     (N103)? mem[573] : 
                     (N105)? mem[588] : 
                     (N107)? mem[603] : 
                     (N109)? mem[618] : 
                     (N111)? mem[633] : 
                     (N113)? mem[648] : 
                     (N115)? mem[663] : 
                     (N117)? mem[678] : 
                     (N119)? mem[693] : 
                     (N121)? mem[708] : 
                     (N123)? mem[723] : 
                     (N125)? mem[738] : 
                     (N127)? mem[753] : 
                     (N129)? mem[768] : 
                     (N131)? mem[783] : 
                     (N133)? mem[798] : 
                     (N135)? mem[813] : 
                     (N137)? mem[828] : 
                     (N139)? mem[843] : 
                     (N141)? mem[858] : 
                     (N143)? mem[873] : 
                     (N145)? mem[888] : 
                     (N147)? mem[903] : 
                     (N149)? mem[918] : 
                     (N151)? mem[933] : 
                     (N153)? mem[948] : 1'b0;
  assign data_o[2] = (N90)? mem[2] : 
                     (N92)? mem[17] : 
                     (N94)? mem[32] : 
                     (N96)? mem[47] : 
                     (N98)? mem[62] : 
                     (N100)? mem[77] : 
                     (N102)? mem[92] : 
                     (N104)? mem[107] : 
                     (N106)? mem[122] : 
                     (N108)? mem[137] : 
                     (N110)? mem[152] : 
                     (N112)? mem[167] : 
                     (N114)? mem[182] : 
                     (N116)? mem[197] : 
                     (N118)? mem[212] : 
                     (N120)? mem[227] : 
                     (N122)? mem[242] : 
                     (N124)? mem[257] : 
                     (N126)? mem[272] : 
                     (N128)? mem[287] : 
                     (N130)? mem[302] : 
                     (N132)? mem[317] : 
                     (N134)? mem[332] : 
                     (N136)? mem[347] : 
                     (N138)? mem[362] : 
                     (N140)? mem[377] : 
                     (N142)? mem[392] : 
                     (N144)? mem[407] : 
                     (N146)? mem[422] : 
                     (N148)? mem[437] : 
                     (N150)? mem[452] : 
                     (N152)? mem[467] : 
                     (N91)? mem[482] : 
                     (N93)? mem[497] : 
                     (N95)? mem[512] : 
                     (N97)? mem[527] : 
                     (N99)? mem[542] : 
                     (N101)? mem[557] : 
                     (N103)? mem[572] : 
                     (N105)? mem[587] : 
                     (N107)? mem[602] : 
                     (N109)? mem[617] : 
                     (N111)? mem[632] : 
                     (N113)? mem[647] : 
                     (N115)? mem[662] : 
                     (N117)? mem[677] : 
                     (N119)? mem[692] : 
                     (N121)? mem[707] : 
                     (N123)? mem[722] : 
                     (N125)? mem[737] : 
                     (N127)? mem[752] : 
                     (N129)? mem[767] : 
                     (N131)? mem[782] : 
                     (N133)? mem[797] : 
                     (N135)? mem[812] : 
                     (N137)? mem[827] : 
                     (N139)? mem[842] : 
                     (N141)? mem[857] : 
                     (N143)? mem[872] : 
                     (N145)? mem[887] : 
                     (N147)? mem[902] : 
                     (N149)? mem[917] : 
                     (N151)? mem[932] : 
                     (N153)? mem[947] : 1'b0;
  assign data_o[1] = (N90)? mem[1] : 
                     (N92)? mem[16] : 
                     (N94)? mem[31] : 
                     (N96)? mem[46] : 
                     (N98)? mem[61] : 
                     (N100)? mem[76] : 
                     (N102)? mem[91] : 
                     (N104)? mem[106] : 
                     (N106)? mem[121] : 
                     (N108)? mem[136] : 
                     (N110)? mem[151] : 
                     (N112)? mem[166] : 
                     (N114)? mem[181] : 
                     (N116)? mem[196] : 
                     (N118)? mem[211] : 
                     (N120)? mem[226] : 
                     (N122)? mem[241] : 
                     (N124)? mem[256] : 
                     (N126)? mem[271] : 
                     (N128)? mem[286] : 
                     (N130)? mem[301] : 
                     (N132)? mem[316] : 
                     (N134)? mem[331] : 
                     (N136)? mem[346] : 
                     (N138)? mem[361] : 
                     (N140)? mem[376] : 
                     (N142)? mem[391] : 
                     (N144)? mem[406] : 
                     (N146)? mem[421] : 
                     (N148)? mem[436] : 
                     (N150)? mem[451] : 
                     (N152)? mem[466] : 
                     (N91)? mem[481] : 
                     (N93)? mem[496] : 
                     (N95)? mem[511] : 
                     (N97)? mem[526] : 
                     (N99)? mem[541] : 
                     (N101)? mem[556] : 
                     (N103)? mem[571] : 
                     (N105)? mem[586] : 
                     (N107)? mem[601] : 
                     (N109)? mem[616] : 
                     (N111)? mem[631] : 
                     (N113)? mem[646] : 
                     (N115)? mem[661] : 
                     (N117)? mem[676] : 
                     (N119)? mem[691] : 
                     (N121)? mem[706] : 
                     (N123)? mem[721] : 
                     (N125)? mem[736] : 
                     (N127)? mem[751] : 
                     (N129)? mem[766] : 
                     (N131)? mem[781] : 
                     (N133)? mem[796] : 
                     (N135)? mem[811] : 
                     (N137)? mem[826] : 
                     (N139)? mem[841] : 
                     (N141)? mem[856] : 
                     (N143)? mem[871] : 
                     (N145)? mem[886] : 
                     (N147)? mem[901] : 
                     (N149)? mem[916] : 
                     (N151)? mem[931] : 
                     (N153)? mem[946] : 1'b0;
  assign data_o[0] = (N90)? mem[0] : 
                     (N92)? mem[15] : 
                     (N94)? mem[30] : 
                     (N96)? mem[45] : 
                     (N98)? mem[60] : 
                     (N100)? mem[75] : 
                     (N102)? mem[90] : 
                     (N104)? mem[105] : 
                     (N106)? mem[120] : 
                     (N108)? mem[135] : 
                     (N110)? mem[150] : 
                     (N112)? mem[165] : 
                     (N114)? mem[180] : 
                     (N116)? mem[195] : 
                     (N118)? mem[210] : 
                     (N120)? mem[225] : 
                     (N122)? mem[240] : 
                     (N124)? mem[255] : 
                     (N126)? mem[270] : 
                     (N128)? mem[285] : 
                     (N130)? mem[300] : 
                     (N132)? mem[315] : 
                     (N134)? mem[330] : 
                     (N136)? mem[345] : 
                     (N138)? mem[360] : 
                     (N140)? mem[375] : 
                     (N142)? mem[390] : 
                     (N144)? mem[405] : 
                     (N146)? mem[420] : 
                     (N148)? mem[435] : 
                     (N150)? mem[450] : 
                     (N152)? mem[465] : 
                     (N91)? mem[480] : 
                     (N93)? mem[495] : 
                     (N95)? mem[510] : 
                     (N97)? mem[525] : 
                     (N99)? mem[540] : 
                     (N101)? mem[555] : 
                     (N103)? mem[570] : 
                     (N105)? mem[585] : 
                     (N107)? mem[600] : 
                     (N109)? mem[615] : 
                     (N111)? mem[630] : 
                     (N113)? mem[645] : 
                     (N115)? mem[660] : 
                     (N117)? mem[675] : 
                     (N119)? mem[690] : 
                     (N121)? mem[705] : 
                     (N123)? mem[720] : 
                     (N125)? mem[735] : 
                     (N127)? mem[750] : 
                     (N129)? mem[765] : 
                     (N131)? mem[780] : 
                     (N133)? mem[795] : 
                     (N135)? mem[810] : 
                     (N137)? mem[825] : 
                     (N139)? mem[840] : 
                     (N141)? mem[855] : 
                     (N143)? mem[870] : 
                     (N145)? mem[885] : 
                     (N147)? mem[900] : 
                     (N149)? mem[915] : 
                     (N151)? mem[930] : 
                     (N153)? mem[945] : 1'b0;

  always @(posedge clk_i) begin
    if(N2248) begin
      mem_959_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2247) begin
      mem_958_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2246) begin
      mem_957_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2245) begin
      mem_956_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2244) begin
      mem_955_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2243) begin
      mem_954_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2242) begin
      mem_953_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2241) begin
      mem_952_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2240) begin
      mem_951_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2239) begin
      mem_950_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2238) begin
      mem_949_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2237) begin
      mem_948_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2236) begin
      mem_947_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2235) begin
      mem_946_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2234) begin
      mem_945_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2233) begin
      mem_944_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2232) begin
      mem_943_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2231) begin
      mem_942_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2230) begin
      mem_941_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2229) begin
      mem_940_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2228) begin
      mem_939_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2227) begin
      mem_938_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2226) begin
      mem_937_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2225) begin
      mem_936_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2224) begin
      mem_935_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2223) begin
      mem_934_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2222) begin
      mem_933_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2221) begin
      mem_932_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2220) begin
      mem_931_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2219) begin
      mem_930_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2218) begin
      mem_929_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2217) begin
      mem_928_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2216) begin
      mem_927_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2215) begin
      mem_926_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2214) begin
      mem_925_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2213) begin
      mem_924_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2212) begin
      mem_923_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2211) begin
      mem_922_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2210) begin
      mem_921_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2209) begin
      mem_920_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2208) begin
      mem_919_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2207) begin
      mem_918_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2206) begin
      mem_917_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2205) begin
      mem_916_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2204) begin
      mem_915_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2203) begin
      mem_914_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2202) begin
      mem_913_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2201) begin
      mem_912_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2200) begin
      mem_911_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2199) begin
      mem_910_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2198) begin
      mem_909_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2197) begin
      mem_908_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2196) begin
      mem_907_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2195) begin
      mem_906_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2194) begin
      mem_905_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2193) begin
      mem_904_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2192) begin
      mem_903_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2191) begin
      mem_902_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2190) begin
      mem_901_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2189) begin
      mem_900_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2188) begin
      mem_899_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2187) begin
      mem_898_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2186) begin
      mem_897_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2185) begin
      mem_896_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2184) begin
      mem_895_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2183) begin
      mem_894_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2182) begin
      mem_893_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2181) begin
      mem_892_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2180) begin
      mem_891_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2179) begin
      mem_890_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2178) begin
      mem_889_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2177) begin
      mem_888_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2176) begin
      mem_887_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2175) begin
      mem_886_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2174) begin
      mem_885_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2173) begin
      mem_884_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2172) begin
      mem_883_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2171) begin
      mem_882_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2170) begin
      mem_881_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2169) begin
      mem_880_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2168) begin
      mem_879_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2167) begin
      mem_878_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2166) begin
      mem_877_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2165) begin
      mem_876_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2164) begin
      mem_875_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2163) begin
      mem_874_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2162) begin
      mem_873_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2161) begin
      mem_872_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2160) begin
      mem_871_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2159) begin
      mem_870_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2158) begin
      mem_869_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2157) begin
      mem_868_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2156) begin
      mem_867_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2155) begin
      mem_866_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2154) begin
      mem_865_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2153) begin
      mem_864_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2152) begin
      mem_863_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2151) begin
      mem_862_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2150) begin
      mem_861_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2149) begin
      mem_860_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2148) begin
      mem_859_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2147) begin
      mem_858_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2146) begin
      mem_857_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2145) begin
      mem_856_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2144) begin
      mem_855_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2143) begin
      mem_854_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2142) begin
      mem_853_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2141) begin
      mem_852_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2140) begin
      mem_851_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2139) begin
      mem_850_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2138) begin
      mem_849_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2137) begin
      mem_848_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2136) begin
      mem_847_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2135) begin
      mem_846_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2134) begin
      mem_845_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2133) begin
      mem_844_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2132) begin
      mem_843_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2131) begin
      mem_842_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2130) begin
      mem_841_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2129) begin
      mem_840_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2128) begin
      mem_839_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2127) begin
      mem_838_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2126) begin
      mem_837_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2125) begin
      mem_836_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2124) begin
      mem_835_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2123) begin
      mem_834_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2122) begin
      mem_833_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2121) begin
      mem_832_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2120) begin
      mem_831_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2119) begin
      mem_830_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2118) begin
      mem_829_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2117) begin
      mem_828_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2116) begin
      mem_827_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2115) begin
      mem_826_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2114) begin
      mem_825_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2113) begin
      mem_824_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2112) begin
      mem_823_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2111) begin
      mem_822_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2110) begin
      mem_821_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2109) begin
      mem_820_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2108) begin
      mem_819_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2107) begin
      mem_818_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2106) begin
      mem_817_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2105) begin
      mem_816_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2104) begin
      mem_815_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2103) begin
      mem_814_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2102) begin
      mem_813_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2101) begin
      mem_812_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2100) begin
      mem_811_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2099) begin
      mem_810_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2098) begin
      mem_809_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2097) begin
      mem_808_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2096) begin
      mem_807_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2095) begin
      mem_806_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2094) begin
      mem_805_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2093) begin
      mem_804_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2092) begin
      mem_803_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2091) begin
      mem_802_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2090) begin
      mem_801_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2089) begin
      mem_800_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2088) begin
      mem_799_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2087) begin
      mem_798_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2086) begin
      mem_797_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2085) begin
      mem_796_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2084) begin
      mem_795_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2083) begin
      mem_794_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2082) begin
      mem_793_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2081) begin
      mem_792_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2080) begin
      mem_791_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2079) begin
      mem_790_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2078) begin
      mem_789_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2077) begin
      mem_788_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2076) begin
      mem_787_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2075) begin
      mem_786_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2074) begin
      mem_785_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2073) begin
      mem_784_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2072) begin
      mem_783_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2071) begin
      mem_782_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2070) begin
      mem_781_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2069) begin
      mem_780_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2068) begin
      mem_779_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2067) begin
      mem_778_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2066) begin
      mem_777_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2065) begin
      mem_776_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2064) begin
      mem_775_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2063) begin
      mem_774_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2062) begin
      mem_773_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2061) begin
      mem_772_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2060) begin
      mem_771_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2059) begin
      mem_770_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2058) begin
      mem_769_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2057) begin
      mem_768_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2056) begin
      mem_767_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2055) begin
      mem_766_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      mem_765_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2053) begin
      mem_764_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2052) begin
      mem_763_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2051) begin
      mem_762_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2050) begin
      mem_761_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2049) begin
      mem_760_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2048) begin
      mem_759_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2047) begin
      mem_758_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2046) begin
      mem_757_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2045) begin
      mem_756_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2044) begin
      mem_755_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2043) begin
      mem_754_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2042) begin
      mem_753_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2041) begin
      mem_752_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2040) begin
      mem_751_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2039) begin
      mem_750_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2038) begin
      mem_749_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2037) begin
      mem_748_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2036) begin
      mem_747_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2035) begin
      mem_746_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2034) begin
      mem_745_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2033) begin
      mem_744_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2032) begin
      mem_743_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2031) begin
      mem_742_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2030) begin
      mem_741_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2029) begin
      mem_740_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2028) begin
      mem_739_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2027) begin
      mem_738_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2026) begin
      mem_737_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2025) begin
      mem_736_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2024) begin
      mem_735_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2023) begin
      mem_734_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2022) begin
      mem_733_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2021) begin
      mem_732_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2020) begin
      mem_731_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2019) begin
      mem_730_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2018) begin
      mem_729_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2017) begin
      mem_728_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2016) begin
      mem_727_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2015) begin
      mem_726_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2014) begin
      mem_725_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2013) begin
      mem_724_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2012) begin
      mem_723_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2011) begin
      mem_722_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2010) begin
      mem_721_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2009) begin
      mem_720_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2008) begin
      mem_719_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2007) begin
      mem_718_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2006) begin
      mem_717_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      mem_716_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2004) begin
      mem_715_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2003) begin
      mem_714_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2002) begin
      mem_713_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2001) begin
      mem_712_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2000) begin
      mem_711_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1999) begin
      mem_710_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1998) begin
      mem_709_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1997) begin
      mem_708_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1996) begin
      mem_707_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1995) begin
      mem_706_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1994) begin
      mem_705_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1993) begin
      mem_704_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1992) begin
      mem_703_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1991) begin
      mem_702_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1990) begin
      mem_701_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1989) begin
      mem_700_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1988) begin
      mem_699_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1987) begin
      mem_698_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1986) begin
      mem_697_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1985) begin
      mem_696_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1984) begin
      mem_695_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1983) begin
      mem_694_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1982) begin
      mem_693_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1981) begin
      mem_692_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1980) begin
      mem_691_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1979) begin
      mem_690_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1978) begin
      mem_689_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1977) begin
      mem_688_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1976) begin
      mem_687_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1975) begin
      mem_686_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1974) begin
      mem_685_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1973) begin
      mem_684_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1972) begin
      mem_683_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1971) begin
      mem_682_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1970) begin
      mem_681_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1969) begin
      mem_680_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1968) begin
      mem_679_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1967) begin
      mem_678_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1966) begin
      mem_677_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1965) begin
      mem_676_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1964) begin
      mem_675_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1963) begin
      mem_674_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1962) begin
      mem_673_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1961) begin
      mem_672_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1960) begin
      mem_671_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1959) begin
      mem_670_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1958) begin
      mem_669_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1957) begin
      mem_668_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      mem_667_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1955) begin
      mem_666_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1954) begin
      mem_665_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1953) begin
      mem_664_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1952) begin
      mem_663_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1951) begin
      mem_662_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1950) begin
      mem_661_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1949) begin
      mem_660_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1948) begin
      mem_659_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1947) begin
      mem_658_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1946) begin
      mem_657_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1945) begin
      mem_656_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1944) begin
      mem_655_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1943) begin
      mem_654_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1942) begin
      mem_653_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1941) begin
      mem_652_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1940) begin
      mem_651_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1939) begin
      mem_650_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1938) begin
      mem_649_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1937) begin
      mem_648_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1936) begin
      mem_647_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1935) begin
      mem_646_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1934) begin
      mem_645_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1933) begin
      mem_644_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1932) begin
      mem_643_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1931) begin
      mem_642_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1930) begin
      mem_641_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1929) begin
      mem_640_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1928) begin
      mem_639_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1927) begin
      mem_638_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1926) begin
      mem_637_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1925) begin
      mem_636_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1924) begin
      mem_635_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1923) begin
      mem_634_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1922) begin
      mem_633_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1921) begin
      mem_632_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1920) begin
      mem_631_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1919) begin
      mem_630_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1918) begin
      mem_629_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1917) begin
      mem_628_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1916) begin
      mem_627_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1915) begin
      mem_626_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1914) begin
      mem_625_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1913) begin
      mem_624_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1912) begin
      mem_623_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1911) begin
      mem_622_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1910) begin
      mem_621_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1909) begin
      mem_620_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1908) begin
      mem_619_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      mem_618_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1906) begin
      mem_617_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1905) begin
      mem_616_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1904) begin
      mem_615_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1903) begin
      mem_614_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1902) begin
      mem_613_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1901) begin
      mem_612_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1900) begin
      mem_611_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1899) begin
      mem_610_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1898) begin
      mem_609_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1897) begin
      mem_608_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1896) begin
      mem_607_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1895) begin
      mem_606_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1894) begin
      mem_605_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1893) begin
      mem_604_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1892) begin
      mem_603_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1891) begin
      mem_602_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1890) begin
      mem_601_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1889) begin
      mem_600_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1888) begin
      mem_599_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1887) begin
      mem_598_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1886) begin
      mem_597_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1885) begin
      mem_596_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1884) begin
      mem_595_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1883) begin
      mem_594_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1882) begin
      mem_593_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1881) begin
      mem_592_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1880) begin
      mem_591_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1879) begin
      mem_590_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1878) begin
      mem_589_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1877) begin
      mem_588_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1876) begin
      mem_587_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1875) begin
      mem_586_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1874) begin
      mem_585_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1873) begin
      mem_584_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1872) begin
      mem_583_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1871) begin
      mem_582_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1870) begin
      mem_581_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1869) begin
      mem_580_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1868) begin
      mem_579_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1867) begin
      mem_578_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1866) begin
      mem_577_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1865) begin
      mem_576_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1864) begin
      mem_575_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1863) begin
      mem_574_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1862) begin
      mem_573_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1861) begin
      mem_572_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1860) begin
      mem_571_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1859) begin
      mem_570_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      mem_569_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1857) begin
      mem_568_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1856) begin
      mem_567_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1855) begin
      mem_566_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1854) begin
      mem_565_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1853) begin
      mem_564_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1852) begin
      mem_563_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1851) begin
      mem_562_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1850) begin
      mem_561_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1849) begin
      mem_560_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1848) begin
      mem_559_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1847) begin
      mem_558_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1846) begin
      mem_557_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1845) begin
      mem_556_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1844) begin
      mem_555_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1843) begin
      mem_554_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1842) begin
      mem_553_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1841) begin
      mem_552_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1840) begin
      mem_551_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1839) begin
      mem_550_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1838) begin
      mem_549_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1837) begin
      mem_548_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1836) begin
      mem_547_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1835) begin
      mem_546_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1834) begin
      mem_545_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1833) begin
      mem_544_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1832) begin
      mem_543_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1831) begin
      mem_542_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1830) begin
      mem_541_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1829) begin
      mem_540_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1828) begin
      mem_539_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1827) begin
      mem_538_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1826) begin
      mem_537_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1825) begin
      mem_536_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1824) begin
      mem_535_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1823) begin
      mem_534_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1822) begin
      mem_533_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1821) begin
      mem_532_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1820) begin
      mem_531_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1819) begin
      mem_530_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1818) begin
      mem_529_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1817) begin
      mem_528_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1816) begin
      mem_527_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1815) begin
      mem_526_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1814) begin
      mem_525_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1813) begin
      mem_524_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1812) begin
      mem_523_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1811) begin
      mem_522_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1810) begin
      mem_521_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      mem_520_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1808) begin
      mem_519_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1807) begin
      mem_518_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1806) begin
      mem_517_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1805) begin
      mem_516_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1804) begin
      mem_515_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1803) begin
      mem_514_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1802) begin
      mem_513_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1801) begin
      mem_512_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1800) begin
      mem_511_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1799) begin
      mem_510_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1798) begin
      mem_509_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1797) begin
      mem_508_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1796) begin
      mem_507_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1795) begin
      mem_506_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1794) begin
      mem_505_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1793) begin
      mem_504_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1792) begin
      mem_503_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1791) begin
      mem_502_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1790) begin
      mem_501_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1789) begin
      mem_500_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1788) begin
      mem_499_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1787) begin
      mem_498_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1786) begin
      mem_497_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1785) begin
      mem_496_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1784) begin
      mem_495_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1783) begin
      mem_494_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1782) begin
      mem_493_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1781) begin
      mem_492_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1780) begin
      mem_491_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1779) begin
      mem_490_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1778) begin
      mem_489_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1777) begin
      mem_488_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1776) begin
      mem_487_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1775) begin
      mem_486_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1774) begin
      mem_485_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1773) begin
      mem_484_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1772) begin
      mem_483_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1771) begin
      mem_482_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1770) begin
      mem_481_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1769) begin
      mem_480_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1768) begin
      mem_479_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1767) begin
      mem_478_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1766) begin
      mem_477_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1765) begin
      mem_476_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1764) begin
      mem_475_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1763) begin
      mem_474_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1762) begin
      mem_473_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1761) begin
      mem_472_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      mem_471_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1759) begin
      mem_470_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1758) begin
      mem_469_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1757) begin
      mem_468_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1756) begin
      mem_467_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1755) begin
      mem_466_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1754) begin
      mem_465_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1753) begin
      mem_464_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1752) begin
      mem_463_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1751) begin
      mem_462_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1750) begin
      mem_461_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1749) begin
      mem_460_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1748) begin
      mem_459_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1747) begin
      mem_458_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1746) begin
      mem_457_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1745) begin
      mem_456_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1744) begin
      mem_455_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1743) begin
      mem_454_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1742) begin
      mem_453_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1741) begin
      mem_452_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1740) begin
      mem_451_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1739) begin
      mem_450_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1738) begin
      mem_449_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1737) begin
      mem_448_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1736) begin
      mem_447_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1735) begin
      mem_446_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1734) begin
      mem_445_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1733) begin
      mem_444_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1732) begin
      mem_443_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1731) begin
      mem_442_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1730) begin
      mem_441_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1729) begin
      mem_440_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1728) begin
      mem_439_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1727) begin
      mem_438_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1726) begin
      mem_437_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1725) begin
      mem_436_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1724) begin
      mem_435_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1723) begin
      mem_434_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1722) begin
      mem_433_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1721) begin
      mem_432_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1720) begin
      mem_431_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1719) begin
      mem_430_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1718) begin
      mem_429_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      mem_428_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1716) begin
      mem_427_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1715) begin
      mem_426_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1714) begin
      mem_425_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1713) begin
      mem_424_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1712) begin
      mem_423_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      mem_422_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1710) begin
      mem_421_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1709) begin
      mem_420_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1708) begin
      mem_419_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1707) begin
      mem_418_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1706) begin
      mem_417_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1705) begin
      mem_416_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1704) begin
      mem_415_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1703) begin
      mem_414_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      mem_413_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1701) begin
      mem_412_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1700) begin
      mem_411_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1699) begin
      mem_410_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1698) begin
      mem_409_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1697) begin
      mem_408_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1696) begin
      mem_407_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1695) begin
      mem_406_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1694) begin
      mem_405_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1693) begin
      mem_404_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1692) begin
      mem_403_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1691) begin
      mem_402_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1690) begin
      mem_401_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1689) begin
      mem_400_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      mem_399_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1687) begin
      mem_398_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1686) begin
      mem_397_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1685) begin
      mem_396_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1684) begin
      mem_395_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1683) begin
      mem_394_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1682) begin
      mem_393_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1681) begin
      mem_392_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1680) begin
      mem_391_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1679) begin
      mem_390_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1678) begin
      mem_389_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1677) begin
      mem_388_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1676) begin
      mem_387_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      mem_386_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1674) begin
      mem_385_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1673) begin
      mem_384_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1672) begin
      mem_383_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1671) begin
      mem_382_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1670) begin
      mem_381_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1669) begin
      mem_380_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1668) begin
      mem_379_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1667) begin
      mem_378_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1666) begin
      mem_377_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1665) begin
      mem_376_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      mem_375_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1663) begin
      mem_374_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      mem_373_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1661) begin
      mem_372_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1660) begin
      mem_371_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1659) begin
      mem_370_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1658) begin
      mem_369_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1657) begin
      mem_368_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1656) begin
      mem_367_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1655) begin
      mem_366_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1654) begin
      mem_365_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1653) begin
      mem_364_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1652) begin
      mem_363_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1651) begin
      mem_362_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1650) begin
      mem_361_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1649) begin
      mem_360_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1648) begin
      mem_359_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1647) begin
      mem_358_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1646) begin
      mem_357_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1645) begin
      mem_356_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1644) begin
      mem_355_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1643) begin
      mem_354_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1642) begin
      mem_353_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1641) begin
      mem_352_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1640) begin
      mem_351_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1639) begin
      mem_350_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1638) begin
      mem_349_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1637) begin
      mem_348_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1636) begin
      mem_347_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1635) begin
      mem_346_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1634) begin
      mem_345_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1633) begin
      mem_344_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1632) begin
      mem_343_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1631) begin
      mem_342_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1630) begin
      mem_341_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1629) begin
      mem_340_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1628) begin
      mem_339_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1627) begin
      mem_338_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1626) begin
      mem_337_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1625) begin
      mem_336_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1624) begin
      mem_335_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1623) begin
      mem_334_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1622) begin
      mem_333_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1621) begin
      mem_332_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1620) begin
      mem_331_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1619) begin
      mem_330_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1618) begin
      mem_329_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1617) begin
      mem_328_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1616) begin
      mem_327_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mem_326_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1614) begin
      mem_325_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1613) begin
      mem_324_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1612) begin
      mem_323_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1611) begin
      mem_322_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1610) begin
      mem_321_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1609) begin
      mem_320_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1608) begin
      mem_319_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1607) begin
      mem_318_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1606) begin
      mem_317_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1605) begin
      mem_316_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1604) begin
      mem_315_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1603) begin
      mem_314_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1602) begin
      mem_313_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1601) begin
      mem_312_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1600) begin
      mem_311_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1599) begin
      mem_310_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1598) begin
      mem_309_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1597) begin
      mem_308_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1596) begin
      mem_307_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1595) begin
      mem_306_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1594) begin
      mem_305_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1593) begin
      mem_304_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1592) begin
      mem_303_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1591) begin
      mem_302_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1590) begin
      mem_301_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1589) begin
      mem_300_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1588) begin
      mem_299_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1587) begin
      mem_298_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1586) begin
      mem_297_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1585) begin
      mem_296_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1584) begin
      mem_295_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1583) begin
      mem_294_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1582) begin
      mem_293_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1581) begin
      mem_292_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1580) begin
      mem_291_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1579) begin
      mem_290_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1578) begin
      mem_289_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1577) begin
      mem_288_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mem_287_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1575) begin
      mem_286_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1574) begin
      mem_285_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1573) begin
      mem_284_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1572) begin
      mem_283_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1571) begin
      mem_282_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1570) begin
      mem_281_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1569) begin
      mem_280_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1568) begin
      mem_279_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1567) begin
      mem_278_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1566) begin
      mem_277_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mem_276_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1564) begin
      mem_275_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1563) begin
      mem_274_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1562) begin
      mem_273_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1561) begin
      mem_272_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1560) begin
      mem_271_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1559) begin
      mem_270_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1558) begin
      mem_269_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1557) begin
      mem_268_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1556) begin
      mem_267_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1555) begin
      mem_266_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1554) begin
      mem_265_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1553) begin
      mem_264_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1552) begin
      mem_263_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1551) begin
      mem_262_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1550) begin
      mem_261_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1549) begin
      mem_260_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1548) begin
      mem_259_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1547) begin
      mem_258_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1546) begin
      mem_257_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1545) begin
      mem_256_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1544) begin
      mem_255_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1543) begin
      mem_254_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1542) begin
      mem_253_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1541) begin
      mem_252_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1540) begin
      mem_251_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1539) begin
      mem_250_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1538) begin
      mem_249_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1537) begin
      mem_248_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1536) begin
      mem_247_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1535) begin
      mem_246_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1534) begin
      mem_245_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1533) begin
      mem_244_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1532) begin
      mem_243_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1531) begin
      mem_242_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1530) begin
      mem_241_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1529) begin
      mem_240_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1528) begin
      mem_239_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1527) begin
      mem_238_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1526) begin
      mem_237_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1525) begin
      mem_236_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1524) begin
      mem_235_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1523) begin
      mem_234_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1522) begin
      mem_233_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1521) begin
      mem_232_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1520) begin
      mem_231_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1519) begin
      mem_230_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1518) begin
      mem_229_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1517) begin
      mem_228_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1516) begin
      mem_227_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1515) begin
      mem_226_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1514) begin
      mem_225_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1513) begin
      mem_224_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1512) begin
      mem_223_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1511) begin
      mem_222_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1510) begin
      mem_221_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1509) begin
      mem_220_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1508) begin
      mem_219_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1507) begin
      mem_218_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1506) begin
      mem_217_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1505) begin
      mem_216_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1504) begin
      mem_215_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1503) begin
      mem_214_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1502) begin
      mem_213_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1501) begin
      mem_212_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1500) begin
      mem_211_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1499) begin
      mem_210_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1498) begin
      mem_209_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1497) begin
      mem_208_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1496) begin
      mem_207_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1495) begin
      mem_206_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1494) begin
      mem_205_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1493) begin
      mem_204_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1492) begin
      mem_203_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1491) begin
      mem_202_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1490) begin
      mem_201_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1489) begin
      mem_200_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1488) begin
      mem_199_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1487) begin
      mem_198_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1486) begin
      mem_197_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1485) begin
      mem_196_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1484) begin
      mem_195_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1483) begin
      mem_194_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1482) begin
      mem_193_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1481) begin
      mem_192_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1480) begin
      mem_191_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1479) begin
      mem_190_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1478) begin
      mem_189_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1477) begin
      mem_188_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1476) begin
      mem_187_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1475) begin
      mem_186_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1474) begin
      mem_185_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1473) begin
      mem_184_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1472) begin
      mem_183_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1471) begin
      mem_182_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1470) begin
      mem_181_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1469) begin
      mem_180_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1468) begin
      mem_179_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1467) begin
      mem_178_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1466) begin
      mem_177_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1465) begin
      mem_176_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1464) begin
      mem_175_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1463) begin
      mem_174_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1462) begin
      mem_173_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1461) begin
      mem_172_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1460) begin
      mem_171_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1459) begin
      mem_170_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1458) begin
      mem_169_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1457) begin
      mem_168_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1456) begin
      mem_167_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1455) begin
      mem_166_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1454) begin
      mem_165_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1453) begin
      mem_164_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1452) begin
      mem_163_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1451) begin
      mem_162_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1450) begin
      mem_161_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1449) begin
      mem_160_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1448) begin
      mem_159_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1447) begin
      mem_158_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1446) begin
      mem_157_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1445) begin
      mem_156_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1444) begin
      mem_155_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1443) begin
      mem_154_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1442) begin
      mem_153_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1441) begin
      mem_152_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1440) begin
      mem_151_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1439) begin
      mem_150_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1438) begin
      mem_149_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1437) begin
      mem_148_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1436) begin
      mem_147_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1435) begin
      mem_146_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1434) begin
      mem_145_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1433) begin
      mem_144_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1432) begin
      mem_143_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1431) begin
      mem_142_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1430) begin
      mem_141_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1429) begin
      mem_140_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1428) begin
      mem_139_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1427) begin
      mem_138_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1426) begin
      mem_137_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1425) begin
      mem_136_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1424) begin
      mem_135_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1423) begin
      mem_134_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1422) begin
      mem_133_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1421) begin
      mem_132_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1420) begin
      mem_131_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1419) begin
      mem_130_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1418) begin
      mem_129_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1417) begin
      mem_128_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1416) begin
      mem_127_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1415) begin
      mem_126_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1414) begin
      mem_125_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1413) begin
      mem_124_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1412) begin
      mem_123_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1411) begin
      mem_122_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1410) begin
      mem_121_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1409) begin
      mem_120_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1408) begin
      mem_119_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1407) begin
      mem_118_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1406) begin
      mem_117_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1405) begin
      mem_116_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1404) begin
      mem_115_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1403) begin
      mem_114_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1402) begin
      mem_113_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1401) begin
      mem_112_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1400) begin
      mem_111_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1399) begin
      mem_110_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1398) begin
      mem_109_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1397) begin
      mem_108_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1396) begin
      mem_107_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1395) begin
      mem_106_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1394) begin
      mem_105_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1393) begin
      mem_104_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1392) begin
      mem_103_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1391) begin
      mem_102_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1390) begin
      mem_101_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1389) begin
      mem_100_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1388) begin
      mem_99_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1387) begin
      mem_98_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1386) begin
      mem_97_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1385) begin
      mem_96_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1384) begin
      mem_95_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1383) begin
      mem_94_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1382) begin
      mem_93_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1381) begin
      mem_92_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1380) begin
      mem_91_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1379) begin
      mem_90_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1378) begin
      mem_89_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1377) begin
      mem_88_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1376) begin
      mem_87_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1375) begin
      mem_86_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1374) begin
      mem_85_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1373) begin
      mem_84_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1372) begin
      mem_83_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1371) begin
      mem_82_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1370) begin
      mem_81_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1369) begin
      mem_80_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1368) begin
      mem_79_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1367) begin
      mem_78_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1366) begin
      mem_77_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1365) begin
      mem_76_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1364) begin
      mem_75_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1363) begin
      mem_74_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1362) begin
      mem_73_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1361) begin
      mem_72_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1360) begin
      mem_71_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1359) begin
      mem_70_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1358) begin
      mem_69_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1357) begin
      mem_68_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1356) begin
      mem_67_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1355) begin
      mem_66_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1354) begin
      mem_65_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1353) begin
      mem_64_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1352) begin
      mem_63_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1351) begin
      mem_62_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1350) begin
      mem_61_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1349) begin
      mem_60_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1348) begin
      mem_59_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1347) begin
      mem_58_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1346) begin
      mem_57_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1345) begin
      mem_56_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1344) begin
      mem_55_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1343) begin
      mem_54_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1342) begin
      mem_53_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1341) begin
      mem_52_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1340) begin
      mem_51_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1339) begin
      mem_50_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1338) begin
      mem_49_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1337) begin
      mem_48_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1336) begin
      mem_47_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1335) begin
      mem_46_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1334) begin
      mem_45_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1333) begin
      mem_44_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1332) begin
      mem_43_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1331) begin
      mem_42_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1330) begin
      mem_41_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1329) begin
      mem_40_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1328) begin
      mem_39_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1327) begin
      mem_38_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1326) begin
      mem_37_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1325) begin
      mem_36_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1324) begin
      mem_35_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1323) begin
      mem_34_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1322) begin
      mem_33_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1321) begin
      mem_32_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1320) begin
      mem_31_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1319) begin
      mem_30_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1318) begin
      mem_29_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1317) begin
      mem_28_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1316) begin
      mem_27_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1315) begin
      mem_26_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1314) begin
      mem_25_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1313) begin
      mem_24_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1312) begin
      mem_23_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1311) begin
      mem_22_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1310) begin
      mem_21_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1309) begin
      mem_20_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1308) begin
      mem_19_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1307) begin
      mem_18_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1306) begin
      mem_17_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1305) begin
      mem_16_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1304) begin
      mem_15_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1303) begin
      mem_14_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N1302) begin
      mem_13_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N1301) begin
      mem_12_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N1300) begin
      mem_11_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N1299) begin
      mem_10_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N1298) begin
      mem_9_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N1297) begin
      mem_8_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N1296) begin
      mem_7_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N1295) begin
      mem_6_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1294) begin
      mem_5_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1293) begin
      mem_4_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1292) begin
      mem_3_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1291) begin
      mem_2_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1290) begin
      mem_1_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1289) begin
      mem_0_sv2v_reg <= data_i[0];
    end 
  end

  assign N2249 = addr_i[5] & N2266;
  assign N2250 = addr_i[5] & N2267;
  assign N2251 = addr_i[5] & N2268;
  assign N2252 = addr_i[2] & N2279;
  assign N2253 = addr_i[2] & N2280;
  assign N2254 = addr_i[2] & N2281;
  assign N325 = N2249 & N2252;
  assign N324 = N2249 & N2253;
  assign N323 = N2249 & N2254;
  assign N322 = N2249 & N2286;
  assign N321 = N2249 & N2287;
  assign N320 = N2249 & N2288;
  assign N319 = N2249 & N2289;
  assign N318 = N2249 & N2290;
  assign N317 = N2250 & N2252;
  assign N316 = N2250 & N2253;
  assign N315 = N2250 & N2254;
  assign N314 = N2250 & N2286;
  assign N313 = N2250 & N2287;
  assign N312 = N2250 & N2288;
  assign N311 = N2250 & N2289;
  assign N310 = N2250 & N2290;
  assign N309 = N2251 & N2252;
  assign N308 = N2251 & N2253;
  assign N307 = N2251 & N2254;
  assign N306 = N2251 & N2286;
  assign N305 = N2251 & N2287;
  assign N304 = N2251 & N2288;
  assign N303 = N2251 & N2289;
  assign N302 = N2251 & N2290;
  assign N301 = N2273 & N2252;
  assign N300 = N2273 & N2253;
  assign N299 = N2273 & N2254;
  assign N298 = N2274 & N2252;
  assign N297 = N2274 & N2253;
  assign N296 = N2274 & N2254;
  assign N295 = N2275 & N2252;
  assign N294 = N2275 & N2253;
  assign N293 = N2275 & N2254;
  assign N292 = N2276 & N2252;
  assign N291 = N2276 & N2253;
  assign N290 = N2276 & N2254;
  assign N289 = N2277 & N2252;
  assign N288 = N2277 & N2253;
  assign N287 = N2277 & N2254;
  assign N2255 = addr_i[5] & N2269;
  assign N2256 = N2265 & N2266;
  assign N2257 = N2265 & N2267;
  assign N2258 = N2265 & N2268;
  assign N2259 = N2265 & N2269;
  assign N2260 = addr_i[2] & N2282;
  assign N2261 = N2278 & N2279;
  assign N2262 = N2278 & N2280;
  assign N2263 = N2278 & N2281;
  assign N2264 = N2278 & N2282;
  assign N1095 = N2270 & N2260;
  assign N1094 = N2270 & N2261;
  assign N1093 = N2270 & N2262;
  assign N1092 = N2270 & N2263;
  assign N1091 = N2270 & N2264;
  assign N1090 = N2271 & N2260;
  assign N1089 = N2271 & N2261;
  assign N1088 = N2271 & N2262;
  assign N1087 = N2271 & N2263;
  assign N1086 = N2271 & N2264;
  assign N1085 = N2272 & N2260;
  assign N1084 = N2272 & N2261;
  assign N1083 = N2272 & N2262;
  assign N1082 = N2272 & N2263;
  assign N1081 = N2272 & N2264;
  assign N1080 = N2255 & N2283;
  assign N1079 = N2255 & N2284;
  assign N1078 = N2255 & N2285;
  assign N1077 = N2255 & N2260;
  assign N1076 = N2255 & N2261;
  assign N1075 = N2255 & N2262;
  assign N1074 = N2255 & N2263;
  assign N1073 = N2255 & N2264;
  assign N1072 = N2256 & N2283;
  assign N1071 = N2256 & N2284;
  assign N1070 = N2256 & N2285;
  assign N1069 = N2256 & N2260;
  assign N1068 = N2256 & N2261;
  assign N1067 = N2256 & N2262;
  assign N1066 = N2256 & N2263;
  assign N1065 = N2256 & N2264;
  assign N1064 = N2257 & N2283;
  assign N1063 = N2257 & N2284;
  assign N1062 = N2257 & N2285;
  assign N1061 = N2257 & N2260;
  assign N1060 = N2257 & N2261;
  assign N1059 = N2257 & N2262;
  assign N1058 = N2257 & N2263;
  assign N1057 = N2257 & N2264;
  assign N1056 = N2258 & N2283;
  assign N1055 = N2258 & N2284;
  assign N1054 = N2258 & N2285;
  assign N1053 = N2258 & N2260;
  assign N1052 = N2258 & N2261;
  assign N1051 = N2258 & N2262;
  assign N1050 = N2258 & N2263;
  assign N1049 = N2258 & N2264;
  assign N1048 = N2259 & N2283;
  assign N1047 = N2259 & N2284;
  assign N1046 = N2259 & N2285;
  assign N1045 = N2259 & N2260;
  assign N1044 = N2259 & N2261;
  assign N1043 = N2259 & N2262;
  assign N1042 = N2259 & N2263;
  assign N1041 = N2259 & N2264;
  assign N2265 = ~addr_i[5];
  assign N2266 = addr_i[3] & addr_i[4];
  assign N2267 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N2268 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N2269 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N2270 = addr_i[5] & N2266;
  assign N2271 = addr_i[5] & N2267;
  assign N2272 = addr_i[5] & N2268;
  assign N2273 = addr_i[5] & N2269;
  assign N2274 = N2265 & N2266;
  assign N2275 = N2265 & N2267;
  assign N2276 = N2265 & N2268;
  assign N2277 = N2265 & N2269;
  assign N2278 = ~addr_i[2];
  assign N2279 = addr_i[0] & addr_i[1];
  assign N2280 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N2281 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N2282 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N2283 = addr_i[2] & N2279;
  assign N2284 = addr_i[2] & N2280;
  assign N2285 = addr_i[2] & N2281;
  assign N2286 = addr_i[2] & N2282;
  assign N2287 = N2278 & N2279;
  assign N2288 = N2278 & N2280;
  assign N2289 = N2278 & N2281;
  assign N2290 = N2278 & N2282;
  assign N1224 = N2270 & N2283;
  assign N1223 = N2270 & N2284;
  assign N1222 = N2270 & N2285;
  assign N1221 = N2270 & N2286;
  assign N1220 = N2270 & N2287;
  assign N1219 = N2270 & N2288;
  assign N1218 = N2270 & N2289;
  assign N1217 = N2270 & N2290;
  assign N1216 = N2271 & N2283;
  assign N1215 = N2271 & N2284;
  assign N1214 = N2271 & N2285;
  assign N1213 = N2271 & N2286;
  assign N1212 = N2271 & N2287;
  assign N1211 = N2271 & N2288;
  assign N1210 = N2271 & N2289;
  assign N1209 = N2271 & N2290;
  assign N1208 = N2272 & N2283;
  assign N1207 = N2272 & N2284;
  assign N1206 = N2272 & N2285;
  assign N1205 = N2272 & N2286;
  assign N1204 = N2272 & N2287;
  assign N1203 = N2272 & N2288;
  assign N1202 = N2272 & N2289;
  assign N1201 = N2272 & N2290;
  assign N1200 = N2273 & N2283;
  assign N1199 = N2273 & N2284;
  assign N1198 = N2273 & N2285;
  assign N1197 = N2273 & N2286;
  assign N1196 = N2273 & N2287;
  assign N1195 = N2273 & N2288;
  assign N1194 = N2273 & N2289;
  assign N1193 = N2273 & N2290;
  assign N1192 = N2274 & N2283;
  assign N1191 = N2274 & N2284;
  assign N1190 = N2274 & N2285;
  assign N1189 = N2274 & N2286;
  assign N1188 = N2274 & N2287;
  assign N1187 = N2274 & N2288;
  assign N1186 = N2274 & N2289;
  assign N1185 = N2274 & N2290;
  assign N1184 = N2275 & N2283;
  assign N1183 = N2275 & N2284;
  assign N1182 = N2275 & N2285;
  assign N1181 = N2275 & N2286;
  assign N1180 = N2275 & N2287;
  assign N1179 = N2275 & N2288;
  assign N1178 = N2275 & N2289;
  assign N1177 = N2275 & N2290;
  assign N1176 = N2276 & N2283;
  assign N1175 = N2276 & N2284;
  assign N1174 = N2276 & N2285;
  assign N1173 = N2276 & N2286;
  assign N1172 = N2276 & N2287;
  assign N1171 = N2276 & N2288;
  assign N1170 = N2276 & N2289;
  assign N1169 = N2276 & N2290;
  assign N1168 = N2277 & N2283;
  assign N1167 = N2277 & N2284;
  assign N1166 = N2277 & N2285;
  assign N1165 = N2277 & N2286;
  assign N1164 = N2277 & N2287;
  assign N1163 = N2277 & N2288;
  assign N1162 = N2277 & N2289;
  assign N1161 = N2277 & N2290;
  assign { N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157 } = (N8)? { N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N1197, N1196, N1195, N1194, N1193, N298, N297, N296, N1189, N1188, N1187, N1186, N1185, N295, N294, N293, N1181, N1180, N1179, N1178, N1177, N292, N291, N290, N1173, N1172, N1171, N1170, N1169, N289, N288, N287, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N156)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222 } = (N9)? { N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N1197, N1196, N1195, N1194, N1193, N298, N297, N296, N1189, N1188, N1187, N1186, N1185, N295, N294, N293, N1181, N1180, N1179, N1178, N1177, N292, N291, N290, N1173, N1172, N1171, N1170, N1169, N289, N288, N287, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N221)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326 } = (N10)? { N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N1197, N1196, N1195, N1194, N1193, N298, N297, N296, N1189, N1188, N1187, N1186, N1185, N295, N294, N293, N1181, N1180, N1179, N1178, N1177, N292, N291, N290, N1173, N1172, N1171, N1170, N1169, N289, N288, N287, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N286)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391 } = (N11)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N390)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456 } = (N12)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N455)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521 } = (N13)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N520)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586 } = (N14)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N585)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651 } = (N15)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N650)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = w_mask_i[7];
  assign { N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716 } = (N16)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N715)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_mask_i[8];
  assign { N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781 } = (N17)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N780)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = w_mask_i[9];
  assign { N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846 } = (N18)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N845)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = w_mask_i[10];
  assign { N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911 } = (N19)? { N1224, N1223, N1222, N1095, N1094, N1093, N1092, N1091, N1216, N1215, N1214, N1090, N1089, N1088, N1087, N1086, N1208, N1207, N1206, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N910)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = w_mask_i[11];
  assign { N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976 } = (N20)? { N1224, N1223, N1222, N1095, N1094, N1093, N1092, N1091, N1216, N1215, N1214, N1090, N1089, N1088, N1087, N1086, N1208, N1207, N1206, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N975)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = w_mask_i[12];
  assign { N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096 } = (N21)? { N1224, N1223, N1222, N1095, N1094, N1093, N1092, N1091, N1216, N1215, N1214, N1090, N1089, N1088, N1087, N1086, N1208, N1207, N1206, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1040)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = w_mask_i[13];
  assign { N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225 } = (N22)? { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1160)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = w_mask_i[14];
  assign { N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289 } = (N23)? { N1288, N1159, N1039, N974, N909, N844, N779, N714, N649, N584, N519, N454, N389, N285, N220, N1287, N1158, N1038, N973, N908, N843, N778, N713, N648, N583, N518, N453, N388, N284, N219, N1286, N1157, N1037, N972, N907, N842, N777, N712, N647, N582, N517, N452, N387, N283, N218, N1285, N1156, N1036, N971, N906, N841, N776, N711, N646, N581, N516, N451, N386, N282, N217, N1284, N1155, N1035, N970, N905, N840, N775, N710, N645, N580, N515, N450, N385, N281, N216, N1283, N1154, N1034, N969, N904, N839, N774, N709, N644, N579, N514, N449, N384, N280, N215, N1282, N1153, N1033, N968, N903, N838, N773, N708, N643, N578, N513, N448, N383, N279, N214, N1281, N1152, N1032, N967, N902, N837, N772, N707, N642, N577, N512, N447, N382, N278, N213, N1280, N1151, N1031, N966, N901, N836, N771, N706, N641, N576, N511, N446, N381, N277, N212, N1279, N1150, N1030, N965, N900, N835, N770, N705, N640, N575, N510, N445, N380, N276, N211, N1278, N1149, N1029, N964, N899, N834, N769, N704, N639, N574, N509, N444, N379, N275, N210, N1277, N1148, N1028, N963, N898, N833, N768, N703, N638, N573, N508, N443, N378, N274, N209, N1276, N1147, N1027, N962, N897, N832, N767, N702, N637, N572, N507, N442, N377, N273, N208, N1275, N1146, N1026, N961, N896, N831, N766, N701, N636, N571, N506, N441, N376, N272, N207, N1274, N1145, N1025, N960, N895, N830, N765, N700, N635, N570, N505, N440, N375, N271, N206, N1273, N1144, N1024, N959, N894, N829, N764, N699, N634, N569, N504, N439, N374, N270, N205, N1272, N1143, N1023, N958, N893, N828, N763, N698, N633, N568, N503, N438, N373, N269, N204, N1271, N1142, N1022, N957, N892, N827, N762, N697, N632, N567, N502, N437, N372, N268, N203, N1270, N1141, N1021, N956, N891, N826, N761, N696, N631, N566, N501, N436, N371, N267, N202, N1269, N1140, N1020, N955, N890, N825, N760, N695, N630, N565, N500, N435, N370, N266, N201, N1268, N1139, N1019, N954, N889, N824, N759, N694, N629, N564, N499, N434, N369, N265, N200, N1267, N1138, N1018, N953, N888, N823, N758, N693, N628, N563, N498, N433, N368, N264, N199, N1266, N1137, N1017, N952, N887, N822, N757, N692, N627, N562, N497, N432, N367, N263, N198, N1265, N1136, N1016, N951, N886, N821, N756, N691, N626, N561, N496, N431, N366, N262, N197, N1264, N1135, N1015, N950, N885, N820, N755, N690, N625, N560, N495, N430, N365, N261, N196, N1263, N1134, N1014, N949, N884, N819, N754, N689, N624, N559, N494, N429, N364, N260, N195, N1262, N1133, N1013, N948, N883, N818, N753, N688, N623, N558, N493, N428, N363, N259, N194, N1261, N1132, N1012, N947, N882, N817, N752, N687, N622, N557, N492, N427, N362, N258, N193, N1260, N1131, N1011, N946, N881, N816, N751, N686, N621, N556, N491, N426, N361, N257, N192, N1259, N1130, N1010, N945, N880, N815, N750, N685, N620, N555, N490, N425, N360, N256, N191, N1258, N1129, N1009, N944, N879, N814, N749, N684, N619, N554, N489, N424, N359, N255, N190, N1257, N1128, N1008, N943, N878, N813, N748, N683, N618, N553, N488, N423, N358, N254, N189, N1256, N1127, N1007, N942, N877, N812, N747, N682, N617, N552, N487, N422, N357, N253, N188, N1255, N1126, N1006, N941, N876, N811, N746, N681, N616, N551, N486, N421, N356, N252, N187, N1254, N1125, N1005, N940, N875, N810, N745, N680, N615, N550, N485, N420, N355, N251, N186, N1253, N1124, N1004, N939, N874, N809, N744, N679, N614, N549, N484, N419, N354, N250, N185, N1252, N1123, N1003, N938, N873, N808, N743, N678, N613, N548, N483, N418, N353, N249, N184, N1251, N1122, N1002, N937, N872, N807, N742, N677, N612, N547, N482, N417, N352, N248, N183, N1250, N1121, N1001, N936, N871, N806, N741, N676, N611, N546, N481, N416, N351, N247, N182, N1249, N1120, N1000, N935, N870, N805, N740, N675, N610, N545, N480, N415, N350, N246, N181, N1248, N1119, N999, N934, N869, N804, N739, N674, N609, N544, N479, N414, N349, N245, N180, N1247, N1118, N998, N933, N868, N803, N738, N673, N608, N543, N478, N413, N348, N244, N179, N1246, N1117, N997, N932, N867, N802, N737, N672, N607, N542, N477, N412, N347, N243, N178, N1245, N1116, N996, N931, N866, N801, N736, N671, N606, N541, N476, N411, N346, N242, N177, N1244, N1115, N995, N930, N865, N800, N735, N670, N605, N540, N475, N410, N345, N241, N176, N1243, N1114, N994, N929, N864, N799, N734, N669, N604, N539, N474, N409, N344, N240, N175, N1242, N1113, N993, N928, N863, N798, N733, N668, N603, N538, N473, N408, N343, N239, N174, N1241, N1112, N992, N927, N862, N797, N732, N667, N602, N537, N472, N407, N342, N238, N173, N1240, N1111, N991, N926, N861, N796, N731, N666, N601, N536, N471, N406, N341, N237, N172, N1239, N1110, N990, N925, N860, N795, N730, N665, N600, N535, N470, N405, N340, N236, N171, N1238, N1109, N989, N924, N859, N794, N729, N664, N599, N534, N469, N404, N339, N235, N170, N1237, N1108, N988, N923, N858, N793, N728, N663, N598, N533, N468, N403, N338, N234, N169, N1236, N1107, N987, N922, N857, N792, N727, N662, N597, N532, N467, N402, N337, N233, N168, N1235, N1106, N986, N921, N856, N791, N726, N661, N596, N531, N466, N401, N336, N232, N167, N1234, N1105, N985, N920, N855, N790, N725, N660, N595, N530, N465, N400, N335, N231, N166, N1233, N1104, N984, N919, N854, N789, N724, N659, N594, N529, N464, N399, N334, N230, N165, N1232, N1103, N983, N918, N853, N788, N723, N658, N593, N528, N463, N398, N333, N229, N164, N1231, N1102, N982, N917, N852, N787, N722, N657, N592, N527, N462, N397, N332, N228, N163, N1230, N1101, N981, N916, N851, N786, N721, N656, N591, N526, N461, N396, N331, N227, N162, N1229, N1100, N980, N915, N850, N785, N720, N655, N590, N525, N460, N395, N330, N226, N161, N1228, N1099, N979, N914, N849, N784, N719, N654, N589, N524, N459, N394, N329, N225, N160, N1227, N1098, N978, N913, N848, N783, N718, N653, N588, N523, N458, N393, N328, N224, N159, N1226, N1097, N977, N912, N847, N782, N717, N652, N587, N522, N457, N392, N327, N223, N158, N1225, N1096, N976, N911, N846, N781, N716, N651, N586, N521, N456, N391, N326, N222, N157 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N155)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = N154;
  assign N24 = ~addr_r[0];
  assign N25 = ~addr_r[1];
  assign N26 = N24 & N25;
  assign N27 = N24 & addr_r[1];
  assign N28 = addr_r[0] & N25;
  assign N29 = addr_r[0] & addr_r[1];
  assign N30 = ~addr_r[2];
  assign N31 = N26 & N30;
  assign N32 = N26 & addr_r[2];
  assign N33 = N28 & N30;
  assign N34 = N28 & addr_r[2];
  assign N35 = N27 & N30;
  assign N36 = N27 & addr_r[2];
  assign N37 = N29 & N30;
  assign N38 = N29 & addr_r[2];
  assign N39 = ~addr_r[3];
  assign N40 = N31 & N39;
  assign N41 = N31 & addr_r[3];
  assign N42 = N33 & N39;
  assign N43 = N33 & addr_r[3];
  assign N44 = N35 & N39;
  assign N45 = N35 & addr_r[3];
  assign N46 = N37 & N39;
  assign N47 = N37 & addr_r[3];
  assign N48 = N32 & N39;
  assign N49 = N32 & addr_r[3];
  assign N50 = N34 & N39;
  assign N51 = N34 & addr_r[3];
  assign N52 = N36 & N39;
  assign N53 = N36 & addr_r[3];
  assign N54 = N38 & N39;
  assign N55 = N38 & addr_r[3];
  assign N56 = ~addr_r[4];
  assign N57 = N40 & N56;
  assign N58 = N40 & addr_r[4];
  assign N59 = N42 & N56;
  assign N60 = N42 & addr_r[4];
  assign N61 = N44 & N56;
  assign N62 = N44 & addr_r[4];
  assign N63 = N46 & N56;
  assign N64 = N46 & addr_r[4];
  assign N65 = N48 & N56;
  assign N66 = N48 & addr_r[4];
  assign N67 = N50 & N56;
  assign N68 = N50 & addr_r[4];
  assign N69 = N52 & N56;
  assign N70 = N52 & addr_r[4];
  assign N71 = N54 & N56;
  assign N72 = N54 & addr_r[4];
  assign N73 = N41 & N56;
  assign N74 = N41 & addr_r[4];
  assign N75 = N43 & N56;
  assign N76 = N43 & addr_r[4];
  assign N77 = N45 & N56;
  assign N78 = N45 & addr_r[4];
  assign N79 = N47 & N56;
  assign N80 = N47 & addr_r[4];
  assign N81 = N49 & N56;
  assign N82 = N49 & addr_r[4];
  assign N83 = N51 & N56;
  assign N84 = N51 & addr_r[4];
  assign N85 = N53 & N56;
  assign N86 = N53 & addr_r[4];
  assign N87 = N55 & N56;
  assign N88 = N55 & addr_r[4];
  assign N89 = ~addr_r[5];
  assign N90 = N57 & N89;
  assign N91 = N57 & addr_r[5];
  assign N92 = N59 & N89;
  assign N93 = N59 & addr_r[5];
  assign N94 = N61 & N89;
  assign N95 = N61 & addr_r[5];
  assign N96 = N63 & N89;
  assign N97 = N63 & addr_r[5];
  assign N98 = N65 & N89;
  assign N99 = N65 & addr_r[5];
  assign N100 = N67 & N89;
  assign N101 = N67 & addr_r[5];
  assign N102 = N69 & N89;
  assign N103 = N69 & addr_r[5];
  assign N104 = N71 & N89;
  assign N105 = N71 & addr_r[5];
  assign N106 = N73 & N89;
  assign N107 = N73 & addr_r[5];
  assign N108 = N75 & N89;
  assign N109 = N75 & addr_r[5];
  assign N110 = N77 & N89;
  assign N111 = N77 & addr_r[5];
  assign N112 = N79 & N89;
  assign N113 = N79 & addr_r[5];
  assign N114 = N81 & N89;
  assign N115 = N81 & addr_r[5];
  assign N116 = N83 & N89;
  assign N117 = N83 & addr_r[5];
  assign N118 = N85 & N89;
  assign N119 = N85 & addr_r[5];
  assign N120 = N87 & N89;
  assign N121 = N87 & addr_r[5];
  assign N122 = N58 & N89;
  assign N123 = N58 & addr_r[5];
  assign N124 = N60 & N89;
  assign N125 = N60 & addr_r[5];
  assign N126 = N62 & N89;
  assign N127 = N62 & addr_r[5];
  assign N128 = N64 & N89;
  assign N129 = N64 & addr_r[5];
  assign N130 = N66 & N89;
  assign N131 = N66 & addr_r[5];
  assign N132 = N68 & N89;
  assign N133 = N68 & addr_r[5];
  assign N134 = N70 & N89;
  assign N135 = N70 & addr_r[5];
  assign N136 = N72 & N89;
  assign N137 = N72 & addr_r[5];
  assign N138 = N74 & N89;
  assign N139 = N74 & addr_r[5];
  assign N140 = N76 & N89;
  assign N141 = N76 & addr_r[5];
  assign N142 = N78 & N89;
  assign N143 = N78 & addr_r[5];
  assign N144 = N80 & N89;
  assign N145 = N80 & addr_r[5];
  assign N146 = N82 & N89;
  assign N147 = N82 & addr_r[5];
  assign N148 = N84 & N89;
  assign N149 = N84 & addr_r[5];
  assign N150 = N86 & N89;
  assign N151 = N86 & addr_r[5];
  assign N152 = N88 & N89;
  assign N153 = N88 & addr_r[5];
  assign N154 = v_i & w_i;
  assign N155 = ~N154;
  assign N156 = ~w_mask_i[0];
  assign N221 = ~w_mask_i[1];
  assign N286 = ~w_mask_i[2];
  assign N390 = ~w_mask_i[3];
  assign N455 = ~w_mask_i[4];
  assign N520 = ~w_mask_i[5];
  assign N585 = ~w_mask_i[6];
  assign N650 = ~w_mask_i[7];
  assign N715 = ~w_mask_i[8];
  assign N780 = ~w_mask_i[9];
  assign N845 = ~w_mask_i[10];
  assign N910 = ~w_mask_i[11];
  assign N975 = ~w_mask_i[12];
  assign N1040 = ~w_mask_i[13];
  assign N1160 = ~w_mask_i[14];

endmodule