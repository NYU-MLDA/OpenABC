module IntSyncCrossingSink_2( // @[:freechips.rocketchip.system.TinyConfig.fir@115330.2]
  input   auto_in_sync_0, // @[:freechips.rocketchip.system.TinyConfig.fir@115333.4]
  output  auto_out_0 // @[:freechips.rocketchip.system.TinyConfig.fir@115333.4]
);
  assign auto_out_0 = auto_in_sync_0; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@115342.4]
endmodule