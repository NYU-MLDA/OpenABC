module bsg_array_concentrate_static_5_62
(
  i,
  o
);

  input [185:0] i;
  output [123:0] o;
  wire [123:0] o;
  assign o[123] = i[185];
  assign o[122] = i[184];
  assign o[121] = i[183];
  assign o[120] = i[182];
  assign o[119] = i[181];
  assign o[118] = i[180];
  assign o[117] = i[179];
  assign o[116] = i[178];
  assign o[115] = i[177];
  assign o[114] = i[176];
  assign o[113] = i[175];
  assign o[112] = i[174];
  assign o[111] = i[173];
  assign o[110] = i[172];
  assign o[109] = i[171];
  assign o[108] = i[170];
  assign o[107] = i[169];
  assign o[106] = i[168];
  assign o[105] = i[167];
  assign o[104] = i[166];
  assign o[103] = i[165];
  assign o[102] = i[164];
  assign o[101] = i[163];
  assign o[100] = i[162];
  assign o[99] = i[161];
  assign o[98] = i[160];
  assign o[97] = i[159];
  assign o[96] = i[158];
  assign o[95] = i[157];
  assign o[94] = i[156];
  assign o[93] = i[155];
  assign o[92] = i[154];
  assign o[91] = i[153];
  assign o[90] = i[152];
  assign o[89] = i[151];
  assign o[88] = i[150];
  assign o[87] = i[149];
  assign o[86] = i[148];
  assign o[85] = i[147];
  assign o[84] = i[146];
  assign o[83] = i[145];
  assign o[82] = i[144];
  assign o[81] = i[143];
  assign o[80] = i[142];
  assign o[79] = i[141];
  assign o[78] = i[140];
  assign o[77] = i[139];
  assign o[76] = i[138];
  assign o[75] = i[137];
  assign o[74] = i[136];
  assign o[73] = i[135];
  assign o[72] = i[134];
  assign o[71] = i[133];
  assign o[70] = i[132];
  assign o[69] = i[131];
  assign o[68] = i[130];
  assign o[67] = i[129];
  assign o[66] = i[128];
  assign o[65] = i[127];
  assign o[64] = i[126];
  assign o[63] = i[125];
  assign o[62] = i[124];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule