module store_buffer
(
  clk_i,
  rst_ni,
  flush_i,
  no_st_pending_o,
  page_offset_i,
  page_offset_matches_o,
  commit_i,
  commit_ready_o,
  ready_o,
  valid_i,
  valid_without_flush_i,
  paddr_i,
  data_i,
  be_i,
  data_size_i,
  req_port_i,
  req_port_o
);

  input [11:0] page_offset_i;
  input [63:0] paddr_i;
  input [63:0] data_i;
  input [7:0] be_i;
  input [1:0] data_size_i;
  input [65:0] req_port_i;
  output [133:0] req_port_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input commit_i;
  input valid_i;
  input valid_without_flush_i;
  output no_st_pending_o;
  output page_offset_matches_o;
  output commit_ready_o;
  output ready_o;
  wire [133:0] req_port_o;
  wire no_st_pending_o,page_offset_matches_o,commit_ready_o,ready_o,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,N107,N108,N109,N110,N111,N112,N113,speculative_queue_n_3__valid_,
  speculative_queue_n_2__valid_,speculative_queue_n_1__valid_,
  speculative_queue_n_0__valid_,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,commit_queue_n_7__valid_,commit_queue_n_6__valid_,commit_queue_n_5__valid_,
  commit_queue_n_4__valid_,commit_queue_n_3__valid_,commit_queue_n_2__valid_,
  commit_queue_n_1__valid_,commit_queue_n_0__valid_,N258,N259,N260,N261,N262,N263,N264,
  N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,
  N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,
  N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,
  N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,
  N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,
  N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,
  N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
  N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,
  N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,
  N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,
  N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,
  N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
  N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,
  N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,
  N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,
  N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,
  N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,
  N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,
  N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,
  N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,
  N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N711,N712,N713,
  N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728;
  wire [1:0] speculative_write_pointer_n;
  wire [2:0] speculative_status_cnt_n;
  wire [3:0] commit_status_cnt_n;
  reg [1:0] speculative_write_pointer_q,speculative_read_pointer_q;
  reg [2:0] speculative_status_cnt_q,commit_write_pointer_q,commit_read_pointer_q;
  reg speculative_queue_q_3__address__55_,speculative_queue_q_3__address__54_,
  speculative_queue_q_3__address__53_,speculative_queue_q_3__address__52_,
  speculative_queue_q_3__address__51_,speculative_queue_q_3__address__50_,
  speculative_queue_q_3__address__49_,speculative_queue_q_3__address__48_,
  speculative_queue_q_3__address__47_,speculative_queue_q_3__address__46_,speculative_queue_q_3__address__45_,
  speculative_queue_q_3__address__44_,speculative_queue_q_3__address__43_,
  speculative_queue_q_3__address__42_,speculative_queue_q_3__address__41_,
  speculative_queue_q_3__address__40_,speculative_queue_q_3__address__39_,
  speculative_queue_q_3__address__38_,speculative_queue_q_3__address__37_,speculative_queue_q_3__address__36_,
  speculative_queue_q_3__address__35_,speculative_queue_q_3__address__34_,
  speculative_queue_q_3__address__33_,speculative_queue_q_3__address__32_,
  speculative_queue_q_3__address__31_,speculative_queue_q_3__address__30_,
  speculative_queue_q_3__address__29_,speculative_queue_q_3__address__28_,
  speculative_queue_q_3__address__27_,speculative_queue_q_3__address__26_,speculative_queue_q_3__address__25_,
  speculative_queue_q_3__address__24_,speculative_queue_q_3__address__23_,
  speculative_queue_q_3__address__22_,speculative_queue_q_3__address__21_,
  speculative_queue_q_3__address__20_,speculative_queue_q_3__address__19_,
  speculative_queue_q_3__address__18_,speculative_queue_q_3__address__17_,speculative_queue_q_3__address__16_,
  speculative_queue_q_3__address__15_,speculative_queue_q_3__address__14_,
  speculative_queue_q_3__address__13_,speculative_queue_q_3__address__12_,
  speculative_queue_q_3__address__11_,speculative_queue_q_3__address__10_,
  speculative_queue_q_3__address__9_,speculative_queue_q_3__address__8_,
  speculative_queue_q_3__address__7_,speculative_queue_q_3__address__6_,speculative_queue_q_3__address__5_,
  speculative_queue_q_3__address__4_,speculative_queue_q_3__address__3_,
  speculative_queue_q_3__address__2_,speculative_queue_q_3__address__1_,
  speculative_queue_q_3__address__0_,speculative_queue_q_3__data__63_,speculative_queue_q_3__data__62_,
  speculative_queue_q_3__data__61_,speculative_queue_q_3__data__60_,
  speculative_queue_q_3__data__59_,speculative_queue_q_3__data__58_,speculative_queue_q_3__data__57_,
  speculative_queue_q_3__data__56_,speculative_queue_q_3__data__55_,
  speculative_queue_q_3__data__54_,speculative_queue_q_3__data__53_,
  speculative_queue_q_3__data__52_,speculative_queue_q_3__data__51_,speculative_queue_q_3__data__50_,
  speculative_queue_q_3__data__49_,speculative_queue_q_3__data__48_,
  speculative_queue_q_3__data__47_,speculative_queue_q_3__data__46_,speculative_queue_q_3__data__45_,
  speculative_queue_q_3__data__44_,speculative_queue_q_3__data__43_,
  speculative_queue_q_3__data__42_,speculative_queue_q_3__data__41_,speculative_queue_q_3__data__40_,
  speculative_queue_q_3__data__39_,speculative_queue_q_3__data__38_,
  speculative_queue_q_3__data__37_,speculative_queue_q_3__data__36_,
  speculative_queue_q_3__data__35_,speculative_queue_q_3__data__34_,speculative_queue_q_3__data__33_,
  speculative_queue_q_3__data__32_,speculative_queue_q_3__data__31_,
  speculative_queue_q_3__data__30_,speculative_queue_q_3__data__29_,speculative_queue_q_3__data__28_,
  speculative_queue_q_3__data__27_,speculative_queue_q_3__data__26_,
  speculative_queue_q_3__data__25_,speculative_queue_q_3__data__24_,speculative_queue_q_3__data__23_,
  speculative_queue_q_3__data__22_,speculative_queue_q_3__data__21_,
  speculative_queue_q_3__data__20_,speculative_queue_q_3__data__19_,
  speculative_queue_q_3__data__18_,speculative_queue_q_3__data__17_,speculative_queue_q_3__data__16_,
  speculative_queue_q_3__data__15_,speculative_queue_q_3__data__14_,
  speculative_queue_q_3__data__13_,speculative_queue_q_3__data__12_,speculative_queue_q_3__data__11_,
  speculative_queue_q_3__data__10_,speculative_queue_q_3__data__9_,
  speculative_queue_q_3__data__8_,speculative_queue_q_3__data__7_,speculative_queue_q_3__data__6_,
  speculative_queue_q_3__data__5_,speculative_queue_q_3__data__4_,
  speculative_queue_q_3__data__3_,speculative_queue_q_3__data__2_,speculative_queue_q_3__data__1_,
  speculative_queue_q_3__data__0_,speculative_queue_q_3__be__7_,
  speculative_queue_q_3__be__6_,speculative_queue_q_3__be__5_,speculative_queue_q_3__be__4_,
  speculative_queue_q_3__be__3_,speculative_queue_q_3__be__2_,speculative_queue_q_3__be__1_,
  speculative_queue_q_3__be__0_,speculative_queue_q_3__data_size__1_,
  speculative_queue_q_3__data_size__0_,speculative_queue_q_3__valid_,
  speculative_queue_q_2__address__55_,speculative_queue_q_2__address__54_,speculative_queue_q_2__address__53_,
  speculative_queue_q_2__address__52_,speculative_queue_q_2__address__51_,
  speculative_queue_q_2__address__50_,speculative_queue_q_2__address__49_,
  speculative_queue_q_2__address__48_,speculative_queue_q_2__address__47_,
  speculative_queue_q_2__address__46_,speculative_queue_q_2__address__45_,
  speculative_queue_q_2__address__44_,speculative_queue_q_2__address__43_,speculative_queue_q_2__address__42_,
  speculative_queue_q_2__address__41_,speculative_queue_q_2__address__40_,
  speculative_queue_q_2__address__39_,speculative_queue_q_2__address__38_,
  speculative_queue_q_2__address__37_,speculative_queue_q_2__address__36_,
  speculative_queue_q_2__address__35_,speculative_queue_q_2__address__34_,speculative_queue_q_2__address__33_,
  speculative_queue_q_2__address__32_,speculative_queue_q_2__address__31_,
  speculative_queue_q_2__address__30_,speculative_queue_q_2__address__29_,
  speculative_queue_q_2__address__28_,speculative_queue_q_2__address__27_,
  speculative_queue_q_2__address__26_,speculative_queue_q_2__address__25_,
  speculative_queue_q_2__address__24_,speculative_queue_q_2__address__23_,speculative_queue_q_2__address__22_,
  speculative_queue_q_2__address__21_,speculative_queue_q_2__address__20_,
  speculative_queue_q_2__address__19_,speculative_queue_q_2__address__18_,
  speculative_queue_q_2__address__17_,speculative_queue_q_2__address__16_,
  speculative_queue_q_2__address__15_,speculative_queue_q_2__address__14_,speculative_queue_q_2__address__13_,
  speculative_queue_q_2__address__12_,speculative_queue_q_2__address__11_,
  speculative_queue_q_2__address__10_,speculative_queue_q_2__address__9_,
  speculative_queue_q_2__address__8_,speculative_queue_q_2__address__7_,
  speculative_queue_q_2__address__6_,speculative_queue_q_2__address__5_,speculative_queue_q_2__address__4_,
  speculative_queue_q_2__address__3_,speculative_queue_q_2__address__2_,
  speculative_queue_q_2__address__1_,speculative_queue_q_2__address__0_,
  speculative_queue_q_2__data__63_,speculative_queue_q_2__data__62_,speculative_queue_q_2__data__61_,
  speculative_queue_q_2__data__60_,speculative_queue_q_2__data__59_,
  speculative_queue_q_2__data__58_,speculative_queue_q_2__data__57_,
  speculative_queue_q_2__data__56_,speculative_queue_q_2__data__55_,speculative_queue_q_2__data__54_,
  speculative_queue_q_2__data__53_,speculative_queue_q_2__data__52_,
  speculative_queue_q_2__data__51_,speculative_queue_q_2__data__50_,speculative_queue_q_2__data__49_,
  speculative_queue_q_2__data__48_,speculative_queue_q_2__data__47_,
  speculative_queue_q_2__data__46_,speculative_queue_q_2__data__45_,speculative_queue_q_2__data__44_,
  speculative_queue_q_2__data__43_,speculative_queue_q_2__data__42_,
  speculative_queue_q_2__data__41_,speculative_queue_q_2__data__40_,
  speculative_queue_q_2__data__39_,speculative_queue_q_2__data__38_,speculative_queue_q_2__data__37_,
  speculative_queue_q_2__data__36_,speculative_queue_q_2__data__35_,
  speculative_queue_q_2__data__34_,speculative_queue_q_2__data__33_,speculative_queue_q_2__data__32_,
  speculative_queue_q_2__data__31_,speculative_queue_q_2__data__30_,
  speculative_queue_q_2__data__29_,speculative_queue_q_2__data__28_,speculative_queue_q_2__data__27_,
  speculative_queue_q_2__data__26_,speculative_queue_q_2__data__25_,
  speculative_queue_q_2__data__24_,speculative_queue_q_2__data__23_,
  speculative_queue_q_2__data__22_,speculative_queue_q_2__data__21_,speculative_queue_q_2__data__20_,
  speculative_queue_q_2__data__19_,speculative_queue_q_2__data__18_,
  speculative_queue_q_2__data__17_,speculative_queue_q_2__data__16_,speculative_queue_q_2__data__15_,
  speculative_queue_q_2__data__14_,speculative_queue_q_2__data__13_,
  speculative_queue_q_2__data__12_,speculative_queue_q_2__data__11_,speculative_queue_q_2__data__10_,
  speculative_queue_q_2__data__9_,speculative_queue_q_2__data__8_,
  speculative_queue_q_2__data__7_,speculative_queue_q_2__data__6_,speculative_queue_q_2__data__5_,
  speculative_queue_q_2__data__4_,speculative_queue_q_2__data__3_,
  speculative_queue_q_2__data__2_,speculative_queue_q_2__data__1_,speculative_queue_q_2__data__0_,
  speculative_queue_q_2__be__7_,speculative_queue_q_2__be__6_,
  speculative_queue_q_2__be__5_,speculative_queue_q_2__be__4_,speculative_queue_q_2__be__3_,
  speculative_queue_q_2__be__2_,speculative_queue_q_2__be__1_,speculative_queue_q_2__be__0_,
  speculative_queue_q_2__data_size__1_,speculative_queue_q_2__data_size__0_,
  speculative_queue_q_2__valid_,speculative_queue_q_1__address__55_,
  speculative_queue_q_1__address__54_,speculative_queue_q_1__address__53_,
  speculative_queue_q_1__address__52_,speculative_queue_q_1__address__51_,speculative_queue_q_1__address__50_,
  speculative_queue_q_1__address__49_,speculative_queue_q_1__address__48_,
  speculative_queue_q_1__address__47_,speculative_queue_q_1__address__46_,
  speculative_queue_q_1__address__45_,speculative_queue_q_1__address__44_,
  speculative_queue_q_1__address__43_,speculative_queue_q_1__address__42_,
  speculative_queue_q_1__address__41_,speculative_queue_q_1__address__40_,speculative_queue_q_1__address__39_,
  speculative_queue_q_1__address__38_,speculative_queue_q_1__address__37_,
  speculative_queue_q_1__address__36_,speculative_queue_q_1__address__35_,
  speculative_queue_q_1__address__34_,speculative_queue_q_1__address__33_,
  speculative_queue_q_1__address__32_,speculative_queue_q_1__address__31_,speculative_queue_q_1__address__30_,
  speculative_queue_q_1__address__29_,speculative_queue_q_1__address__28_,
  speculative_queue_q_1__address__27_,speculative_queue_q_1__address__26_,
  speculative_queue_q_1__address__25_,speculative_queue_q_1__address__24_,
  speculative_queue_q_1__address__23_,speculative_queue_q_1__address__22_,
  speculative_queue_q_1__address__21_,speculative_queue_q_1__address__20_,speculative_queue_q_1__address__19_,
  speculative_queue_q_1__address__18_,speculative_queue_q_1__address__17_,
  speculative_queue_q_1__address__16_,speculative_queue_q_1__address__15_,
  speculative_queue_q_1__address__14_,speculative_queue_q_1__address__13_,
  speculative_queue_q_1__address__12_,speculative_queue_q_1__address__11_,speculative_queue_q_1__address__10_,
  speculative_queue_q_1__address__9_,speculative_queue_q_1__address__8_,
  speculative_queue_q_1__address__7_,speculative_queue_q_1__address__6_,
  speculative_queue_q_1__address__5_,speculative_queue_q_1__address__4_,
  speculative_queue_q_1__address__3_,speculative_queue_q_1__address__2_,speculative_queue_q_1__address__1_,
  speculative_queue_q_1__address__0_,speculative_queue_q_1__data__63_,
  speculative_queue_q_1__data__62_,speculative_queue_q_1__data__61_,
  speculative_queue_q_1__data__60_,speculative_queue_q_1__data__59_,speculative_queue_q_1__data__58_,
  speculative_queue_q_1__data__57_,speculative_queue_q_1__data__56_,
  speculative_queue_q_1__data__55_,speculative_queue_q_1__data__54_,speculative_queue_q_1__data__53_,
  speculative_queue_q_1__data__52_,speculative_queue_q_1__data__51_,
  speculative_queue_q_1__data__50_,speculative_queue_q_1__data__49_,speculative_queue_q_1__data__48_,
  speculative_queue_q_1__data__47_,speculative_queue_q_1__data__46_,
  speculative_queue_q_1__data__45_,speculative_queue_q_1__data__44_,
  speculative_queue_q_1__data__43_,speculative_queue_q_1__data__42_,speculative_queue_q_1__data__41_,
  speculative_queue_q_1__data__40_,speculative_queue_q_1__data__39_,
  speculative_queue_q_1__data__38_,speculative_queue_q_1__data__37_,speculative_queue_q_1__data__36_,
  speculative_queue_q_1__data__35_,speculative_queue_q_1__data__34_,
  speculative_queue_q_1__data__33_,speculative_queue_q_1__data__32_,speculative_queue_q_1__data__31_,
  speculative_queue_q_1__data__30_,speculative_queue_q_1__data__29_,
  speculative_queue_q_1__data__28_,speculative_queue_q_1__data__27_,
  speculative_queue_q_1__data__26_,speculative_queue_q_1__data__25_,speculative_queue_q_1__data__24_,
  speculative_queue_q_1__data__23_,speculative_queue_q_1__data__22_,
  speculative_queue_q_1__data__21_,speculative_queue_q_1__data__20_,speculative_queue_q_1__data__19_,
  speculative_queue_q_1__data__18_,speculative_queue_q_1__data__17_,
  speculative_queue_q_1__data__16_,speculative_queue_q_1__data__15_,speculative_queue_q_1__data__14_,
  speculative_queue_q_1__data__13_,speculative_queue_q_1__data__12_,
  speculative_queue_q_1__data__11_,speculative_queue_q_1__data__10_,
  speculative_queue_q_1__data__9_,speculative_queue_q_1__data__8_,speculative_queue_q_1__data__7_,
  speculative_queue_q_1__data__6_,speculative_queue_q_1__data__5_,
  speculative_queue_q_1__data__4_,speculative_queue_q_1__data__3_,speculative_queue_q_1__data__2_,
  speculative_queue_q_1__data__1_,speculative_queue_q_1__data__0_,
  speculative_queue_q_1__be__7_,speculative_queue_q_1__be__6_,speculative_queue_q_1__be__5_,
  speculative_queue_q_1__be__4_,speculative_queue_q_1__be__3_,speculative_queue_q_1__be__2_,
  speculative_queue_q_1__be__1_,speculative_queue_q_1__be__0_,
  speculative_queue_q_1__data_size__1_,speculative_queue_q_1__data_size__0_,speculative_queue_q_1__valid_,
  speculative_queue_q_0__address__55_,speculative_queue_q_0__address__54_,
  speculative_queue_q_0__address__53_,speculative_queue_q_0__address__52_,
  speculative_queue_q_0__address__51_,speculative_queue_q_0__address__50_,
  speculative_queue_q_0__address__49_,speculative_queue_q_0__address__48_,speculative_queue_q_0__address__47_,
  speculative_queue_q_0__address__46_,speculative_queue_q_0__address__45_,
  speculative_queue_q_0__address__44_,speculative_queue_q_0__address__43_,
  speculative_queue_q_0__address__42_,speculative_queue_q_0__address__41_,
  speculative_queue_q_0__address__40_,speculative_queue_q_0__address__39_,
  speculative_queue_q_0__address__38_,speculative_queue_q_0__address__37_,speculative_queue_q_0__address__36_,
  speculative_queue_q_0__address__35_,speculative_queue_q_0__address__34_,
  speculative_queue_q_0__address__33_,speculative_queue_q_0__address__32_,
  speculative_queue_q_0__address__31_,speculative_queue_q_0__address__30_,
  speculative_queue_q_0__address__29_,speculative_queue_q_0__address__28_,speculative_queue_q_0__address__27_,
  speculative_queue_q_0__address__26_,speculative_queue_q_0__address__25_,
  speculative_queue_q_0__address__24_,speculative_queue_q_0__address__23_,
  speculative_queue_q_0__address__22_,speculative_queue_q_0__address__21_,
  speculative_queue_q_0__address__20_,speculative_queue_q_0__address__19_,
  speculative_queue_q_0__address__18_,speculative_queue_q_0__address__17_,speculative_queue_q_0__address__16_,
  speculative_queue_q_0__address__15_,speculative_queue_q_0__address__14_,
  speculative_queue_q_0__address__13_,speculative_queue_q_0__address__12_,
  speculative_queue_q_0__address__11_,speculative_queue_q_0__address__10_,
  speculative_queue_q_0__address__9_,speculative_queue_q_0__address__8_,speculative_queue_q_0__address__7_,
  speculative_queue_q_0__address__6_,speculative_queue_q_0__address__5_,
  speculative_queue_q_0__address__4_,speculative_queue_q_0__address__3_,
  speculative_queue_q_0__address__2_,speculative_queue_q_0__address__1_,
  speculative_queue_q_0__address__0_,speculative_queue_q_0__data__63_,speculative_queue_q_0__data__62_,
  speculative_queue_q_0__data__61_,speculative_queue_q_0__data__60_,
  speculative_queue_q_0__data__59_,speculative_queue_q_0__data__58_,speculative_queue_q_0__data__57_,
  speculative_queue_q_0__data__56_,speculative_queue_q_0__data__55_,
  speculative_queue_q_0__data__54_,speculative_queue_q_0__data__53_,speculative_queue_q_0__data__52_,
  speculative_queue_q_0__data__51_,speculative_queue_q_0__data__50_,
  speculative_queue_q_0__data__49_,speculative_queue_q_0__data__48_,
  speculative_queue_q_0__data__47_,speculative_queue_q_0__data__46_,speculative_queue_q_0__data__45_,
  speculative_queue_q_0__data__44_,speculative_queue_q_0__data__43_,
  speculative_queue_q_0__data__42_,speculative_queue_q_0__data__41_,speculative_queue_q_0__data__40_,
  speculative_queue_q_0__data__39_,speculative_queue_q_0__data__38_,
  speculative_queue_q_0__data__37_,speculative_queue_q_0__data__36_,speculative_queue_q_0__data__35_,
  speculative_queue_q_0__data__34_,speculative_queue_q_0__data__33_,
  speculative_queue_q_0__data__32_,speculative_queue_q_0__data__31_,
  speculative_queue_q_0__data__30_,speculative_queue_q_0__data__29_,speculative_queue_q_0__data__28_,
  speculative_queue_q_0__data__27_,speculative_queue_q_0__data__26_,
  speculative_queue_q_0__data__25_,speculative_queue_q_0__data__24_,speculative_queue_q_0__data__23_,
  speculative_queue_q_0__data__22_,speculative_queue_q_0__data__21_,
  speculative_queue_q_0__data__20_,speculative_queue_q_0__data__19_,speculative_queue_q_0__data__18_,
  speculative_queue_q_0__data__17_,speculative_queue_q_0__data__16_,
  speculative_queue_q_0__data__15_,speculative_queue_q_0__data__14_,
  speculative_queue_q_0__data__13_,speculative_queue_q_0__data__12_,speculative_queue_q_0__data__11_,
  speculative_queue_q_0__data__10_,speculative_queue_q_0__data__9_,
  speculative_queue_q_0__data__8_,speculative_queue_q_0__data__7_,speculative_queue_q_0__data__6_,
  speculative_queue_q_0__data__5_,speculative_queue_q_0__data__4_,
  speculative_queue_q_0__data__3_,speculative_queue_q_0__data__2_,speculative_queue_q_0__data__1_,
  speculative_queue_q_0__data__0_,speculative_queue_q_0__be__7_,
  speculative_queue_q_0__be__6_,speculative_queue_q_0__be__5_,speculative_queue_q_0__be__4_,
  speculative_queue_q_0__be__3_,speculative_queue_q_0__be__2_,speculative_queue_q_0__be__1_,
  speculative_queue_q_0__be__0_,speculative_queue_q_0__data_size__1_,
  speculative_queue_q_0__data_size__0_,speculative_queue_q_0__valid_,commit_queue_q_7__address__55_,
  commit_queue_q_7__address__54_,commit_queue_q_7__address__53_,
  commit_queue_q_7__address__52_,commit_queue_q_7__address__51_,commit_queue_q_7__address__50_,
  commit_queue_q_7__address__49_,commit_queue_q_7__address__48_,
  commit_queue_q_7__address__47_,commit_queue_q_7__address__46_,commit_queue_q_7__address__45_,
  commit_queue_q_7__address__44_,commit_queue_q_7__address__43_,
  commit_queue_q_7__address__42_,commit_queue_q_7__address__41_,commit_queue_q_7__address__40_,
  commit_queue_q_7__address__39_,commit_queue_q_7__address__38_,commit_queue_q_7__address__37_,
  commit_queue_q_7__address__36_,commit_queue_q_7__address__35_,
  commit_queue_q_7__address__34_,commit_queue_q_7__address__33_,commit_queue_q_7__address__32_,
  commit_queue_q_7__address__31_,commit_queue_q_7__address__30_,
  commit_queue_q_7__address__29_,commit_queue_q_7__address__28_,commit_queue_q_7__address__27_,
  commit_queue_q_7__address__26_,commit_queue_q_7__address__25_,commit_queue_q_7__address__24_,
  commit_queue_q_7__address__23_,commit_queue_q_7__address__22_,
  commit_queue_q_7__address__21_,commit_queue_q_7__address__20_,commit_queue_q_7__address__19_,
  commit_queue_q_7__address__18_,commit_queue_q_7__address__17_,
  commit_queue_q_7__address__16_,commit_queue_q_7__address__15_,commit_queue_q_7__address__14_,
  commit_queue_q_7__address__13_,commit_queue_q_7__address__12_,
  commit_queue_q_7__address__11_,commit_queue_q_7__address__10_,commit_queue_q_7__address__9_,
  commit_queue_q_7__address__8_,commit_queue_q_7__address__7_,commit_queue_q_7__address__6_,
  commit_queue_q_7__address__5_,commit_queue_q_7__address__4_,
  commit_queue_q_7__address__3_,commit_queue_q_7__address__2_,commit_queue_q_7__address__1_,
  commit_queue_q_7__address__0_,commit_queue_q_7__data__63_,commit_queue_q_7__data__62_,
  commit_queue_q_7__data__61_,commit_queue_q_7__data__60_,commit_queue_q_7__data__59_,
  commit_queue_q_7__data__58_,commit_queue_q_7__data__57_,commit_queue_q_7__data__56_,
  commit_queue_q_7__data__55_,commit_queue_q_7__data__54_,
  commit_queue_q_7__data__53_,commit_queue_q_7__data__52_,commit_queue_q_7__data__51_,
  commit_queue_q_7__data__50_,commit_queue_q_7__data__49_,commit_queue_q_7__data__48_,
  commit_queue_q_7__data__47_,commit_queue_q_7__data__46_,commit_queue_q_7__data__45_,
  commit_queue_q_7__data__44_,commit_queue_q_7__data__43_,commit_queue_q_7__data__42_,
  commit_queue_q_7__data__41_,commit_queue_q_7__data__40_,commit_queue_q_7__data__39_,
  commit_queue_q_7__data__38_,commit_queue_q_7__data__37_,commit_queue_q_7__data__36_,
  commit_queue_q_7__data__35_,commit_queue_q_7__data__34_,
  commit_queue_q_7__data__33_,commit_queue_q_7__data__32_,commit_queue_q_7__data__31_,
  commit_queue_q_7__data__30_,commit_queue_q_7__data__29_,commit_queue_q_7__data__28_,
  commit_queue_q_7__data__27_,commit_queue_q_7__data__26_,commit_queue_q_7__data__25_,
  commit_queue_q_7__data__24_,commit_queue_q_7__data__23_,commit_queue_q_7__data__22_,
  commit_queue_q_7__data__21_,commit_queue_q_7__data__20_,commit_queue_q_7__data__19_,
  commit_queue_q_7__data__18_,commit_queue_q_7__data__17_,commit_queue_q_7__data__16_,
  commit_queue_q_7__data__15_,commit_queue_q_7__data__14_,
  commit_queue_q_7__data__13_,commit_queue_q_7__data__12_,commit_queue_q_7__data__11_,
  commit_queue_q_7__data__10_,commit_queue_q_7__data__9_,commit_queue_q_7__data__8_,
  commit_queue_q_7__data__7_,commit_queue_q_7__data__6_,commit_queue_q_7__data__5_,
  commit_queue_q_7__data__4_,commit_queue_q_7__data__3_,commit_queue_q_7__data__2_,
  commit_queue_q_7__data__1_,commit_queue_q_7__data__0_,commit_queue_q_7__be__7_,
  commit_queue_q_7__be__6_,commit_queue_q_7__be__5_,commit_queue_q_7__be__4_,
  commit_queue_q_7__be__3_,commit_queue_q_7__be__2_,commit_queue_q_7__be__1_,commit_queue_q_7__be__0_,
  commit_queue_q_7__data_size__1_,commit_queue_q_7__data_size__0_,
  commit_queue_q_7__valid_,commit_queue_q_6__address__55_,commit_queue_q_6__address__54_,
  commit_queue_q_6__address__53_,commit_queue_q_6__address__52_,commit_queue_q_6__address__51_,
  commit_queue_q_6__address__50_,commit_queue_q_6__address__49_,
  commit_queue_q_6__address__48_,commit_queue_q_6__address__47_,commit_queue_q_6__address__46_,
  commit_queue_q_6__address__45_,commit_queue_q_6__address__44_,
  commit_queue_q_6__address__43_,commit_queue_q_6__address__42_,commit_queue_q_6__address__41_,
  commit_queue_q_6__address__40_,commit_queue_q_6__address__39_,
  commit_queue_q_6__address__38_,commit_queue_q_6__address__37_,commit_queue_q_6__address__36_,
  commit_queue_q_6__address__35_,commit_queue_q_6__address__34_,commit_queue_q_6__address__33_,
  commit_queue_q_6__address__32_,commit_queue_q_6__address__31_,
  commit_queue_q_6__address__30_,commit_queue_q_6__address__29_,commit_queue_q_6__address__28_,
  commit_queue_q_6__address__27_,commit_queue_q_6__address__26_,
  commit_queue_q_6__address__25_,commit_queue_q_6__address__24_,commit_queue_q_6__address__23_,
  commit_queue_q_6__address__22_,commit_queue_q_6__address__21_,
  commit_queue_q_6__address__20_,commit_queue_q_6__address__19_,commit_queue_q_6__address__18_,
  commit_queue_q_6__address__17_,commit_queue_q_6__address__16_,commit_queue_q_6__address__15_,
  commit_queue_q_6__address__14_,commit_queue_q_6__address__13_,
  commit_queue_q_6__address__12_,commit_queue_q_6__address__11_,commit_queue_q_6__address__10_,
  commit_queue_q_6__address__9_,commit_queue_q_6__address__8_,
  commit_queue_q_6__address__7_,commit_queue_q_6__address__6_,commit_queue_q_6__address__5_,
  commit_queue_q_6__address__4_,commit_queue_q_6__address__3_,commit_queue_q_6__address__2_,
  commit_queue_q_6__address__1_,commit_queue_q_6__address__0_,commit_queue_q_6__data__63_,
  commit_queue_q_6__data__62_,commit_queue_q_6__data__61_,
  commit_queue_q_6__data__60_,commit_queue_q_6__data__59_,commit_queue_q_6__data__58_,
  commit_queue_q_6__data__57_,commit_queue_q_6__data__56_,commit_queue_q_6__data__55_,
  commit_queue_q_6__data__54_,commit_queue_q_6__data__53_,commit_queue_q_6__data__52_,
  commit_queue_q_6__data__51_,commit_queue_q_6__data__50_,commit_queue_q_6__data__49_,
  commit_queue_q_6__data__48_,commit_queue_q_6__data__47_,commit_queue_q_6__data__46_,
  commit_queue_q_6__data__45_,commit_queue_q_6__data__44_,commit_queue_q_6__data__43_,
  commit_queue_q_6__data__42_,commit_queue_q_6__data__41_,
  commit_queue_q_6__data__40_,commit_queue_q_6__data__39_,commit_queue_q_6__data__38_,
  commit_queue_q_6__data__37_,commit_queue_q_6__data__36_,commit_queue_q_6__data__35_,
  commit_queue_q_6__data__34_,commit_queue_q_6__data__33_,commit_queue_q_6__data__32_,
  commit_queue_q_6__data__31_,commit_queue_q_6__data__30_,commit_queue_q_6__data__29_,
  commit_queue_q_6__data__28_,commit_queue_q_6__data__27_,commit_queue_q_6__data__26_,
  commit_queue_q_6__data__25_,commit_queue_q_6__data__24_,commit_queue_q_6__data__23_,
  commit_queue_q_6__data__22_,commit_queue_q_6__data__21_,
  commit_queue_q_6__data__20_,commit_queue_q_6__data__19_,commit_queue_q_6__data__18_,
  commit_queue_q_6__data__17_,commit_queue_q_6__data__16_,commit_queue_q_6__data__15_,
  commit_queue_q_6__data__14_,commit_queue_q_6__data__13_,commit_queue_q_6__data__12_,
  commit_queue_q_6__data__11_,commit_queue_q_6__data__10_,commit_queue_q_6__data__9_,
  commit_queue_q_6__data__8_,commit_queue_q_6__data__7_,commit_queue_q_6__data__6_,
  commit_queue_q_6__data__5_,commit_queue_q_6__data__4_,commit_queue_q_6__data__3_,
  commit_queue_q_6__data__2_,commit_queue_q_6__data__1_,commit_queue_q_6__data__0_,
  commit_queue_q_6__be__7_,commit_queue_q_6__be__6_,commit_queue_q_6__be__5_,
  commit_queue_q_6__be__4_,commit_queue_q_6__be__3_,commit_queue_q_6__be__2_,
  commit_queue_q_6__be__1_,commit_queue_q_6__be__0_,commit_queue_q_6__data_size__1_,
  commit_queue_q_6__data_size__0_,commit_queue_q_6__valid_,commit_queue_q_5__address__55_,
  commit_queue_q_5__address__54_,commit_queue_q_5__address__53_,
  commit_queue_q_5__address__52_,commit_queue_q_5__address__51_,commit_queue_q_5__address__50_,
  commit_queue_q_5__address__49_,commit_queue_q_5__address__48_,
  commit_queue_q_5__address__47_,commit_queue_q_5__address__46_,commit_queue_q_5__address__45_,
  commit_queue_q_5__address__44_,commit_queue_q_5__address__43_,commit_queue_q_5__address__42_,
  commit_queue_q_5__address__41_,commit_queue_q_5__address__40_,
  commit_queue_q_5__address__39_,commit_queue_q_5__address__38_,commit_queue_q_5__address__37_,
  commit_queue_q_5__address__36_,commit_queue_q_5__address__35_,
  commit_queue_q_5__address__34_,commit_queue_q_5__address__33_,commit_queue_q_5__address__32_,
  commit_queue_q_5__address__31_,commit_queue_q_5__address__30_,commit_queue_q_5__address__29_,
  commit_queue_q_5__address__28_,commit_queue_q_5__address__27_,
  commit_queue_q_5__address__26_,commit_queue_q_5__address__25_,commit_queue_q_5__address__24_,
  commit_queue_q_5__address__23_,commit_queue_q_5__address__22_,
  commit_queue_q_5__address__21_,commit_queue_q_5__address__20_,commit_queue_q_5__address__19_,
  commit_queue_q_5__address__18_,commit_queue_q_5__address__17_,
  commit_queue_q_5__address__16_,commit_queue_q_5__address__15_,commit_queue_q_5__address__14_,
  commit_queue_q_5__address__13_,commit_queue_q_5__address__12_,commit_queue_q_5__address__11_,
  commit_queue_q_5__address__10_,commit_queue_q_5__address__9_,
  commit_queue_q_5__address__8_,commit_queue_q_5__address__7_,commit_queue_q_5__address__6_,
  commit_queue_q_5__address__5_,commit_queue_q_5__address__4_,commit_queue_q_5__address__3_,
  commit_queue_q_5__address__2_,commit_queue_q_5__address__1_,
  commit_queue_q_5__address__0_,commit_queue_q_5__data__63_,commit_queue_q_5__data__62_,
  commit_queue_q_5__data__61_,commit_queue_q_5__data__60_,commit_queue_q_5__data__59_,
  commit_queue_q_5__data__58_,commit_queue_q_5__data__57_,commit_queue_q_5__data__56_,
  commit_queue_q_5__data__55_,commit_queue_q_5__data__54_,commit_queue_q_5__data__53_,
  commit_queue_q_5__data__52_,commit_queue_q_5__data__51_,commit_queue_q_5__data__50_,
  commit_queue_q_5__data__49_,commit_queue_q_5__data__48_,
  commit_queue_q_5__data__47_,commit_queue_q_5__data__46_,commit_queue_q_5__data__45_,
  commit_queue_q_5__data__44_,commit_queue_q_5__data__43_,commit_queue_q_5__data__42_,
  commit_queue_q_5__data__41_,commit_queue_q_5__data__40_,commit_queue_q_5__data__39_,
  commit_queue_q_5__data__38_,commit_queue_q_5__data__37_,commit_queue_q_5__data__36_,
  commit_queue_q_5__data__35_,commit_queue_q_5__data__34_,commit_queue_q_5__data__33_,
  commit_queue_q_5__data__32_,commit_queue_q_5__data__31_,commit_queue_q_5__data__30_,
  commit_queue_q_5__data__29_,commit_queue_q_5__data__28_,
  commit_queue_q_5__data__27_,commit_queue_q_5__data__26_,commit_queue_q_5__data__25_,
  commit_queue_q_5__data__24_,commit_queue_q_5__data__23_,commit_queue_q_5__data__22_,
  commit_queue_q_5__data__21_,commit_queue_q_5__data__20_,commit_queue_q_5__data__19_,
  commit_queue_q_5__data__18_,commit_queue_q_5__data__17_,commit_queue_q_5__data__16_,
  commit_queue_q_5__data__15_,commit_queue_q_5__data__14_,commit_queue_q_5__data__13_,
  commit_queue_q_5__data__12_,commit_queue_q_5__data__11_,commit_queue_q_5__data__10_,
  commit_queue_q_5__data__9_,commit_queue_q_5__data__8_,
  commit_queue_q_5__data__7_,commit_queue_q_5__data__6_,commit_queue_q_5__data__5_,
  commit_queue_q_5__data__4_,commit_queue_q_5__data__3_,commit_queue_q_5__data__2_,
  commit_queue_q_5__data__1_,commit_queue_q_5__data__0_,commit_queue_q_5__be__7_,commit_queue_q_5__be__6_,
  commit_queue_q_5__be__5_,commit_queue_q_5__be__4_,commit_queue_q_5__be__3_,
  commit_queue_q_5__be__2_,commit_queue_q_5__be__1_,commit_queue_q_5__be__0_,
  commit_queue_q_5__data_size__1_,commit_queue_q_5__data_size__0_,commit_queue_q_5__valid_,
  commit_queue_q_4__address__55_,commit_queue_q_4__address__54_,
  commit_queue_q_4__address__53_,commit_queue_q_4__address__52_,commit_queue_q_4__address__51_,
  commit_queue_q_4__address__50_,commit_queue_q_4__address__49_,
  commit_queue_q_4__address__48_,commit_queue_q_4__address__47_,commit_queue_q_4__address__46_,
  commit_queue_q_4__address__45_,commit_queue_q_4__address__44_,
  commit_queue_q_4__address__43_,commit_queue_q_4__address__42_,commit_queue_q_4__address__41_,
  commit_queue_q_4__address__40_,commit_queue_q_4__address__39_,commit_queue_q_4__address__38_,
  commit_queue_q_4__address__37_,commit_queue_q_4__address__36_,
  commit_queue_q_4__address__35_,commit_queue_q_4__address__34_,commit_queue_q_4__address__33_,
  commit_queue_q_4__address__32_,commit_queue_q_4__address__31_,
  commit_queue_q_4__address__30_,commit_queue_q_4__address__29_,commit_queue_q_4__address__28_,
  commit_queue_q_4__address__27_,commit_queue_q_4__address__26_,commit_queue_q_4__address__25_,
  commit_queue_q_4__address__24_,commit_queue_q_4__address__23_,
  commit_queue_q_4__address__22_,commit_queue_q_4__address__21_,commit_queue_q_4__address__20_,
  commit_queue_q_4__address__19_,commit_queue_q_4__address__18_,
  commit_queue_q_4__address__17_,commit_queue_q_4__address__16_,commit_queue_q_4__address__15_,
  commit_queue_q_4__address__14_,commit_queue_q_4__address__13_,
  commit_queue_q_4__address__12_,commit_queue_q_4__address__11_,commit_queue_q_4__address__10_,
  commit_queue_q_4__address__9_,commit_queue_q_4__address__8_,commit_queue_q_4__address__7_,
  commit_queue_q_4__address__6_,commit_queue_q_4__address__5_,
  commit_queue_q_4__address__4_,commit_queue_q_4__address__3_,commit_queue_q_4__address__2_,
  commit_queue_q_4__address__1_,commit_queue_q_4__address__0_,commit_queue_q_4__data__63_,
  commit_queue_q_4__data__62_,commit_queue_q_4__data__61_,commit_queue_q_4__data__60_,
  commit_queue_q_4__data__59_,commit_queue_q_4__data__58_,
  commit_queue_q_4__data__57_,commit_queue_q_4__data__56_,commit_queue_q_4__data__55_,
  commit_queue_q_4__data__54_,commit_queue_q_4__data__53_,commit_queue_q_4__data__52_,
  commit_queue_q_4__data__51_,commit_queue_q_4__data__50_,commit_queue_q_4__data__49_,
  commit_queue_q_4__data__48_,commit_queue_q_4__data__47_,commit_queue_q_4__data__46_,
  commit_queue_q_4__data__45_,commit_queue_q_4__data__44_,commit_queue_q_4__data__43_,
  commit_queue_q_4__data__42_,commit_queue_q_4__data__41_,commit_queue_q_4__data__40_,
  commit_queue_q_4__data__39_,commit_queue_q_4__data__38_,
  commit_queue_q_4__data__37_,commit_queue_q_4__data__36_,commit_queue_q_4__data__35_,
  commit_queue_q_4__data__34_,commit_queue_q_4__data__33_,commit_queue_q_4__data__32_,
  commit_queue_q_4__data__31_,commit_queue_q_4__data__30_,commit_queue_q_4__data__29_,
  commit_queue_q_4__data__28_,commit_queue_q_4__data__27_,commit_queue_q_4__data__26_,
  commit_queue_q_4__data__25_,commit_queue_q_4__data__24_,commit_queue_q_4__data__23_,
  commit_queue_q_4__data__22_,commit_queue_q_4__data__21_,commit_queue_q_4__data__20_,
  commit_queue_q_4__data__19_,commit_queue_q_4__data__18_,
  commit_queue_q_4__data__17_,commit_queue_q_4__data__16_,commit_queue_q_4__data__15_,
  commit_queue_q_4__data__14_,commit_queue_q_4__data__13_,commit_queue_q_4__data__12_,
  commit_queue_q_4__data__11_,commit_queue_q_4__data__10_,commit_queue_q_4__data__9_,
  commit_queue_q_4__data__8_,commit_queue_q_4__data__7_,commit_queue_q_4__data__6_,
  commit_queue_q_4__data__5_,commit_queue_q_4__data__4_,commit_queue_q_4__data__3_,
  commit_queue_q_4__data__2_,commit_queue_q_4__data__1_,commit_queue_q_4__data__0_,
  commit_queue_q_4__be__7_,commit_queue_q_4__be__6_,commit_queue_q_4__be__5_,
  commit_queue_q_4__be__4_,commit_queue_q_4__be__3_,commit_queue_q_4__be__2_,
  commit_queue_q_4__be__1_,commit_queue_q_4__be__0_,commit_queue_q_4__data_size__1_,
  commit_queue_q_4__data_size__0_,commit_queue_q_4__valid_,commit_queue_q_3__address__55_,
  commit_queue_q_3__address__54_,commit_queue_q_3__address__53_,commit_queue_q_3__address__52_,
  commit_queue_q_3__address__51_,commit_queue_q_3__address__50_,
  commit_queue_q_3__address__49_,commit_queue_q_3__address__48_,commit_queue_q_3__address__47_,
  commit_queue_q_3__address__46_,commit_queue_q_3__address__45_,
  commit_queue_q_3__address__44_,commit_queue_q_3__address__43_,commit_queue_q_3__address__42_,
  commit_queue_q_3__address__41_,commit_queue_q_3__address__40_,
  commit_queue_q_3__address__39_,commit_queue_q_3__address__38_,commit_queue_q_3__address__37_,
  commit_queue_q_3__address__36_,commit_queue_q_3__address__35_,commit_queue_q_3__address__34_,
  commit_queue_q_3__address__33_,commit_queue_q_3__address__32_,
  commit_queue_q_3__address__31_,commit_queue_q_3__address__30_,commit_queue_q_3__address__29_,
  commit_queue_q_3__address__28_,commit_queue_q_3__address__27_,
  commit_queue_q_3__address__26_,commit_queue_q_3__address__25_,commit_queue_q_3__address__24_,
  commit_queue_q_3__address__23_,commit_queue_q_3__address__22_,
  commit_queue_q_3__address__21_,commit_queue_q_3__address__20_,commit_queue_q_3__address__19_,
  commit_queue_q_3__address__18_,commit_queue_q_3__address__17_,commit_queue_q_3__address__16_,
  commit_queue_q_3__address__15_,commit_queue_q_3__address__14_,
  commit_queue_q_3__address__13_,commit_queue_q_3__address__12_,commit_queue_q_3__address__11_,
  commit_queue_q_3__address__10_,commit_queue_q_3__address__9_,
  commit_queue_q_3__address__8_,commit_queue_q_3__address__7_,commit_queue_q_3__address__6_,
  commit_queue_q_3__address__5_,commit_queue_q_3__address__4_,commit_queue_q_3__address__3_,
  commit_queue_q_3__address__2_,commit_queue_q_3__address__1_,
  commit_queue_q_3__address__0_,commit_queue_q_3__data__63_,commit_queue_q_3__data__62_,
  commit_queue_q_3__data__61_,commit_queue_q_3__data__60_,commit_queue_q_3__data__59_,
  commit_queue_q_3__data__58_,commit_queue_q_3__data__57_,commit_queue_q_3__data__56_,
  commit_queue_q_3__data__55_,commit_queue_q_3__data__54_,commit_queue_q_3__data__53_,
  commit_queue_q_3__data__52_,commit_queue_q_3__data__51_,commit_queue_q_3__data__50_,
  commit_queue_q_3__data__49_,commit_queue_q_3__data__48_,commit_queue_q_3__data__47_,
  commit_queue_q_3__data__46_,commit_queue_q_3__data__45_,
  commit_queue_q_3__data__44_,commit_queue_q_3__data__43_,commit_queue_q_3__data__42_,
  commit_queue_q_3__data__41_,commit_queue_q_3__data__40_,commit_queue_q_3__data__39_,
  commit_queue_q_3__data__38_,commit_queue_q_3__data__37_,commit_queue_q_3__data__36_,
  commit_queue_q_3__data__35_,commit_queue_q_3__data__34_,commit_queue_q_3__data__33_,
  commit_queue_q_3__data__32_,commit_queue_q_3__data__31_,commit_queue_q_3__data__30_,
  commit_queue_q_3__data__29_,commit_queue_q_3__data__28_,commit_queue_q_3__data__27_,
  commit_queue_q_3__data__26_,commit_queue_q_3__data__25_,
  commit_queue_q_3__data__24_,commit_queue_q_3__data__23_,commit_queue_q_3__data__22_,
  commit_queue_q_3__data__21_,commit_queue_q_3__data__20_,commit_queue_q_3__data__19_,
  commit_queue_q_3__data__18_,commit_queue_q_3__data__17_,commit_queue_q_3__data__16_,
  commit_queue_q_3__data__15_,commit_queue_q_3__data__14_,commit_queue_q_3__data__13_,
  commit_queue_q_3__data__12_,commit_queue_q_3__data__11_,commit_queue_q_3__data__10_,
  commit_queue_q_3__data__9_,commit_queue_q_3__data__8_,commit_queue_q_3__data__7_,
  commit_queue_q_3__data__6_,commit_queue_q_3__data__5_,commit_queue_q_3__data__4_,
  commit_queue_q_3__data__3_,commit_queue_q_3__data__2_,commit_queue_q_3__data__1_,
  commit_queue_q_3__data__0_,commit_queue_q_3__be__7_,commit_queue_q_3__be__6_,
  commit_queue_q_3__be__5_,commit_queue_q_3__be__4_,commit_queue_q_3__be__3_,
  commit_queue_q_3__be__2_,commit_queue_q_3__be__1_,commit_queue_q_3__be__0_,
  commit_queue_q_3__data_size__1_,commit_queue_q_3__data_size__0_,commit_queue_q_3__valid_,
  commit_queue_q_2__address__55_,commit_queue_q_2__address__54_,
  commit_queue_q_2__address__53_,commit_queue_q_2__address__52_,commit_queue_q_2__address__51_,
  commit_queue_q_2__address__50_,commit_queue_q_2__address__49_,
  commit_queue_q_2__address__48_,commit_queue_q_2__address__47_,commit_queue_q_2__address__46_,
  commit_queue_q_2__address__45_,commit_queue_q_2__address__44_,commit_queue_q_2__address__43_,
  commit_queue_q_2__address__42_,commit_queue_q_2__address__41_,
  commit_queue_q_2__address__40_,commit_queue_q_2__address__39_,commit_queue_q_2__address__38_,
  commit_queue_q_2__address__37_,commit_queue_q_2__address__36_,
  commit_queue_q_2__address__35_,commit_queue_q_2__address__34_,commit_queue_q_2__address__33_,
  commit_queue_q_2__address__32_,commit_queue_q_2__address__31_,commit_queue_q_2__address__30_,
  commit_queue_q_2__address__29_,commit_queue_q_2__address__28_,
  commit_queue_q_2__address__27_,commit_queue_q_2__address__26_,commit_queue_q_2__address__25_,
  commit_queue_q_2__address__24_,commit_queue_q_2__address__23_,
  commit_queue_q_2__address__22_,commit_queue_q_2__address__21_,commit_queue_q_2__address__20_,
  commit_queue_q_2__address__19_,commit_queue_q_2__address__18_,
  commit_queue_q_2__address__17_,commit_queue_q_2__address__16_,commit_queue_q_2__address__15_,
  commit_queue_q_2__address__14_,commit_queue_q_2__address__13_,commit_queue_q_2__address__12_,
  commit_queue_q_2__address__11_,commit_queue_q_2__address__10_,
  commit_queue_q_2__address__9_,commit_queue_q_2__address__8_,commit_queue_q_2__address__7_,
  commit_queue_q_2__address__6_,commit_queue_q_2__address__5_,commit_queue_q_2__address__4_,
  commit_queue_q_2__address__3_,commit_queue_q_2__address__2_,
  commit_queue_q_2__address__1_,commit_queue_q_2__address__0_,commit_queue_q_2__data__63_,
  commit_queue_q_2__data__62_,commit_queue_q_2__data__61_,commit_queue_q_2__data__60_,
  commit_queue_q_2__data__59_,commit_queue_q_2__data__58_,commit_queue_q_2__data__57_,
  commit_queue_q_2__data__56_,commit_queue_q_2__data__55_,commit_queue_q_2__data__54_,
  commit_queue_q_2__data__53_,commit_queue_q_2__data__52_,
  commit_queue_q_2__data__51_,commit_queue_q_2__data__50_,commit_queue_q_2__data__49_,
  commit_queue_q_2__data__48_,commit_queue_q_2__data__47_,commit_queue_q_2__data__46_,
  commit_queue_q_2__data__45_,commit_queue_q_2__data__44_,commit_queue_q_2__data__43_,
  commit_queue_q_2__data__42_,commit_queue_q_2__data__41_,commit_queue_q_2__data__40_,
  commit_queue_q_2__data__39_,commit_queue_q_2__data__38_,commit_queue_q_2__data__37_,
  commit_queue_q_2__data__36_,commit_queue_q_2__data__35_,commit_queue_q_2__data__34_,
  commit_queue_q_2__data__33_,commit_queue_q_2__data__32_,
  commit_queue_q_2__data__31_,commit_queue_q_2__data__30_,commit_queue_q_2__data__29_,
  commit_queue_q_2__data__28_,commit_queue_q_2__data__27_,commit_queue_q_2__data__26_,
  commit_queue_q_2__data__25_,commit_queue_q_2__data__24_,commit_queue_q_2__data__23_,
  commit_queue_q_2__data__22_,commit_queue_q_2__data__21_,commit_queue_q_2__data__20_,
  commit_queue_q_2__data__19_,commit_queue_q_2__data__18_,commit_queue_q_2__data__17_,
  commit_queue_q_2__data__16_,commit_queue_q_2__data__15_,commit_queue_q_2__data__14_,
  commit_queue_q_2__data__13_,commit_queue_q_2__data__12_,
  commit_queue_q_2__data__11_,commit_queue_q_2__data__10_,commit_queue_q_2__data__9_,
  commit_queue_q_2__data__8_,commit_queue_q_2__data__7_,commit_queue_q_2__data__6_,
  commit_queue_q_2__data__5_,commit_queue_q_2__data__4_,commit_queue_q_2__data__3_,
  commit_queue_q_2__data__2_,commit_queue_q_2__data__1_,commit_queue_q_2__data__0_,
  commit_queue_q_2__be__7_,commit_queue_q_2__be__6_,commit_queue_q_2__be__5_,
  commit_queue_q_2__be__4_,commit_queue_q_2__be__3_,commit_queue_q_2__be__2_,commit_queue_q_2__be__1_,
  commit_queue_q_2__be__0_,commit_queue_q_2__data_size__1_,
  commit_queue_q_2__data_size__0_,commit_queue_q_2__valid_,commit_queue_q_1__address__55_,
  commit_queue_q_1__address__54_,commit_queue_q_1__address__53_,commit_queue_q_1__address__52_,
  commit_queue_q_1__address__51_,commit_queue_q_1__address__50_,
  commit_queue_q_1__address__49_,commit_queue_q_1__address__48_,commit_queue_q_1__address__47_,
  commit_queue_q_1__address__46_,commit_queue_q_1__address__45_,
  commit_queue_q_1__address__44_,commit_queue_q_1__address__43_,commit_queue_q_1__address__42_,
  commit_queue_q_1__address__41_,commit_queue_q_1__address__40_,commit_queue_q_1__address__39_,
  commit_queue_q_1__address__38_,commit_queue_q_1__address__37_,
  commit_queue_q_1__address__36_,commit_queue_q_1__address__35_,commit_queue_q_1__address__34_,
  commit_queue_q_1__address__33_,commit_queue_q_1__address__32_,
  commit_queue_q_1__address__31_,commit_queue_q_1__address__30_,commit_queue_q_1__address__29_,
  commit_queue_q_1__address__28_,commit_queue_q_1__address__27_,commit_queue_q_1__address__26_,
  commit_queue_q_1__address__25_,commit_queue_q_1__address__24_,
  commit_queue_q_1__address__23_,commit_queue_q_1__address__22_,commit_queue_q_1__address__21_,
  commit_queue_q_1__address__20_,commit_queue_q_1__address__19_,
  commit_queue_q_1__address__18_,commit_queue_q_1__address__17_,commit_queue_q_1__address__16_,
  commit_queue_q_1__address__15_,commit_queue_q_1__address__14_,
  commit_queue_q_1__address__13_,commit_queue_q_1__address__12_,commit_queue_q_1__address__11_,
  commit_queue_q_1__address__10_,commit_queue_q_1__address__9_,commit_queue_q_1__address__8_,
  commit_queue_q_1__address__7_,commit_queue_q_1__address__6_,
  commit_queue_q_1__address__5_,commit_queue_q_1__address__4_,commit_queue_q_1__address__3_,
  commit_queue_q_1__address__2_,commit_queue_q_1__address__1_,commit_queue_q_1__address__0_,
  commit_queue_q_1__data__63_,commit_queue_q_1__data__62_,commit_queue_q_1__data__61_,
  commit_queue_q_1__data__60_,commit_queue_q_1__data__59_,
  commit_queue_q_1__data__58_,commit_queue_q_1__data__57_,commit_queue_q_1__data__56_,
  commit_queue_q_1__data__55_,commit_queue_q_1__data__54_,commit_queue_q_1__data__53_,
  commit_queue_q_1__data__52_,commit_queue_q_1__data__51_,commit_queue_q_1__data__50_,
  commit_queue_q_1__data__49_,commit_queue_q_1__data__48_,commit_queue_q_1__data__47_,
  commit_queue_q_1__data__46_,commit_queue_q_1__data__45_,commit_queue_q_1__data__44_,
  commit_queue_q_1__data__43_,commit_queue_q_1__data__42_,commit_queue_q_1__data__41_,
  commit_queue_q_1__data__40_,commit_queue_q_1__data__39_,
  commit_queue_q_1__data__38_,commit_queue_q_1__data__37_,commit_queue_q_1__data__36_,
  commit_queue_q_1__data__35_,commit_queue_q_1__data__34_,commit_queue_q_1__data__33_,
  commit_queue_q_1__data__32_,commit_queue_q_1__data__31_,commit_queue_q_1__data__30_,
  commit_queue_q_1__data__29_,commit_queue_q_1__data__28_,commit_queue_q_1__data__27_,
  commit_queue_q_1__data__26_,commit_queue_q_1__data__25_,commit_queue_q_1__data__24_,
  commit_queue_q_1__data__23_,commit_queue_q_1__data__22_,commit_queue_q_1__data__21_,
  commit_queue_q_1__data__20_,commit_queue_q_1__data__19_,
  commit_queue_q_1__data__18_,commit_queue_q_1__data__17_,commit_queue_q_1__data__16_,
  commit_queue_q_1__data__15_,commit_queue_q_1__data__14_,commit_queue_q_1__data__13_,
  commit_queue_q_1__data__12_,commit_queue_q_1__data__11_,commit_queue_q_1__data__10_,
  commit_queue_q_1__data__9_,commit_queue_q_1__data__8_,commit_queue_q_1__data__7_,
  commit_queue_q_1__data__6_,commit_queue_q_1__data__5_,commit_queue_q_1__data__4_,
  commit_queue_q_1__data__3_,commit_queue_q_1__data__2_,commit_queue_q_1__data__1_,
  commit_queue_q_1__data__0_,commit_queue_q_1__be__7_,commit_queue_q_1__be__6_,
  commit_queue_q_1__be__5_,commit_queue_q_1__be__4_,commit_queue_q_1__be__3_,
  commit_queue_q_1__be__2_,commit_queue_q_1__be__1_,commit_queue_q_1__be__0_,
  commit_queue_q_1__data_size__1_,commit_queue_q_1__data_size__0_,commit_queue_q_1__valid_,
  commit_queue_q_0__address__55_,commit_queue_q_0__address__54_,commit_queue_q_0__address__53_,
  commit_queue_q_0__address__52_,commit_queue_q_0__address__51_,
  commit_queue_q_0__address__50_,commit_queue_q_0__address__49_,commit_queue_q_0__address__48_,
  commit_queue_q_0__address__47_,commit_queue_q_0__address__46_,
  commit_queue_q_0__address__45_,commit_queue_q_0__address__44_,commit_queue_q_0__address__43_,
  commit_queue_q_0__address__42_,commit_queue_q_0__address__41_,
  commit_queue_q_0__address__40_,commit_queue_q_0__address__39_,commit_queue_q_0__address__38_,
  commit_queue_q_0__address__37_,commit_queue_q_0__address__36_,commit_queue_q_0__address__35_,
  commit_queue_q_0__address__34_,commit_queue_q_0__address__33_,
  commit_queue_q_0__address__32_,commit_queue_q_0__address__31_,commit_queue_q_0__address__30_,
  commit_queue_q_0__address__29_,commit_queue_q_0__address__28_,
  commit_queue_q_0__address__27_,commit_queue_q_0__address__26_,commit_queue_q_0__address__25_,
  commit_queue_q_0__address__24_,commit_queue_q_0__address__23_,
  commit_queue_q_0__address__22_,commit_queue_q_0__address__21_,commit_queue_q_0__address__20_,
  commit_queue_q_0__address__19_,commit_queue_q_0__address__18_,commit_queue_q_0__address__17_,
  commit_queue_q_0__address__16_,commit_queue_q_0__address__15_,
  commit_queue_q_0__address__14_,commit_queue_q_0__address__13_,commit_queue_q_0__address__12_,
  commit_queue_q_0__address__11_,commit_queue_q_0__address__10_,
  commit_queue_q_0__address__9_,commit_queue_q_0__address__8_,commit_queue_q_0__address__7_,
  commit_queue_q_0__address__6_,commit_queue_q_0__address__5_,commit_queue_q_0__address__4_,
  commit_queue_q_0__address__3_,commit_queue_q_0__address__2_,
  commit_queue_q_0__address__1_,commit_queue_q_0__address__0_,commit_queue_q_0__data__63_,
  commit_queue_q_0__data__62_,commit_queue_q_0__data__61_,commit_queue_q_0__data__60_,
  commit_queue_q_0__data__59_,commit_queue_q_0__data__58_,commit_queue_q_0__data__57_,
  commit_queue_q_0__data__56_,commit_queue_q_0__data__55_,commit_queue_q_0__data__54_,
  commit_queue_q_0__data__53_,commit_queue_q_0__data__52_,commit_queue_q_0__data__51_,
  commit_queue_q_0__data__50_,commit_queue_q_0__data__49_,
  commit_queue_q_0__data__48_,commit_queue_q_0__data__47_,commit_queue_q_0__data__46_,
  commit_queue_q_0__data__45_,commit_queue_q_0__data__44_,commit_queue_q_0__data__43_,
  commit_queue_q_0__data__42_,commit_queue_q_0__data__41_,commit_queue_q_0__data__40_,
  commit_queue_q_0__data__39_,commit_queue_q_0__data__38_,commit_queue_q_0__data__37_,
  commit_queue_q_0__data__36_,commit_queue_q_0__data__35_,commit_queue_q_0__data__34_,
  commit_queue_q_0__data__33_,commit_queue_q_0__data__32_,commit_queue_q_0__data__31_,
  commit_queue_q_0__data__30_,commit_queue_q_0__data__29_,
  commit_queue_q_0__data__28_,commit_queue_q_0__data__27_,commit_queue_q_0__data__26_,
  commit_queue_q_0__data__25_,commit_queue_q_0__data__24_,commit_queue_q_0__data__23_,
  commit_queue_q_0__data__22_,commit_queue_q_0__data__21_,commit_queue_q_0__data__20_,
  commit_queue_q_0__data__19_,commit_queue_q_0__data__18_,commit_queue_q_0__data__17_,
  commit_queue_q_0__data__16_,commit_queue_q_0__data__15_,commit_queue_q_0__data__14_,
  commit_queue_q_0__data__13_,commit_queue_q_0__data__12_,commit_queue_q_0__data__11_,
  commit_queue_q_0__data__10_,commit_queue_q_0__data__9_,commit_queue_q_0__data__8_,
  commit_queue_q_0__data__7_,commit_queue_q_0__data__6_,commit_queue_q_0__data__5_,
  commit_queue_q_0__data__4_,commit_queue_q_0__data__3_,
  commit_queue_q_0__data__2_,commit_queue_q_0__data__1_,commit_queue_q_0__data__0_,commit_queue_q_0__be__7_,
  commit_queue_q_0__be__6_,commit_queue_q_0__be__5_,commit_queue_q_0__be__4_,
  commit_queue_q_0__be__3_,commit_queue_q_0__be__2_,commit_queue_q_0__be__1_,
  commit_queue_q_0__be__0_,commit_queue_q_0__data_size__1_,commit_queue_q_0__data_size__0_,
  commit_queue_q_0__valid_;
  reg [3:0] commit_status_cnt_q;
  assign req_port_o[12] = 1'b1;
  assign req_port_o[0] = 1'b0;
  assign req_port_o[1] = 1'b0;
  assign N113 = speculative_status_cnt_q < { 1'b1, 1'b1 };
  assign req_port_o[133] = (N202)? commit_queue_q_0__address__11_ : 
                           (N204)? commit_queue_q_1__address__11_ : 
                           (N206)? commit_queue_q_2__address__11_ : 
                           (N208)? commit_queue_q_3__address__11_ : 
                           (N203)? commit_queue_q_4__address__11_ : 
                           (N205)? commit_queue_q_5__address__11_ : 
                           (N207)? commit_queue_q_6__address__11_ : 
                           (N209)? commit_queue_q_7__address__11_ : 1'b0;
  assign req_port_o[132] = (N202)? commit_queue_q_0__address__10_ : 
                           (N204)? commit_queue_q_1__address__10_ : 
                           (N206)? commit_queue_q_2__address__10_ : 
                           (N208)? commit_queue_q_3__address__10_ : 
                           (N203)? commit_queue_q_4__address__10_ : 
                           (N205)? commit_queue_q_5__address__10_ : 
                           (N207)? commit_queue_q_6__address__10_ : 
                           (N209)? commit_queue_q_7__address__10_ : 1'b0;
  assign req_port_o[131] = (N202)? commit_queue_q_0__address__9_ : 
                           (N204)? commit_queue_q_1__address__9_ : 
                           (N206)? commit_queue_q_2__address__9_ : 
                           (N208)? commit_queue_q_3__address__9_ : 
                           (N203)? commit_queue_q_4__address__9_ : 
                           (N205)? commit_queue_q_5__address__9_ : 
                           (N207)? commit_queue_q_6__address__9_ : 
                           (N209)? commit_queue_q_7__address__9_ : 1'b0;
  assign req_port_o[130] = (N202)? commit_queue_q_0__address__8_ : 
                           (N204)? commit_queue_q_1__address__8_ : 
                           (N206)? commit_queue_q_2__address__8_ : 
                           (N208)? commit_queue_q_3__address__8_ : 
                           (N203)? commit_queue_q_4__address__8_ : 
                           (N205)? commit_queue_q_5__address__8_ : 
                           (N207)? commit_queue_q_6__address__8_ : 
                           (N209)? commit_queue_q_7__address__8_ : 1'b0;
  assign req_port_o[129] = (N202)? commit_queue_q_0__address__7_ : 
                           (N204)? commit_queue_q_1__address__7_ : 
                           (N206)? commit_queue_q_2__address__7_ : 
                           (N208)? commit_queue_q_3__address__7_ : 
                           (N203)? commit_queue_q_4__address__7_ : 
                           (N205)? commit_queue_q_5__address__7_ : 
                           (N207)? commit_queue_q_6__address__7_ : 
                           (N209)? commit_queue_q_7__address__7_ : 1'b0;
  assign req_port_o[128] = (N202)? commit_queue_q_0__address__6_ : 
                           (N204)? commit_queue_q_1__address__6_ : 
                           (N206)? commit_queue_q_2__address__6_ : 
                           (N208)? commit_queue_q_3__address__6_ : 
                           (N203)? commit_queue_q_4__address__6_ : 
                           (N205)? commit_queue_q_5__address__6_ : 
                           (N207)? commit_queue_q_6__address__6_ : 
                           (N209)? commit_queue_q_7__address__6_ : 1'b0;
  assign req_port_o[127] = (N202)? commit_queue_q_0__address__5_ : 
                           (N204)? commit_queue_q_1__address__5_ : 
                           (N206)? commit_queue_q_2__address__5_ : 
                           (N208)? commit_queue_q_3__address__5_ : 
                           (N203)? commit_queue_q_4__address__5_ : 
                           (N205)? commit_queue_q_5__address__5_ : 
                           (N207)? commit_queue_q_6__address__5_ : 
                           (N209)? commit_queue_q_7__address__5_ : 1'b0;
  assign req_port_o[126] = (N202)? commit_queue_q_0__address__4_ : 
                           (N204)? commit_queue_q_1__address__4_ : 
                           (N206)? commit_queue_q_2__address__4_ : 
                           (N208)? commit_queue_q_3__address__4_ : 
                           (N203)? commit_queue_q_4__address__4_ : 
                           (N205)? commit_queue_q_5__address__4_ : 
                           (N207)? commit_queue_q_6__address__4_ : 
                           (N209)? commit_queue_q_7__address__4_ : 1'b0;
  assign req_port_o[125] = (N202)? commit_queue_q_0__address__3_ : 
                           (N204)? commit_queue_q_1__address__3_ : 
                           (N206)? commit_queue_q_2__address__3_ : 
                           (N208)? commit_queue_q_3__address__3_ : 
                           (N203)? commit_queue_q_4__address__3_ : 
                           (N205)? commit_queue_q_5__address__3_ : 
                           (N207)? commit_queue_q_6__address__3_ : 
                           (N209)? commit_queue_q_7__address__3_ : 1'b0;
  assign req_port_o[124] = (N202)? commit_queue_q_0__address__2_ : 
                           (N204)? commit_queue_q_1__address__2_ : 
                           (N206)? commit_queue_q_2__address__2_ : 
                           (N208)? commit_queue_q_3__address__2_ : 
                           (N203)? commit_queue_q_4__address__2_ : 
                           (N205)? commit_queue_q_5__address__2_ : 
                           (N207)? commit_queue_q_6__address__2_ : 
                           (N209)? commit_queue_q_7__address__2_ : 1'b0;
  assign req_port_o[123] = (N202)? commit_queue_q_0__address__1_ : 
                           (N204)? commit_queue_q_1__address__1_ : 
                           (N206)? commit_queue_q_2__address__1_ : 
                           (N208)? commit_queue_q_3__address__1_ : 
                           (N203)? commit_queue_q_4__address__1_ : 
                           (N205)? commit_queue_q_5__address__1_ : 
                           (N207)? commit_queue_q_6__address__1_ : 
                           (N209)? commit_queue_q_7__address__1_ : 1'b0;
  assign req_port_o[122] = (N202)? commit_queue_q_0__address__0_ : 
                           (N204)? commit_queue_q_1__address__0_ : 
                           (N206)? commit_queue_q_2__address__0_ : 
                           (N208)? commit_queue_q_3__address__0_ : 
                           (N203)? commit_queue_q_4__address__0_ : 
                           (N205)? commit_queue_q_5__address__0_ : 
                           (N207)? commit_queue_q_6__address__0_ : 
                           (N209)? commit_queue_q_7__address__0_ : 1'b0;
  assign req_port_o[121] = (N214)? commit_queue_q_0__address__55_ : 
                           (N216)? commit_queue_q_1__address__55_ : 
                           (N218)? commit_queue_q_2__address__55_ : 
                           (N220)? commit_queue_q_3__address__55_ : 
                           (N215)? commit_queue_q_4__address__55_ : 
                           (N217)? commit_queue_q_5__address__55_ : 
                           (N219)? commit_queue_q_6__address__55_ : 
                           (N221)? commit_queue_q_7__address__55_ : 1'b0;
  assign req_port_o[120] = (N214)? commit_queue_q_0__address__54_ : 
                           (N216)? commit_queue_q_1__address__54_ : 
                           (N218)? commit_queue_q_2__address__54_ : 
                           (N220)? commit_queue_q_3__address__54_ : 
                           (N215)? commit_queue_q_4__address__54_ : 
                           (N217)? commit_queue_q_5__address__54_ : 
                           (N219)? commit_queue_q_6__address__54_ : 
                           (N221)? commit_queue_q_7__address__54_ : 1'b0;
  assign req_port_o[119] = (N214)? commit_queue_q_0__address__53_ : 
                           (N216)? commit_queue_q_1__address__53_ : 
                           (N218)? commit_queue_q_2__address__53_ : 
                           (N220)? commit_queue_q_3__address__53_ : 
                           (N215)? commit_queue_q_4__address__53_ : 
                           (N217)? commit_queue_q_5__address__53_ : 
                           (N219)? commit_queue_q_6__address__53_ : 
                           (N221)? commit_queue_q_7__address__53_ : 1'b0;
  assign req_port_o[118] = (N214)? commit_queue_q_0__address__52_ : 
                           (N216)? commit_queue_q_1__address__52_ : 
                           (N218)? commit_queue_q_2__address__52_ : 
                           (N220)? commit_queue_q_3__address__52_ : 
                           (N215)? commit_queue_q_4__address__52_ : 
                           (N217)? commit_queue_q_5__address__52_ : 
                           (N219)? commit_queue_q_6__address__52_ : 
                           (N221)? commit_queue_q_7__address__52_ : 1'b0;
  assign req_port_o[117] = (N214)? commit_queue_q_0__address__51_ : 
                           (N216)? commit_queue_q_1__address__51_ : 
                           (N218)? commit_queue_q_2__address__51_ : 
                           (N220)? commit_queue_q_3__address__51_ : 
                           (N215)? commit_queue_q_4__address__51_ : 
                           (N217)? commit_queue_q_5__address__51_ : 
                           (N219)? commit_queue_q_6__address__51_ : 
                           (N221)? commit_queue_q_7__address__51_ : 1'b0;
  assign req_port_o[116] = (N214)? commit_queue_q_0__address__50_ : 
                           (N216)? commit_queue_q_1__address__50_ : 
                           (N218)? commit_queue_q_2__address__50_ : 
                           (N220)? commit_queue_q_3__address__50_ : 
                           (N215)? commit_queue_q_4__address__50_ : 
                           (N217)? commit_queue_q_5__address__50_ : 
                           (N219)? commit_queue_q_6__address__50_ : 
                           (N221)? commit_queue_q_7__address__50_ : 1'b0;
  assign req_port_o[115] = (N214)? commit_queue_q_0__address__49_ : 
                           (N216)? commit_queue_q_1__address__49_ : 
                           (N218)? commit_queue_q_2__address__49_ : 
                           (N220)? commit_queue_q_3__address__49_ : 
                           (N215)? commit_queue_q_4__address__49_ : 
                           (N217)? commit_queue_q_5__address__49_ : 
                           (N219)? commit_queue_q_6__address__49_ : 
                           (N221)? commit_queue_q_7__address__49_ : 1'b0;
  assign req_port_o[114] = (N214)? commit_queue_q_0__address__48_ : 
                           (N216)? commit_queue_q_1__address__48_ : 
                           (N218)? commit_queue_q_2__address__48_ : 
                           (N220)? commit_queue_q_3__address__48_ : 
                           (N215)? commit_queue_q_4__address__48_ : 
                           (N217)? commit_queue_q_5__address__48_ : 
                           (N219)? commit_queue_q_6__address__48_ : 
                           (N221)? commit_queue_q_7__address__48_ : 1'b0;
  assign req_port_o[113] = (N214)? commit_queue_q_0__address__47_ : 
                           (N216)? commit_queue_q_1__address__47_ : 
                           (N218)? commit_queue_q_2__address__47_ : 
                           (N220)? commit_queue_q_3__address__47_ : 
                           (N215)? commit_queue_q_4__address__47_ : 
                           (N217)? commit_queue_q_5__address__47_ : 
                           (N219)? commit_queue_q_6__address__47_ : 
                           (N221)? commit_queue_q_7__address__47_ : 1'b0;
  assign req_port_o[112] = (N214)? commit_queue_q_0__address__46_ : 
                           (N216)? commit_queue_q_1__address__46_ : 
                           (N218)? commit_queue_q_2__address__46_ : 
                           (N220)? commit_queue_q_3__address__46_ : 
                           (N215)? commit_queue_q_4__address__46_ : 
                           (N217)? commit_queue_q_5__address__46_ : 
                           (N219)? commit_queue_q_6__address__46_ : 
                           (N221)? commit_queue_q_7__address__46_ : 1'b0;
  assign req_port_o[111] = (N214)? commit_queue_q_0__address__45_ : 
                           (N216)? commit_queue_q_1__address__45_ : 
                           (N218)? commit_queue_q_2__address__45_ : 
                           (N220)? commit_queue_q_3__address__45_ : 
                           (N215)? commit_queue_q_4__address__45_ : 
                           (N217)? commit_queue_q_5__address__45_ : 
                           (N219)? commit_queue_q_6__address__45_ : 
                           (N221)? commit_queue_q_7__address__45_ : 1'b0;
  assign req_port_o[110] = (N214)? commit_queue_q_0__address__44_ : 
                           (N216)? commit_queue_q_1__address__44_ : 
                           (N218)? commit_queue_q_2__address__44_ : 
                           (N220)? commit_queue_q_3__address__44_ : 
                           (N215)? commit_queue_q_4__address__44_ : 
                           (N217)? commit_queue_q_5__address__44_ : 
                           (N219)? commit_queue_q_6__address__44_ : 
                           (N221)? commit_queue_q_7__address__44_ : 1'b0;
  assign req_port_o[109] = (N214)? commit_queue_q_0__address__43_ : 
                           (N216)? commit_queue_q_1__address__43_ : 
                           (N218)? commit_queue_q_2__address__43_ : 
                           (N220)? commit_queue_q_3__address__43_ : 
                           (N215)? commit_queue_q_4__address__43_ : 
                           (N217)? commit_queue_q_5__address__43_ : 
                           (N219)? commit_queue_q_6__address__43_ : 
                           (N221)? commit_queue_q_7__address__43_ : 1'b0;
  assign req_port_o[108] = (N214)? commit_queue_q_0__address__42_ : 
                           (N216)? commit_queue_q_1__address__42_ : 
                           (N218)? commit_queue_q_2__address__42_ : 
                           (N220)? commit_queue_q_3__address__42_ : 
                           (N215)? commit_queue_q_4__address__42_ : 
                           (N217)? commit_queue_q_5__address__42_ : 
                           (N219)? commit_queue_q_6__address__42_ : 
                           (N221)? commit_queue_q_7__address__42_ : 1'b0;
  assign req_port_o[107] = (N214)? commit_queue_q_0__address__41_ : 
                           (N216)? commit_queue_q_1__address__41_ : 
                           (N218)? commit_queue_q_2__address__41_ : 
                           (N220)? commit_queue_q_3__address__41_ : 
                           (N215)? commit_queue_q_4__address__41_ : 
                           (N217)? commit_queue_q_5__address__41_ : 
                           (N219)? commit_queue_q_6__address__41_ : 
                           (N221)? commit_queue_q_7__address__41_ : 1'b0;
  assign req_port_o[106] = (N214)? commit_queue_q_0__address__40_ : 
                           (N216)? commit_queue_q_1__address__40_ : 
                           (N218)? commit_queue_q_2__address__40_ : 
                           (N220)? commit_queue_q_3__address__40_ : 
                           (N215)? commit_queue_q_4__address__40_ : 
                           (N217)? commit_queue_q_5__address__40_ : 
                           (N219)? commit_queue_q_6__address__40_ : 
                           (N221)? commit_queue_q_7__address__40_ : 1'b0;
  assign req_port_o[105] = (N214)? commit_queue_q_0__address__39_ : 
                           (N216)? commit_queue_q_1__address__39_ : 
                           (N218)? commit_queue_q_2__address__39_ : 
                           (N220)? commit_queue_q_3__address__39_ : 
                           (N215)? commit_queue_q_4__address__39_ : 
                           (N217)? commit_queue_q_5__address__39_ : 
                           (N219)? commit_queue_q_6__address__39_ : 
                           (N221)? commit_queue_q_7__address__39_ : 1'b0;
  assign req_port_o[104] = (N214)? commit_queue_q_0__address__38_ : 
                           (N216)? commit_queue_q_1__address__38_ : 
                           (N218)? commit_queue_q_2__address__38_ : 
                           (N220)? commit_queue_q_3__address__38_ : 
                           (N215)? commit_queue_q_4__address__38_ : 
                           (N217)? commit_queue_q_5__address__38_ : 
                           (N219)? commit_queue_q_6__address__38_ : 
                           (N221)? commit_queue_q_7__address__38_ : 1'b0;
  assign req_port_o[103] = (N214)? commit_queue_q_0__address__37_ : 
                           (N216)? commit_queue_q_1__address__37_ : 
                           (N218)? commit_queue_q_2__address__37_ : 
                           (N220)? commit_queue_q_3__address__37_ : 
                           (N215)? commit_queue_q_4__address__37_ : 
                           (N217)? commit_queue_q_5__address__37_ : 
                           (N219)? commit_queue_q_6__address__37_ : 
                           (N221)? commit_queue_q_7__address__37_ : 1'b0;
  assign req_port_o[102] = (N214)? commit_queue_q_0__address__36_ : 
                           (N216)? commit_queue_q_1__address__36_ : 
                           (N218)? commit_queue_q_2__address__36_ : 
                           (N220)? commit_queue_q_3__address__36_ : 
                           (N215)? commit_queue_q_4__address__36_ : 
                           (N217)? commit_queue_q_5__address__36_ : 
                           (N219)? commit_queue_q_6__address__36_ : 
                           (N221)? commit_queue_q_7__address__36_ : 1'b0;
  assign req_port_o[101] = (N214)? commit_queue_q_0__address__35_ : 
                           (N216)? commit_queue_q_1__address__35_ : 
                           (N218)? commit_queue_q_2__address__35_ : 
                           (N220)? commit_queue_q_3__address__35_ : 
                           (N215)? commit_queue_q_4__address__35_ : 
                           (N217)? commit_queue_q_5__address__35_ : 
                           (N219)? commit_queue_q_6__address__35_ : 
                           (N221)? commit_queue_q_7__address__35_ : 1'b0;
  assign req_port_o[100] = (N214)? commit_queue_q_0__address__34_ : 
                           (N216)? commit_queue_q_1__address__34_ : 
                           (N218)? commit_queue_q_2__address__34_ : 
                           (N220)? commit_queue_q_3__address__34_ : 
                           (N215)? commit_queue_q_4__address__34_ : 
                           (N217)? commit_queue_q_5__address__34_ : 
                           (N219)? commit_queue_q_6__address__34_ : 
                           (N221)? commit_queue_q_7__address__34_ : 1'b0;
  assign req_port_o[99] = (N214)? commit_queue_q_0__address__33_ : 
                          (N216)? commit_queue_q_1__address__33_ : 
                          (N218)? commit_queue_q_2__address__33_ : 
                          (N220)? commit_queue_q_3__address__33_ : 
                          (N215)? commit_queue_q_4__address__33_ : 
                          (N217)? commit_queue_q_5__address__33_ : 
                          (N219)? commit_queue_q_6__address__33_ : 
                          (N221)? commit_queue_q_7__address__33_ : 1'b0;
  assign req_port_o[98] = (N214)? commit_queue_q_0__address__32_ : 
                          (N216)? commit_queue_q_1__address__32_ : 
                          (N218)? commit_queue_q_2__address__32_ : 
                          (N220)? commit_queue_q_3__address__32_ : 
                          (N215)? commit_queue_q_4__address__32_ : 
                          (N217)? commit_queue_q_5__address__32_ : 
                          (N219)? commit_queue_q_6__address__32_ : 
                          (N221)? commit_queue_q_7__address__32_ : 1'b0;
  assign req_port_o[97] = (N214)? commit_queue_q_0__address__31_ : 
                          (N216)? commit_queue_q_1__address__31_ : 
                          (N218)? commit_queue_q_2__address__31_ : 
                          (N220)? commit_queue_q_3__address__31_ : 
                          (N215)? commit_queue_q_4__address__31_ : 
                          (N217)? commit_queue_q_5__address__31_ : 
                          (N219)? commit_queue_q_6__address__31_ : 
                          (N221)? commit_queue_q_7__address__31_ : 1'b0;
  assign req_port_o[96] = (N214)? commit_queue_q_0__address__30_ : 
                          (N216)? commit_queue_q_1__address__30_ : 
                          (N218)? commit_queue_q_2__address__30_ : 
                          (N220)? commit_queue_q_3__address__30_ : 
                          (N215)? commit_queue_q_4__address__30_ : 
                          (N217)? commit_queue_q_5__address__30_ : 
                          (N219)? commit_queue_q_6__address__30_ : 
                          (N221)? commit_queue_q_7__address__30_ : 1'b0;
  assign req_port_o[95] = (N214)? commit_queue_q_0__address__29_ : 
                          (N216)? commit_queue_q_1__address__29_ : 
                          (N218)? commit_queue_q_2__address__29_ : 
                          (N220)? commit_queue_q_3__address__29_ : 
                          (N215)? commit_queue_q_4__address__29_ : 
                          (N217)? commit_queue_q_5__address__29_ : 
                          (N219)? commit_queue_q_6__address__29_ : 
                          (N221)? commit_queue_q_7__address__29_ : 1'b0;
  assign req_port_o[94] = (N214)? commit_queue_q_0__address__28_ : 
                          (N216)? commit_queue_q_1__address__28_ : 
                          (N218)? commit_queue_q_2__address__28_ : 
                          (N220)? commit_queue_q_3__address__28_ : 
                          (N215)? commit_queue_q_4__address__28_ : 
                          (N217)? commit_queue_q_5__address__28_ : 
                          (N219)? commit_queue_q_6__address__28_ : 
                          (N221)? commit_queue_q_7__address__28_ : 1'b0;
  assign req_port_o[93] = (N214)? commit_queue_q_0__address__27_ : 
                          (N216)? commit_queue_q_1__address__27_ : 
                          (N218)? commit_queue_q_2__address__27_ : 
                          (N220)? commit_queue_q_3__address__27_ : 
                          (N215)? commit_queue_q_4__address__27_ : 
                          (N217)? commit_queue_q_5__address__27_ : 
                          (N219)? commit_queue_q_6__address__27_ : 
                          (N221)? commit_queue_q_7__address__27_ : 1'b0;
  assign req_port_o[92] = (N214)? commit_queue_q_0__address__26_ : 
                          (N216)? commit_queue_q_1__address__26_ : 
                          (N218)? commit_queue_q_2__address__26_ : 
                          (N220)? commit_queue_q_3__address__26_ : 
                          (N215)? commit_queue_q_4__address__26_ : 
                          (N217)? commit_queue_q_5__address__26_ : 
                          (N219)? commit_queue_q_6__address__26_ : 
                          (N221)? commit_queue_q_7__address__26_ : 1'b0;
  assign req_port_o[91] = (N214)? commit_queue_q_0__address__25_ : 
                          (N216)? commit_queue_q_1__address__25_ : 
                          (N218)? commit_queue_q_2__address__25_ : 
                          (N220)? commit_queue_q_3__address__25_ : 
                          (N215)? commit_queue_q_4__address__25_ : 
                          (N217)? commit_queue_q_5__address__25_ : 
                          (N219)? commit_queue_q_6__address__25_ : 
                          (N221)? commit_queue_q_7__address__25_ : 1'b0;
  assign req_port_o[90] = (N214)? commit_queue_q_0__address__24_ : 
                          (N216)? commit_queue_q_1__address__24_ : 
                          (N218)? commit_queue_q_2__address__24_ : 
                          (N220)? commit_queue_q_3__address__24_ : 
                          (N215)? commit_queue_q_4__address__24_ : 
                          (N217)? commit_queue_q_5__address__24_ : 
                          (N219)? commit_queue_q_6__address__24_ : 
                          (N221)? commit_queue_q_7__address__24_ : 1'b0;
  assign req_port_o[89] = (N214)? commit_queue_q_0__address__23_ : 
                          (N216)? commit_queue_q_1__address__23_ : 
                          (N218)? commit_queue_q_2__address__23_ : 
                          (N220)? commit_queue_q_3__address__23_ : 
                          (N215)? commit_queue_q_4__address__23_ : 
                          (N217)? commit_queue_q_5__address__23_ : 
                          (N219)? commit_queue_q_6__address__23_ : 
                          (N221)? commit_queue_q_7__address__23_ : 1'b0;
  assign req_port_o[88] = (N214)? commit_queue_q_0__address__22_ : 
                          (N216)? commit_queue_q_1__address__22_ : 
                          (N218)? commit_queue_q_2__address__22_ : 
                          (N220)? commit_queue_q_3__address__22_ : 
                          (N215)? commit_queue_q_4__address__22_ : 
                          (N217)? commit_queue_q_5__address__22_ : 
                          (N219)? commit_queue_q_6__address__22_ : 
                          (N221)? commit_queue_q_7__address__22_ : 1'b0;
  assign req_port_o[87] = (N214)? commit_queue_q_0__address__21_ : 
                          (N216)? commit_queue_q_1__address__21_ : 
                          (N218)? commit_queue_q_2__address__21_ : 
                          (N220)? commit_queue_q_3__address__21_ : 
                          (N215)? commit_queue_q_4__address__21_ : 
                          (N217)? commit_queue_q_5__address__21_ : 
                          (N219)? commit_queue_q_6__address__21_ : 
                          (N221)? commit_queue_q_7__address__21_ : 1'b0;
  assign req_port_o[86] = (N214)? commit_queue_q_0__address__20_ : 
                          (N216)? commit_queue_q_1__address__20_ : 
                          (N218)? commit_queue_q_2__address__20_ : 
                          (N220)? commit_queue_q_3__address__20_ : 
                          (N215)? commit_queue_q_4__address__20_ : 
                          (N217)? commit_queue_q_5__address__20_ : 
                          (N219)? commit_queue_q_6__address__20_ : 
                          (N221)? commit_queue_q_7__address__20_ : 1'b0;
  assign req_port_o[85] = (N214)? commit_queue_q_0__address__19_ : 
                          (N216)? commit_queue_q_1__address__19_ : 
                          (N218)? commit_queue_q_2__address__19_ : 
                          (N220)? commit_queue_q_3__address__19_ : 
                          (N215)? commit_queue_q_4__address__19_ : 
                          (N217)? commit_queue_q_5__address__19_ : 
                          (N219)? commit_queue_q_6__address__19_ : 
                          (N221)? commit_queue_q_7__address__19_ : 1'b0;
  assign req_port_o[84] = (N214)? commit_queue_q_0__address__18_ : 
                          (N216)? commit_queue_q_1__address__18_ : 
                          (N218)? commit_queue_q_2__address__18_ : 
                          (N220)? commit_queue_q_3__address__18_ : 
                          (N215)? commit_queue_q_4__address__18_ : 
                          (N217)? commit_queue_q_5__address__18_ : 
                          (N219)? commit_queue_q_6__address__18_ : 
                          (N221)? commit_queue_q_7__address__18_ : 1'b0;
  assign req_port_o[83] = (N214)? commit_queue_q_0__address__17_ : 
                          (N216)? commit_queue_q_1__address__17_ : 
                          (N218)? commit_queue_q_2__address__17_ : 
                          (N220)? commit_queue_q_3__address__17_ : 
                          (N215)? commit_queue_q_4__address__17_ : 
                          (N217)? commit_queue_q_5__address__17_ : 
                          (N219)? commit_queue_q_6__address__17_ : 
                          (N221)? commit_queue_q_7__address__17_ : 1'b0;
  assign req_port_o[82] = (N214)? commit_queue_q_0__address__16_ : 
                          (N216)? commit_queue_q_1__address__16_ : 
                          (N218)? commit_queue_q_2__address__16_ : 
                          (N220)? commit_queue_q_3__address__16_ : 
                          (N215)? commit_queue_q_4__address__16_ : 
                          (N217)? commit_queue_q_5__address__16_ : 
                          (N219)? commit_queue_q_6__address__16_ : 
                          (N221)? commit_queue_q_7__address__16_ : 1'b0;
  assign req_port_o[81] = (N214)? commit_queue_q_0__address__15_ : 
                          (N216)? commit_queue_q_1__address__15_ : 
                          (N218)? commit_queue_q_2__address__15_ : 
                          (N220)? commit_queue_q_3__address__15_ : 
                          (N215)? commit_queue_q_4__address__15_ : 
                          (N217)? commit_queue_q_5__address__15_ : 
                          (N219)? commit_queue_q_6__address__15_ : 
                          (N221)? commit_queue_q_7__address__15_ : 1'b0;
  assign req_port_o[80] = (N214)? commit_queue_q_0__address__14_ : 
                          (N216)? commit_queue_q_1__address__14_ : 
                          (N218)? commit_queue_q_2__address__14_ : 
                          (N220)? commit_queue_q_3__address__14_ : 
                          (N215)? commit_queue_q_4__address__14_ : 
                          (N217)? commit_queue_q_5__address__14_ : 
                          (N219)? commit_queue_q_6__address__14_ : 
                          (N221)? commit_queue_q_7__address__14_ : 1'b0;
  assign req_port_o[79] = (N214)? commit_queue_q_0__address__13_ : 
                          (N216)? commit_queue_q_1__address__13_ : 
                          (N218)? commit_queue_q_2__address__13_ : 
                          (N220)? commit_queue_q_3__address__13_ : 
                          (N215)? commit_queue_q_4__address__13_ : 
                          (N217)? commit_queue_q_5__address__13_ : 
                          (N219)? commit_queue_q_6__address__13_ : 
                          (N221)? commit_queue_q_7__address__13_ : 1'b0;
  assign req_port_o[78] = (N214)? commit_queue_q_0__address__12_ : 
                          (N216)? commit_queue_q_1__address__12_ : 
                          (N218)? commit_queue_q_2__address__12_ : 
                          (N220)? commit_queue_q_3__address__12_ : 
                          (N215)? commit_queue_q_4__address__12_ : 
                          (N217)? commit_queue_q_5__address__12_ : 
                          (N219)? commit_queue_q_6__address__12_ : 
                          (N221)? commit_queue_q_7__address__12_ : 1'b0;
  assign req_port_o[77] = (N226)? commit_queue_q_0__data__63_ : 
                          (N228)? commit_queue_q_1__data__63_ : 
                          (N230)? commit_queue_q_2__data__63_ : 
                          (N232)? commit_queue_q_3__data__63_ : 
                          (N227)? commit_queue_q_4__data__63_ : 
                          (N229)? commit_queue_q_5__data__63_ : 
                          (N231)? commit_queue_q_6__data__63_ : 
                          (N233)? commit_queue_q_7__data__63_ : 1'b0;
  assign req_port_o[76] = (N226)? commit_queue_q_0__data__62_ : 
                          (N228)? commit_queue_q_1__data__62_ : 
                          (N230)? commit_queue_q_2__data__62_ : 
                          (N232)? commit_queue_q_3__data__62_ : 
                          (N227)? commit_queue_q_4__data__62_ : 
                          (N229)? commit_queue_q_5__data__62_ : 
                          (N231)? commit_queue_q_6__data__62_ : 
                          (N233)? commit_queue_q_7__data__62_ : 1'b0;
  assign req_port_o[75] = (N226)? commit_queue_q_0__data__61_ : 
                          (N228)? commit_queue_q_1__data__61_ : 
                          (N230)? commit_queue_q_2__data__61_ : 
                          (N232)? commit_queue_q_3__data__61_ : 
                          (N227)? commit_queue_q_4__data__61_ : 
                          (N229)? commit_queue_q_5__data__61_ : 
                          (N231)? commit_queue_q_6__data__61_ : 
                          (N233)? commit_queue_q_7__data__61_ : 1'b0;
  assign req_port_o[74] = (N226)? commit_queue_q_0__data__60_ : 
                          (N228)? commit_queue_q_1__data__60_ : 
                          (N230)? commit_queue_q_2__data__60_ : 
                          (N232)? commit_queue_q_3__data__60_ : 
                          (N227)? commit_queue_q_4__data__60_ : 
                          (N229)? commit_queue_q_5__data__60_ : 
                          (N231)? commit_queue_q_6__data__60_ : 
                          (N233)? commit_queue_q_7__data__60_ : 1'b0;
  assign req_port_o[73] = (N226)? commit_queue_q_0__data__59_ : 
                          (N228)? commit_queue_q_1__data__59_ : 
                          (N230)? commit_queue_q_2__data__59_ : 
                          (N232)? commit_queue_q_3__data__59_ : 
                          (N227)? commit_queue_q_4__data__59_ : 
                          (N229)? commit_queue_q_5__data__59_ : 
                          (N231)? commit_queue_q_6__data__59_ : 
                          (N233)? commit_queue_q_7__data__59_ : 1'b0;
  assign req_port_o[72] = (N226)? commit_queue_q_0__data__58_ : 
                          (N228)? commit_queue_q_1__data__58_ : 
                          (N230)? commit_queue_q_2__data__58_ : 
                          (N232)? commit_queue_q_3__data__58_ : 
                          (N227)? commit_queue_q_4__data__58_ : 
                          (N229)? commit_queue_q_5__data__58_ : 
                          (N231)? commit_queue_q_6__data__58_ : 
                          (N233)? commit_queue_q_7__data__58_ : 1'b0;
  assign req_port_o[71] = (N226)? commit_queue_q_0__data__57_ : 
                          (N228)? commit_queue_q_1__data__57_ : 
                          (N230)? commit_queue_q_2__data__57_ : 
                          (N232)? commit_queue_q_3__data__57_ : 
                          (N227)? commit_queue_q_4__data__57_ : 
                          (N229)? commit_queue_q_5__data__57_ : 
                          (N231)? commit_queue_q_6__data__57_ : 
                          (N233)? commit_queue_q_7__data__57_ : 1'b0;
  assign req_port_o[70] = (N226)? commit_queue_q_0__data__56_ : 
                          (N228)? commit_queue_q_1__data__56_ : 
                          (N230)? commit_queue_q_2__data__56_ : 
                          (N232)? commit_queue_q_3__data__56_ : 
                          (N227)? commit_queue_q_4__data__56_ : 
                          (N229)? commit_queue_q_5__data__56_ : 
                          (N231)? commit_queue_q_6__data__56_ : 
                          (N233)? commit_queue_q_7__data__56_ : 1'b0;
  assign req_port_o[69] = (N226)? commit_queue_q_0__data__55_ : 
                          (N228)? commit_queue_q_1__data__55_ : 
                          (N230)? commit_queue_q_2__data__55_ : 
                          (N232)? commit_queue_q_3__data__55_ : 
                          (N227)? commit_queue_q_4__data__55_ : 
                          (N229)? commit_queue_q_5__data__55_ : 
                          (N231)? commit_queue_q_6__data__55_ : 
                          (N233)? commit_queue_q_7__data__55_ : 1'b0;
  assign req_port_o[68] = (N226)? commit_queue_q_0__data__54_ : 
                          (N228)? commit_queue_q_1__data__54_ : 
                          (N230)? commit_queue_q_2__data__54_ : 
                          (N232)? commit_queue_q_3__data__54_ : 
                          (N227)? commit_queue_q_4__data__54_ : 
                          (N229)? commit_queue_q_5__data__54_ : 
                          (N231)? commit_queue_q_6__data__54_ : 
                          (N233)? commit_queue_q_7__data__54_ : 1'b0;
  assign req_port_o[67] = (N226)? commit_queue_q_0__data__53_ : 
                          (N228)? commit_queue_q_1__data__53_ : 
                          (N230)? commit_queue_q_2__data__53_ : 
                          (N232)? commit_queue_q_3__data__53_ : 
                          (N227)? commit_queue_q_4__data__53_ : 
                          (N229)? commit_queue_q_5__data__53_ : 
                          (N231)? commit_queue_q_6__data__53_ : 
                          (N233)? commit_queue_q_7__data__53_ : 1'b0;
  assign req_port_o[66] = (N226)? commit_queue_q_0__data__52_ : 
                          (N228)? commit_queue_q_1__data__52_ : 
                          (N230)? commit_queue_q_2__data__52_ : 
                          (N232)? commit_queue_q_3__data__52_ : 
                          (N227)? commit_queue_q_4__data__52_ : 
                          (N229)? commit_queue_q_5__data__52_ : 
                          (N231)? commit_queue_q_6__data__52_ : 
                          (N233)? commit_queue_q_7__data__52_ : 1'b0;
  assign req_port_o[65] = (N226)? commit_queue_q_0__data__51_ : 
                          (N228)? commit_queue_q_1__data__51_ : 
                          (N230)? commit_queue_q_2__data__51_ : 
                          (N232)? commit_queue_q_3__data__51_ : 
                          (N227)? commit_queue_q_4__data__51_ : 
                          (N229)? commit_queue_q_5__data__51_ : 
                          (N231)? commit_queue_q_6__data__51_ : 
                          (N233)? commit_queue_q_7__data__51_ : 1'b0;
  assign req_port_o[64] = (N226)? commit_queue_q_0__data__50_ : 
                          (N228)? commit_queue_q_1__data__50_ : 
                          (N230)? commit_queue_q_2__data__50_ : 
                          (N232)? commit_queue_q_3__data__50_ : 
                          (N227)? commit_queue_q_4__data__50_ : 
                          (N229)? commit_queue_q_5__data__50_ : 
                          (N231)? commit_queue_q_6__data__50_ : 
                          (N233)? commit_queue_q_7__data__50_ : 1'b0;
  assign req_port_o[63] = (N226)? commit_queue_q_0__data__49_ : 
                          (N228)? commit_queue_q_1__data__49_ : 
                          (N230)? commit_queue_q_2__data__49_ : 
                          (N232)? commit_queue_q_3__data__49_ : 
                          (N227)? commit_queue_q_4__data__49_ : 
                          (N229)? commit_queue_q_5__data__49_ : 
                          (N231)? commit_queue_q_6__data__49_ : 
                          (N233)? commit_queue_q_7__data__49_ : 1'b0;
  assign req_port_o[62] = (N226)? commit_queue_q_0__data__48_ : 
                          (N228)? commit_queue_q_1__data__48_ : 
                          (N230)? commit_queue_q_2__data__48_ : 
                          (N232)? commit_queue_q_3__data__48_ : 
                          (N227)? commit_queue_q_4__data__48_ : 
                          (N229)? commit_queue_q_5__data__48_ : 
                          (N231)? commit_queue_q_6__data__48_ : 
                          (N233)? commit_queue_q_7__data__48_ : 1'b0;
  assign req_port_o[61] = (N226)? commit_queue_q_0__data__47_ : 
                          (N228)? commit_queue_q_1__data__47_ : 
                          (N230)? commit_queue_q_2__data__47_ : 
                          (N232)? commit_queue_q_3__data__47_ : 
                          (N227)? commit_queue_q_4__data__47_ : 
                          (N229)? commit_queue_q_5__data__47_ : 
                          (N231)? commit_queue_q_6__data__47_ : 
                          (N233)? commit_queue_q_7__data__47_ : 1'b0;
  assign req_port_o[60] = (N226)? commit_queue_q_0__data__46_ : 
                          (N228)? commit_queue_q_1__data__46_ : 
                          (N230)? commit_queue_q_2__data__46_ : 
                          (N232)? commit_queue_q_3__data__46_ : 
                          (N227)? commit_queue_q_4__data__46_ : 
                          (N229)? commit_queue_q_5__data__46_ : 
                          (N231)? commit_queue_q_6__data__46_ : 
                          (N233)? commit_queue_q_7__data__46_ : 1'b0;
  assign req_port_o[59] = (N226)? commit_queue_q_0__data__45_ : 
                          (N228)? commit_queue_q_1__data__45_ : 
                          (N230)? commit_queue_q_2__data__45_ : 
                          (N232)? commit_queue_q_3__data__45_ : 
                          (N227)? commit_queue_q_4__data__45_ : 
                          (N229)? commit_queue_q_5__data__45_ : 
                          (N231)? commit_queue_q_6__data__45_ : 
                          (N233)? commit_queue_q_7__data__45_ : 1'b0;
  assign req_port_o[58] = (N226)? commit_queue_q_0__data__44_ : 
                          (N228)? commit_queue_q_1__data__44_ : 
                          (N230)? commit_queue_q_2__data__44_ : 
                          (N232)? commit_queue_q_3__data__44_ : 
                          (N227)? commit_queue_q_4__data__44_ : 
                          (N229)? commit_queue_q_5__data__44_ : 
                          (N231)? commit_queue_q_6__data__44_ : 
                          (N233)? commit_queue_q_7__data__44_ : 1'b0;
  assign req_port_o[57] = (N226)? commit_queue_q_0__data__43_ : 
                          (N228)? commit_queue_q_1__data__43_ : 
                          (N230)? commit_queue_q_2__data__43_ : 
                          (N232)? commit_queue_q_3__data__43_ : 
                          (N227)? commit_queue_q_4__data__43_ : 
                          (N229)? commit_queue_q_5__data__43_ : 
                          (N231)? commit_queue_q_6__data__43_ : 
                          (N233)? commit_queue_q_7__data__43_ : 1'b0;
  assign req_port_o[56] = (N226)? commit_queue_q_0__data__42_ : 
                          (N228)? commit_queue_q_1__data__42_ : 
                          (N230)? commit_queue_q_2__data__42_ : 
                          (N232)? commit_queue_q_3__data__42_ : 
                          (N227)? commit_queue_q_4__data__42_ : 
                          (N229)? commit_queue_q_5__data__42_ : 
                          (N231)? commit_queue_q_6__data__42_ : 
                          (N233)? commit_queue_q_7__data__42_ : 1'b0;
  assign req_port_o[55] = (N226)? commit_queue_q_0__data__41_ : 
                          (N228)? commit_queue_q_1__data__41_ : 
                          (N230)? commit_queue_q_2__data__41_ : 
                          (N232)? commit_queue_q_3__data__41_ : 
                          (N227)? commit_queue_q_4__data__41_ : 
                          (N229)? commit_queue_q_5__data__41_ : 
                          (N231)? commit_queue_q_6__data__41_ : 
                          (N233)? commit_queue_q_7__data__41_ : 1'b0;
  assign req_port_o[54] = (N226)? commit_queue_q_0__data__40_ : 
                          (N228)? commit_queue_q_1__data__40_ : 
                          (N230)? commit_queue_q_2__data__40_ : 
                          (N232)? commit_queue_q_3__data__40_ : 
                          (N227)? commit_queue_q_4__data__40_ : 
                          (N229)? commit_queue_q_5__data__40_ : 
                          (N231)? commit_queue_q_6__data__40_ : 
                          (N233)? commit_queue_q_7__data__40_ : 1'b0;
  assign req_port_o[53] = (N226)? commit_queue_q_0__data__39_ : 
                          (N228)? commit_queue_q_1__data__39_ : 
                          (N230)? commit_queue_q_2__data__39_ : 
                          (N232)? commit_queue_q_3__data__39_ : 
                          (N227)? commit_queue_q_4__data__39_ : 
                          (N229)? commit_queue_q_5__data__39_ : 
                          (N231)? commit_queue_q_6__data__39_ : 
                          (N233)? commit_queue_q_7__data__39_ : 1'b0;
  assign req_port_o[52] = (N226)? commit_queue_q_0__data__38_ : 
                          (N228)? commit_queue_q_1__data__38_ : 
                          (N230)? commit_queue_q_2__data__38_ : 
                          (N232)? commit_queue_q_3__data__38_ : 
                          (N227)? commit_queue_q_4__data__38_ : 
                          (N229)? commit_queue_q_5__data__38_ : 
                          (N231)? commit_queue_q_6__data__38_ : 
                          (N233)? commit_queue_q_7__data__38_ : 1'b0;
  assign req_port_o[51] = (N226)? commit_queue_q_0__data__37_ : 
                          (N228)? commit_queue_q_1__data__37_ : 
                          (N230)? commit_queue_q_2__data__37_ : 
                          (N232)? commit_queue_q_3__data__37_ : 
                          (N227)? commit_queue_q_4__data__37_ : 
                          (N229)? commit_queue_q_5__data__37_ : 
                          (N231)? commit_queue_q_6__data__37_ : 
                          (N233)? commit_queue_q_7__data__37_ : 1'b0;
  assign req_port_o[50] = (N226)? commit_queue_q_0__data__36_ : 
                          (N228)? commit_queue_q_1__data__36_ : 
                          (N230)? commit_queue_q_2__data__36_ : 
                          (N232)? commit_queue_q_3__data__36_ : 
                          (N227)? commit_queue_q_4__data__36_ : 
                          (N229)? commit_queue_q_5__data__36_ : 
                          (N231)? commit_queue_q_6__data__36_ : 
                          (N233)? commit_queue_q_7__data__36_ : 1'b0;
  assign req_port_o[49] = (N226)? commit_queue_q_0__data__35_ : 
                          (N228)? commit_queue_q_1__data__35_ : 
                          (N230)? commit_queue_q_2__data__35_ : 
                          (N232)? commit_queue_q_3__data__35_ : 
                          (N227)? commit_queue_q_4__data__35_ : 
                          (N229)? commit_queue_q_5__data__35_ : 
                          (N231)? commit_queue_q_6__data__35_ : 
                          (N233)? commit_queue_q_7__data__35_ : 1'b0;
  assign req_port_o[48] = (N226)? commit_queue_q_0__data__34_ : 
                          (N228)? commit_queue_q_1__data__34_ : 
                          (N230)? commit_queue_q_2__data__34_ : 
                          (N232)? commit_queue_q_3__data__34_ : 
                          (N227)? commit_queue_q_4__data__34_ : 
                          (N229)? commit_queue_q_5__data__34_ : 
                          (N231)? commit_queue_q_6__data__34_ : 
                          (N233)? commit_queue_q_7__data__34_ : 1'b0;
  assign req_port_o[47] = (N226)? commit_queue_q_0__data__33_ : 
                          (N228)? commit_queue_q_1__data__33_ : 
                          (N230)? commit_queue_q_2__data__33_ : 
                          (N232)? commit_queue_q_3__data__33_ : 
                          (N227)? commit_queue_q_4__data__33_ : 
                          (N229)? commit_queue_q_5__data__33_ : 
                          (N231)? commit_queue_q_6__data__33_ : 
                          (N233)? commit_queue_q_7__data__33_ : 1'b0;
  assign req_port_o[46] = (N226)? commit_queue_q_0__data__32_ : 
                          (N228)? commit_queue_q_1__data__32_ : 
                          (N230)? commit_queue_q_2__data__32_ : 
                          (N232)? commit_queue_q_3__data__32_ : 
                          (N227)? commit_queue_q_4__data__32_ : 
                          (N229)? commit_queue_q_5__data__32_ : 
                          (N231)? commit_queue_q_6__data__32_ : 
                          (N233)? commit_queue_q_7__data__32_ : 1'b0;
  assign req_port_o[45] = (N226)? commit_queue_q_0__data__31_ : 
                          (N228)? commit_queue_q_1__data__31_ : 
                          (N230)? commit_queue_q_2__data__31_ : 
                          (N232)? commit_queue_q_3__data__31_ : 
                          (N227)? commit_queue_q_4__data__31_ : 
                          (N229)? commit_queue_q_5__data__31_ : 
                          (N231)? commit_queue_q_6__data__31_ : 
                          (N233)? commit_queue_q_7__data__31_ : 1'b0;
  assign req_port_o[44] = (N226)? commit_queue_q_0__data__30_ : 
                          (N228)? commit_queue_q_1__data__30_ : 
                          (N230)? commit_queue_q_2__data__30_ : 
                          (N232)? commit_queue_q_3__data__30_ : 
                          (N227)? commit_queue_q_4__data__30_ : 
                          (N229)? commit_queue_q_5__data__30_ : 
                          (N231)? commit_queue_q_6__data__30_ : 
                          (N233)? commit_queue_q_7__data__30_ : 1'b0;
  assign req_port_o[43] = (N226)? commit_queue_q_0__data__29_ : 
                          (N228)? commit_queue_q_1__data__29_ : 
                          (N230)? commit_queue_q_2__data__29_ : 
                          (N232)? commit_queue_q_3__data__29_ : 
                          (N227)? commit_queue_q_4__data__29_ : 
                          (N229)? commit_queue_q_5__data__29_ : 
                          (N231)? commit_queue_q_6__data__29_ : 
                          (N233)? commit_queue_q_7__data__29_ : 1'b0;
  assign req_port_o[42] = (N226)? commit_queue_q_0__data__28_ : 
                          (N228)? commit_queue_q_1__data__28_ : 
                          (N230)? commit_queue_q_2__data__28_ : 
                          (N232)? commit_queue_q_3__data__28_ : 
                          (N227)? commit_queue_q_4__data__28_ : 
                          (N229)? commit_queue_q_5__data__28_ : 
                          (N231)? commit_queue_q_6__data__28_ : 
                          (N233)? commit_queue_q_7__data__28_ : 1'b0;
  assign req_port_o[41] = (N226)? commit_queue_q_0__data__27_ : 
                          (N228)? commit_queue_q_1__data__27_ : 
                          (N230)? commit_queue_q_2__data__27_ : 
                          (N232)? commit_queue_q_3__data__27_ : 
                          (N227)? commit_queue_q_4__data__27_ : 
                          (N229)? commit_queue_q_5__data__27_ : 
                          (N231)? commit_queue_q_6__data__27_ : 
                          (N233)? commit_queue_q_7__data__27_ : 1'b0;
  assign req_port_o[40] = (N226)? commit_queue_q_0__data__26_ : 
                          (N228)? commit_queue_q_1__data__26_ : 
                          (N230)? commit_queue_q_2__data__26_ : 
                          (N232)? commit_queue_q_3__data__26_ : 
                          (N227)? commit_queue_q_4__data__26_ : 
                          (N229)? commit_queue_q_5__data__26_ : 
                          (N231)? commit_queue_q_6__data__26_ : 
                          (N233)? commit_queue_q_7__data__26_ : 1'b0;
  assign req_port_o[39] = (N226)? commit_queue_q_0__data__25_ : 
                          (N228)? commit_queue_q_1__data__25_ : 
                          (N230)? commit_queue_q_2__data__25_ : 
                          (N232)? commit_queue_q_3__data__25_ : 
                          (N227)? commit_queue_q_4__data__25_ : 
                          (N229)? commit_queue_q_5__data__25_ : 
                          (N231)? commit_queue_q_6__data__25_ : 
                          (N233)? commit_queue_q_7__data__25_ : 1'b0;
  assign req_port_o[38] = (N226)? commit_queue_q_0__data__24_ : 
                          (N228)? commit_queue_q_1__data__24_ : 
                          (N230)? commit_queue_q_2__data__24_ : 
                          (N232)? commit_queue_q_3__data__24_ : 
                          (N227)? commit_queue_q_4__data__24_ : 
                          (N229)? commit_queue_q_5__data__24_ : 
                          (N231)? commit_queue_q_6__data__24_ : 
                          (N233)? commit_queue_q_7__data__24_ : 1'b0;
  assign req_port_o[37] = (N226)? commit_queue_q_0__data__23_ : 
                          (N228)? commit_queue_q_1__data__23_ : 
                          (N230)? commit_queue_q_2__data__23_ : 
                          (N232)? commit_queue_q_3__data__23_ : 
                          (N227)? commit_queue_q_4__data__23_ : 
                          (N229)? commit_queue_q_5__data__23_ : 
                          (N231)? commit_queue_q_6__data__23_ : 
                          (N233)? commit_queue_q_7__data__23_ : 1'b0;
  assign req_port_o[36] = (N226)? commit_queue_q_0__data__22_ : 
                          (N228)? commit_queue_q_1__data__22_ : 
                          (N230)? commit_queue_q_2__data__22_ : 
                          (N232)? commit_queue_q_3__data__22_ : 
                          (N227)? commit_queue_q_4__data__22_ : 
                          (N229)? commit_queue_q_5__data__22_ : 
                          (N231)? commit_queue_q_6__data__22_ : 
                          (N233)? commit_queue_q_7__data__22_ : 1'b0;
  assign req_port_o[35] = (N226)? commit_queue_q_0__data__21_ : 
                          (N228)? commit_queue_q_1__data__21_ : 
                          (N230)? commit_queue_q_2__data__21_ : 
                          (N232)? commit_queue_q_3__data__21_ : 
                          (N227)? commit_queue_q_4__data__21_ : 
                          (N229)? commit_queue_q_5__data__21_ : 
                          (N231)? commit_queue_q_6__data__21_ : 
                          (N233)? commit_queue_q_7__data__21_ : 1'b0;
  assign req_port_o[34] = (N226)? commit_queue_q_0__data__20_ : 
                          (N228)? commit_queue_q_1__data__20_ : 
                          (N230)? commit_queue_q_2__data__20_ : 
                          (N232)? commit_queue_q_3__data__20_ : 
                          (N227)? commit_queue_q_4__data__20_ : 
                          (N229)? commit_queue_q_5__data__20_ : 
                          (N231)? commit_queue_q_6__data__20_ : 
                          (N233)? commit_queue_q_7__data__20_ : 1'b0;
  assign req_port_o[33] = (N226)? commit_queue_q_0__data__19_ : 
                          (N228)? commit_queue_q_1__data__19_ : 
                          (N230)? commit_queue_q_2__data__19_ : 
                          (N232)? commit_queue_q_3__data__19_ : 
                          (N227)? commit_queue_q_4__data__19_ : 
                          (N229)? commit_queue_q_5__data__19_ : 
                          (N231)? commit_queue_q_6__data__19_ : 
                          (N233)? commit_queue_q_7__data__19_ : 1'b0;
  assign req_port_o[32] = (N226)? commit_queue_q_0__data__18_ : 
                          (N228)? commit_queue_q_1__data__18_ : 
                          (N230)? commit_queue_q_2__data__18_ : 
                          (N232)? commit_queue_q_3__data__18_ : 
                          (N227)? commit_queue_q_4__data__18_ : 
                          (N229)? commit_queue_q_5__data__18_ : 
                          (N231)? commit_queue_q_6__data__18_ : 
                          (N233)? commit_queue_q_7__data__18_ : 1'b0;
  assign req_port_o[31] = (N226)? commit_queue_q_0__data__17_ : 
                          (N228)? commit_queue_q_1__data__17_ : 
                          (N230)? commit_queue_q_2__data__17_ : 
                          (N232)? commit_queue_q_3__data__17_ : 
                          (N227)? commit_queue_q_4__data__17_ : 
                          (N229)? commit_queue_q_5__data__17_ : 
                          (N231)? commit_queue_q_6__data__17_ : 
                          (N233)? commit_queue_q_7__data__17_ : 1'b0;
  assign req_port_o[30] = (N226)? commit_queue_q_0__data__16_ : 
                          (N228)? commit_queue_q_1__data__16_ : 
                          (N230)? commit_queue_q_2__data__16_ : 
                          (N232)? commit_queue_q_3__data__16_ : 
                          (N227)? commit_queue_q_4__data__16_ : 
                          (N229)? commit_queue_q_5__data__16_ : 
                          (N231)? commit_queue_q_6__data__16_ : 
                          (N233)? commit_queue_q_7__data__16_ : 1'b0;
  assign req_port_o[29] = (N226)? commit_queue_q_0__data__15_ : 
                          (N228)? commit_queue_q_1__data__15_ : 
                          (N230)? commit_queue_q_2__data__15_ : 
                          (N232)? commit_queue_q_3__data__15_ : 
                          (N227)? commit_queue_q_4__data__15_ : 
                          (N229)? commit_queue_q_5__data__15_ : 
                          (N231)? commit_queue_q_6__data__15_ : 
                          (N233)? commit_queue_q_7__data__15_ : 1'b0;
  assign req_port_o[28] = (N226)? commit_queue_q_0__data__14_ : 
                          (N228)? commit_queue_q_1__data__14_ : 
                          (N230)? commit_queue_q_2__data__14_ : 
                          (N232)? commit_queue_q_3__data__14_ : 
                          (N227)? commit_queue_q_4__data__14_ : 
                          (N229)? commit_queue_q_5__data__14_ : 
                          (N231)? commit_queue_q_6__data__14_ : 
                          (N233)? commit_queue_q_7__data__14_ : 1'b0;
  assign req_port_o[27] = (N226)? commit_queue_q_0__data__13_ : 
                          (N228)? commit_queue_q_1__data__13_ : 
                          (N230)? commit_queue_q_2__data__13_ : 
                          (N232)? commit_queue_q_3__data__13_ : 
                          (N227)? commit_queue_q_4__data__13_ : 
                          (N229)? commit_queue_q_5__data__13_ : 
                          (N231)? commit_queue_q_6__data__13_ : 
                          (N233)? commit_queue_q_7__data__13_ : 1'b0;
  assign req_port_o[26] = (N226)? commit_queue_q_0__data__12_ : 
                          (N228)? commit_queue_q_1__data__12_ : 
                          (N230)? commit_queue_q_2__data__12_ : 
                          (N232)? commit_queue_q_3__data__12_ : 
                          (N227)? commit_queue_q_4__data__12_ : 
                          (N229)? commit_queue_q_5__data__12_ : 
                          (N231)? commit_queue_q_6__data__12_ : 
                          (N233)? commit_queue_q_7__data__12_ : 1'b0;
  assign req_port_o[25] = (N226)? commit_queue_q_0__data__11_ : 
                          (N228)? commit_queue_q_1__data__11_ : 
                          (N230)? commit_queue_q_2__data__11_ : 
                          (N232)? commit_queue_q_3__data__11_ : 
                          (N227)? commit_queue_q_4__data__11_ : 
                          (N229)? commit_queue_q_5__data__11_ : 
                          (N231)? commit_queue_q_6__data__11_ : 
                          (N233)? commit_queue_q_7__data__11_ : 1'b0;
  assign req_port_o[24] = (N226)? commit_queue_q_0__data__10_ : 
                          (N228)? commit_queue_q_1__data__10_ : 
                          (N230)? commit_queue_q_2__data__10_ : 
                          (N232)? commit_queue_q_3__data__10_ : 
                          (N227)? commit_queue_q_4__data__10_ : 
                          (N229)? commit_queue_q_5__data__10_ : 
                          (N231)? commit_queue_q_6__data__10_ : 
                          (N233)? commit_queue_q_7__data__10_ : 1'b0;
  assign req_port_o[23] = (N226)? commit_queue_q_0__data__9_ : 
                          (N228)? commit_queue_q_1__data__9_ : 
                          (N230)? commit_queue_q_2__data__9_ : 
                          (N232)? commit_queue_q_3__data__9_ : 
                          (N227)? commit_queue_q_4__data__9_ : 
                          (N229)? commit_queue_q_5__data__9_ : 
                          (N231)? commit_queue_q_6__data__9_ : 
                          (N233)? commit_queue_q_7__data__9_ : 1'b0;
  assign req_port_o[22] = (N226)? commit_queue_q_0__data__8_ : 
                          (N228)? commit_queue_q_1__data__8_ : 
                          (N230)? commit_queue_q_2__data__8_ : 
                          (N232)? commit_queue_q_3__data__8_ : 
                          (N227)? commit_queue_q_4__data__8_ : 
                          (N229)? commit_queue_q_5__data__8_ : 
                          (N231)? commit_queue_q_6__data__8_ : 
                          (N233)? commit_queue_q_7__data__8_ : 1'b0;
  assign req_port_o[21] = (N226)? commit_queue_q_0__data__7_ : 
                          (N228)? commit_queue_q_1__data__7_ : 
                          (N230)? commit_queue_q_2__data__7_ : 
                          (N232)? commit_queue_q_3__data__7_ : 
                          (N227)? commit_queue_q_4__data__7_ : 
                          (N229)? commit_queue_q_5__data__7_ : 
                          (N231)? commit_queue_q_6__data__7_ : 
                          (N233)? commit_queue_q_7__data__7_ : 1'b0;
  assign req_port_o[20] = (N226)? commit_queue_q_0__data__6_ : 
                          (N228)? commit_queue_q_1__data__6_ : 
                          (N230)? commit_queue_q_2__data__6_ : 
                          (N232)? commit_queue_q_3__data__6_ : 
                          (N227)? commit_queue_q_4__data__6_ : 
                          (N229)? commit_queue_q_5__data__6_ : 
                          (N231)? commit_queue_q_6__data__6_ : 
                          (N233)? commit_queue_q_7__data__6_ : 1'b0;
  assign req_port_o[19] = (N226)? commit_queue_q_0__data__5_ : 
                          (N228)? commit_queue_q_1__data__5_ : 
                          (N230)? commit_queue_q_2__data__5_ : 
                          (N232)? commit_queue_q_3__data__5_ : 
                          (N227)? commit_queue_q_4__data__5_ : 
                          (N229)? commit_queue_q_5__data__5_ : 
                          (N231)? commit_queue_q_6__data__5_ : 
                          (N233)? commit_queue_q_7__data__5_ : 1'b0;
  assign req_port_o[18] = (N226)? commit_queue_q_0__data__4_ : 
                          (N228)? commit_queue_q_1__data__4_ : 
                          (N230)? commit_queue_q_2__data__4_ : 
                          (N232)? commit_queue_q_3__data__4_ : 
                          (N227)? commit_queue_q_4__data__4_ : 
                          (N229)? commit_queue_q_5__data__4_ : 
                          (N231)? commit_queue_q_6__data__4_ : 
                          (N233)? commit_queue_q_7__data__4_ : 1'b0;
  assign req_port_o[17] = (N226)? commit_queue_q_0__data__3_ : 
                          (N228)? commit_queue_q_1__data__3_ : 
                          (N230)? commit_queue_q_2__data__3_ : 
                          (N232)? commit_queue_q_3__data__3_ : 
                          (N227)? commit_queue_q_4__data__3_ : 
                          (N229)? commit_queue_q_5__data__3_ : 
                          (N231)? commit_queue_q_6__data__3_ : 
                          (N233)? commit_queue_q_7__data__3_ : 1'b0;
  assign req_port_o[16] = (N226)? commit_queue_q_0__data__2_ : 
                          (N228)? commit_queue_q_1__data__2_ : 
                          (N230)? commit_queue_q_2__data__2_ : 
                          (N232)? commit_queue_q_3__data__2_ : 
                          (N227)? commit_queue_q_4__data__2_ : 
                          (N229)? commit_queue_q_5__data__2_ : 
                          (N231)? commit_queue_q_6__data__2_ : 
                          (N233)? commit_queue_q_7__data__2_ : 1'b0;
  assign req_port_o[15] = (N226)? commit_queue_q_0__data__1_ : 
                          (N228)? commit_queue_q_1__data__1_ : 
                          (N230)? commit_queue_q_2__data__1_ : 
                          (N232)? commit_queue_q_3__data__1_ : 
                          (N227)? commit_queue_q_4__data__1_ : 
                          (N229)? commit_queue_q_5__data__1_ : 
                          (N231)? commit_queue_q_6__data__1_ : 
                          (N233)? commit_queue_q_7__data__1_ : 1'b0;
  assign req_port_o[14] = (N226)? commit_queue_q_0__data__0_ : 
                          (N228)? commit_queue_q_1__data__0_ : 
                          (N230)? commit_queue_q_2__data__0_ : 
                          (N232)? commit_queue_q_3__data__0_ : 
                          (N227)? commit_queue_q_4__data__0_ : 
                          (N229)? commit_queue_q_5__data__0_ : 
                          (N231)? commit_queue_q_6__data__0_ : 
                          (N233)? commit_queue_q_7__data__0_ : 1'b0;
  assign req_port_o[11] = (N238)? commit_queue_q_0__be__7_ : 
                          (N240)? commit_queue_q_1__be__7_ : 
                          (N242)? commit_queue_q_2__be__7_ : 
                          (N244)? commit_queue_q_3__be__7_ : 
                          (N239)? commit_queue_q_4__be__7_ : 
                          (N241)? commit_queue_q_5__be__7_ : 
                          (N243)? commit_queue_q_6__be__7_ : 
                          (N245)? commit_queue_q_7__be__7_ : 1'b0;
  assign req_port_o[10] = (N238)? commit_queue_q_0__be__6_ : 
                          (N240)? commit_queue_q_1__be__6_ : 
                          (N242)? commit_queue_q_2__be__6_ : 
                          (N244)? commit_queue_q_3__be__6_ : 
                          (N239)? commit_queue_q_4__be__6_ : 
                          (N241)? commit_queue_q_5__be__6_ : 
                          (N243)? commit_queue_q_6__be__6_ : 
                          (N245)? commit_queue_q_7__be__6_ : 1'b0;
  assign req_port_o[9] = (N238)? commit_queue_q_0__be__5_ : 
                         (N240)? commit_queue_q_1__be__5_ : 
                         (N242)? commit_queue_q_2__be__5_ : 
                         (N244)? commit_queue_q_3__be__5_ : 
                         (N239)? commit_queue_q_4__be__5_ : 
                         (N241)? commit_queue_q_5__be__5_ : 
                         (N243)? commit_queue_q_6__be__5_ : 
                         (N245)? commit_queue_q_7__be__5_ : 1'b0;
  assign req_port_o[8] = (N238)? commit_queue_q_0__be__4_ : 
                         (N240)? commit_queue_q_1__be__4_ : 
                         (N242)? commit_queue_q_2__be__4_ : 
                         (N244)? commit_queue_q_3__be__4_ : 
                         (N239)? commit_queue_q_4__be__4_ : 
                         (N241)? commit_queue_q_5__be__4_ : 
                         (N243)? commit_queue_q_6__be__4_ : 
                         (N245)? commit_queue_q_7__be__4_ : 1'b0;
  assign req_port_o[7] = (N238)? commit_queue_q_0__be__3_ : 
                         (N240)? commit_queue_q_1__be__3_ : 
                         (N242)? commit_queue_q_2__be__3_ : 
                         (N244)? commit_queue_q_3__be__3_ : 
                         (N239)? commit_queue_q_4__be__3_ : 
                         (N241)? commit_queue_q_5__be__3_ : 
                         (N243)? commit_queue_q_6__be__3_ : 
                         (N245)? commit_queue_q_7__be__3_ : 1'b0;
  assign req_port_o[6] = (N238)? commit_queue_q_0__be__2_ : 
                         (N240)? commit_queue_q_1__be__2_ : 
                         (N242)? commit_queue_q_2__be__2_ : 
                         (N244)? commit_queue_q_3__be__2_ : 
                         (N239)? commit_queue_q_4__be__2_ : 
                         (N241)? commit_queue_q_5__be__2_ : 
                         (N243)? commit_queue_q_6__be__2_ : 
                         (N245)? commit_queue_q_7__be__2_ : 1'b0;
  assign req_port_o[5] = (N238)? commit_queue_q_0__be__1_ : 
                         (N240)? commit_queue_q_1__be__1_ : 
                         (N242)? commit_queue_q_2__be__1_ : 
                         (N244)? commit_queue_q_3__be__1_ : 
                         (N239)? commit_queue_q_4__be__1_ : 
                         (N241)? commit_queue_q_5__be__1_ : 
                         (N243)? commit_queue_q_6__be__1_ : 
                         (N245)? commit_queue_q_7__be__1_ : 1'b0;
  assign req_port_o[4] = (N238)? commit_queue_q_0__be__0_ : 
                         (N240)? commit_queue_q_1__be__0_ : 
                         (N242)? commit_queue_q_2__be__0_ : 
                         (N244)? commit_queue_q_3__be__0_ : 
                         (N239)? commit_queue_q_4__be__0_ : 
                         (N241)? commit_queue_q_5__be__0_ : 
                         (N243)? commit_queue_q_6__be__0_ : 
                         (N245)? commit_queue_q_7__be__0_ : 1'b0;
  assign req_port_o[3] = (N250)? commit_queue_q_0__data_size__1_ : 
                         (N252)? commit_queue_q_1__data_size__1_ : 
                         (N254)? commit_queue_q_2__data_size__1_ : 
                         (N256)? commit_queue_q_3__data_size__1_ : 
                         (N251)? commit_queue_q_4__data_size__1_ : 
                         (N253)? commit_queue_q_5__data_size__1_ : 
                         (N255)? commit_queue_q_6__data_size__1_ : 
                         (N257)? commit_queue_q_7__data_size__1_ : 1'b0;
  assign req_port_o[2] = (N250)? commit_queue_q_0__data_size__0_ : 
                         (N252)? commit_queue_q_1__data_size__0_ : 
                         (N254)? commit_queue_q_2__data_size__0_ : 
                         (N256)? commit_queue_q_3__data_size__0_ : 
                         (N251)? commit_queue_q_4__data_size__0_ : 
                         (N253)? commit_queue_q_5__data_size__0_ : 
                         (N255)? commit_queue_q_6__data_size__0_ : 
                         (N257)? commit_queue_q_7__data_size__0_ : 1'b0;
  assign N270 = (N262)? commit_queue_q_0__valid_ : 
                (N264)? commit_queue_q_1__valid_ : 
                (N266)? commit_queue_q_2__valid_ : 
                (N268)? commit_queue_q_3__valid_ : 
                (N263)? commit_queue_q_4__valid_ : 
                (N265)? commit_queue_q_5__valid_ : 
                (N267)? commit_queue_q_6__valid_ : 
                (N269)? commit_queue_q_7__valid_ : 1'b0;
  assign N328 = (N324)? speculative_queue_q_0__address__55_ : 
                (N326)? speculative_queue_q_1__address__55_ : 
                (N325)? speculative_queue_q_2__address__55_ : 
                (N327)? speculative_queue_q_3__address__55_ : 1'b0;
  assign N329 = (N324)? speculative_queue_q_0__address__54_ : 
                (N326)? speculative_queue_q_1__address__54_ : 
                (N325)? speculative_queue_q_2__address__54_ : 
                (N327)? speculative_queue_q_3__address__54_ : 1'b0;
  assign N330 = (N324)? speculative_queue_q_0__address__53_ : 
                (N326)? speculative_queue_q_1__address__53_ : 
                (N325)? speculative_queue_q_2__address__53_ : 
                (N327)? speculative_queue_q_3__address__53_ : 1'b0;
  assign N331 = (N324)? speculative_queue_q_0__address__52_ : 
                (N326)? speculative_queue_q_1__address__52_ : 
                (N325)? speculative_queue_q_2__address__52_ : 
                (N327)? speculative_queue_q_3__address__52_ : 1'b0;
  assign N332 = (N324)? speculative_queue_q_0__address__51_ : 
                (N326)? speculative_queue_q_1__address__51_ : 
                (N325)? speculative_queue_q_2__address__51_ : 
                (N327)? speculative_queue_q_3__address__51_ : 1'b0;
  assign N333 = (N324)? speculative_queue_q_0__address__50_ : 
                (N326)? speculative_queue_q_1__address__50_ : 
                (N325)? speculative_queue_q_2__address__50_ : 
                (N327)? speculative_queue_q_3__address__50_ : 1'b0;
  assign N334 = (N324)? speculative_queue_q_0__address__49_ : 
                (N326)? speculative_queue_q_1__address__49_ : 
                (N325)? speculative_queue_q_2__address__49_ : 
                (N327)? speculative_queue_q_3__address__49_ : 1'b0;
  assign N335 = (N324)? speculative_queue_q_0__address__48_ : 
                (N326)? speculative_queue_q_1__address__48_ : 
                (N325)? speculative_queue_q_2__address__48_ : 
                (N327)? speculative_queue_q_3__address__48_ : 1'b0;
  assign N336 = (N324)? speculative_queue_q_0__address__47_ : 
                (N326)? speculative_queue_q_1__address__47_ : 
                (N325)? speculative_queue_q_2__address__47_ : 
                (N327)? speculative_queue_q_3__address__47_ : 1'b0;
  assign N337 = (N324)? speculative_queue_q_0__address__46_ : 
                (N326)? speculative_queue_q_1__address__46_ : 
                (N325)? speculative_queue_q_2__address__46_ : 
                (N327)? speculative_queue_q_3__address__46_ : 1'b0;
  assign N338 = (N324)? speculative_queue_q_0__address__45_ : 
                (N326)? speculative_queue_q_1__address__45_ : 
                (N325)? speculative_queue_q_2__address__45_ : 
                (N327)? speculative_queue_q_3__address__45_ : 1'b0;
  assign N339 = (N324)? speculative_queue_q_0__address__44_ : 
                (N326)? speculative_queue_q_1__address__44_ : 
                (N325)? speculative_queue_q_2__address__44_ : 
                (N327)? speculative_queue_q_3__address__44_ : 1'b0;
  assign N340 = (N324)? speculative_queue_q_0__address__43_ : 
                (N326)? speculative_queue_q_1__address__43_ : 
                (N325)? speculative_queue_q_2__address__43_ : 
                (N327)? speculative_queue_q_3__address__43_ : 1'b0;
  assign N341 = (N324)? speculative_queue_q_0__address__42_ : 
                (N326)? speculative_queue_q_1__address__42_ : 
                (N325)? speculative_queue_q_2__address__42_ : 
                (N327)? speculative_queue_q_3__address__42_ : 1'b0;
  assign N342 = (N324)? speculative_queue_q_0__address__41_ : 
                (N326)? speculative_queue_q_1__address__41_ : 
                (N325)? speculative_queue_q_2__address__41_ : 
                (N327)? speculative_queue_q_3__address__41_ : 1'b0;
  assign N343 = (N324)? speculative_queue_q_0__address__40_ : 
                (N326)? speculative_queue_q_1__address__40_ : 
                (N325)? speculative_queue_q_2__address__40_ : 
                (N327)? speculative_queue_q_3__address__40_ : 1'b0;
  assign N344 = (N324)? speculative_queue_q_0__address__39_ : 
                (N326)? speculative_queue_q_1__address__39_ : 
                (N325)? speculative_queue_q_2__address__39_ : 
                (N327)? speculative_queue_q_3__address__39_ : 1'b0;
  assign N345 = (N324)? speculative_queue_q_0__address__38_ : 
                (N326)? speculative_queue_q_1__address__38_ : 
                (N325)? speculative_queue_q_2__address__38_ : 
                (N327)? speculative_queue_q_3__address__38_ : 1'b0;
  assign N346 = (N324)? speculative_queue_q_0__address__37_ : 
                (N326)? speculative_queue_q_1__address__37_ : 
                (N325)? speculative_queue_q_2__address__37_ : 
                (N327)? speculative_queue_q_3__address__37_ : 1'b0;
  assign N347 = (N324)? speculative_queue_q_0__address__36_ : 
                (N326)? speculative_queue_q_1__address__36_ : 
                (N325)? speculative_queue_q_2__address__36_ : 
                (N327)? speculative_queue_q_3__address__36_ : 1'b0;
  assign N348 = (N324)? speculative_queue_q_0__address__35_ : 
                (N326)? speculative_queue_q_1__address__35_ : 
                (N325)? speculative_queue_q_2__address__35_ : 
                (N327)? speculative_queue_q_3__address__35_ : 1'b0;
  assign N349 = (N324)? speculative_queue_q_0__address__34_ : 
                (N326)? speculative_queue_q_1__address__34_ : 
                (N325)? speculative_queue_q_2__address__34_ : 
                (N327)? speculative_queue_q_3__address__34_ : 1'b0;
  assign N350 = (N324)? speculative_queue_q_0__address__33_ : 
                (N326)? speculative_queue_q_1__address__33_ : 
                (N325)? speculative_queue_q_2__address__33_ : 
                (N327)? speculative_queue_q_3__address__33_ : 1'b0;
  assign N351 = (N324)? speculative_queue_q_0__address__32_ : 
                (N326)? speculative_queue_q_1__address__32_ : 
                (N325)? speculative_queue_q_2__address__32_ : 
                (N327)? speculative_queue_q_3__address__32_ : 1'b0;
  assign N352 = (N324)? speculative_queue_q_0__address__31_ : 
                (N326)? speculative_queue_q_1__address__31_ : 
                (N325)? speculative_queue_q_2__address__31_ : 
                (N327)? speculative_queue_q_3__address__31_ : 1'b0;
  assign N353 = (N324)? speculative_queue_q_0__address__30_ : 
                (N326)? speculative_queue_q_1__address__30_ : 
                (N325)? speculative_queue_q_2__address__30_ : 
                (N327)? speculative_queue_q_3__address__30_ : 1'b0;
  assign N354 = (N324)? speculative_queue_q_0__address__29_ : 
                (N326)? speculative_queue_q_1__address__29_ : 
                (N325)? speculative_queue_q_2__address__29_ : 
                (N327)? speculative_queue_q_3__address__29_ : 1'b0;
  assign N355 = (N324)? speculative_queue_q_0__address__28_ : 
                (N326)? speculative_queue_q_1__address__28_ : 
                (N325)? speculative_queue_q_2__address__28_ : 
                (N327)? speculative_queue_q_3__address__28_ : 1'b0;
  assign N356 = (N324)? speculative_queue_q_0__address__27_ : 
                (N326)? speculative_queue_q_1__address__27_ : 
                (N325)? speculative_queue_q_2__address__27_ : 
                (N327)? speculative_queue_q_3__address__27_ : 1'b0;
  assign N357 = (N324)? speculative_queue_q_0__address__26_ : 
                (N326)? speculative_queue_q_1__address__26_ : 
                (N325)? speculative_queue_q_2__address__26_ : 
                (N327)? speculative_queue_q_3__address__26_ : 1'b0;
  assign N358 = (N324)? speculative_queue_q_0__address__25_ : 
                (N326)? speculative_queue_q_1__address__25_ : 
                (N325)? speculative_queue_q_2__address__25_ : 
                (N327)? speculative_queue_q_3__address__25_ : 1'b0;
  assign N359 = (N324)? speculative_queue_q_0__address__24_ : 
                (N326)? speculative_queue_q_1__address__24_ : 
                (N325)? speculative_queue_q_2__address__24_ : 
                (N327)? speculative_queue_q_3__address__24_ : 1'b0;
  assign N360 = (N324)? speculative_queue_q_0__address__23_ : 
                (N326)? speculative_queue_q_1__address__23_ : 
                (N325)? speculative_queue_q_2__address__23_ : 
                (N327)? speculative_queue_q_3__address__23_ : 1'b0;
  assign N361 = (N324)? speculative_queue_q_0__address__22_ : 
                (N326)? speculative_queue_q_1__address__22_ : 
                (N325)? speculative_queue_q_2__address__22_ : 
                (N327)? speculative_queue_q_3__address__22_ : 1'b0;
  assign N362 = (N324)? speculative_queue_q_0__address__21_ : 
                (N326)? speculative_queue_q_1__address__21_ : 
                (N325)? speculative_queue_q_2__address__21_ : 
                (N327)? speculative_queue_q_3__address__21_ : 1'b0;
  assign N363 = (N324)? speculative_queue_q_0__address__20_ : 
                (N326)? speculative_queue_q_1__address__20_ : 
                (N325)? speculative_queue_q_2__address__20_ : 
                (N327)? speculative_queue_q_3__address__20_ : 1'b0;
  assign N364 = (N324)? speculative_queue_q_0__address__19_ : 
                (N326)? speculative_queue_q_1__address__19_ : 
                (N325)? speculative_queue_q_2__address__19_ : 
                (N327)? speculative_queue_q_3__address__19_ : 1'b0;
  assign N365 = (N324)? speculative_queue_q_0__address__18_ : 
                (N326)? speculative_queue_q_1__address__18_ : 
                (N325)? speculative_queue_q_2__address__18_ : 
                (N327)? speculative_queue_q_3__address__18_ : 1'b0;
  assign N366 = (N324)? speculative_queue_q_0__address__17_ : 
                (N326)? speculative_queue_q_1__address__17_ : 
                (N325)? speculative_queue_q_2__address__17_ : 
                (N327)? speculative_queue_q_3__address__17_ : 1'b0;
  assign N367 = (N324)? speculative_queue_q_0__address__16_ : 
                (N326)? speculative_queue_q_1__address__16_ : 
                (N325)? speculative_queue_q_2__address__16_ : 
                (N327)? speculative_queue_q_3__address__16_ : 1'b0;
  assign N368 = (N324)? speculative_queue_q_0__address__15_ : 
                (N326)? speculative_queue_q_1__address__15_ : 
                (N325)? speculative_queue_q_2__address__15_ : 
                (N327)? speculative_queue_q_3__address__15_ : 1'b0;
  assign N369 = (N324)? speculative_queue_q_0__address__14_ : 
                (N326)? speculative_queue_q_1__address__14_ : 
                (N325)? speculative_queue_q_2__address__14_ : 
                (N327)? speculative_queue_q_3__address__14_ : 1'b0;
  assign N370 = (N324)? speculative_queue_q_0__address__13_ : 
                (N326)? speculative_queue_q_1__address__13_ : 
                (N325)? speculative_queue_q_2__address__13_ : 
                (N327)? speculative_queue_q_3__address__13_ : 1'b0;
  assign N371 = (N324)? speculative_queue_q_0__address__12_ : 
                (N326)? speculative_queue_q_1__address__12_ : 
                (N325)? speculative_queue_q_2__address__12_ : 
                (N327)? speculative_queue_q_3__address__12_ : 1'b0;
  assign N372 = (N324)? speculative_queue_q_0__address__11_ : 
                (N326)? speculative_queue_q_1__address__11_ : 
                (N325)? speculative_queue_q_2__address__11_ : 
                (N327)? speculative_queue_q_3__address__11_ : 1'b0;
  assign N373 = (N324)? speculative_queue_q_0__address__10_ : 
                (N326)? speculative_queue_q_1__address__10_ : 
                (N325)? speculative_queue_q_2__address__10_ : 
                (N327)? speculative_queue_q_3__address__10_ : 1'b0;
  assign N374 = (N324)? speculative_queue_q_0__address__9_ : 
                (N326)? speculative_queue_q_1__address__9_ : 
                (N325)? speculative_queue_q_2__address__9_ : 
                (N327)? speculative_queue_q_3__address__9_ : 1'b0;
  assign N375 = (N324)? speculative_queue_q_0__address__8_ : 
                (N326)? speculative_queue_q_1__address__8_ : 
                (N325)? speculative_queue_q_2__address__8_ : 
                (N327)? speculative_queue_q_3__address__8_ : 1'b0;
  assign N376 = (N324)? speculative_queue_q_0__address__7_ : 
                (N326)? speculative_queue_q_1__address__7_ : 
                (N325)? speculative_queue_q_2__address__7_ : 
                (N327)? speculative_queue_q_3__address__7_ : 1'b0;
  assign N377 = (N324)? speculative_queue_q_0__address__6_ : 
                (N326)? speculative_queue_q_1__address__6_ : 
                (N325)? speculative_queue_q_2__address__6_ : 
                (N327)? speculative_queue_q_3__address__6_ : 1'b0;
  assign N378 = (N324)? speculative_queue_q_0__address__5_ : 
                (N326)? speculative_queue_q_1__address__5_ : 
                (N325)? speculative_queue_q_2__address__5_ : 
                (N327)? speculative_queue_q_3__address__5_ : 1'b0;
  assign N379 = (N324)? speculative_queue_q_0__address__4_ : 
                (N326)? speculative_queue_q_1__address__4_ : 
                (N325)? speculative_queue_q_2__address__4_ : 
                (N327)? speculative_queue_q_3__address__4_ : 1'b0;
  assign N380 = (N324)? speculative_queue_q_0__address__3_ : 
                (N326)? speculative_queue_q_1__address__3_ : 
                (N325)? speculative_queue_q_2__address__3_ : 
                (N327)? speculative_queue_q_3__address__3_ : 1'b0;
  assign N381 = (N324)? speculative_queue_q_0__address__2_ : 
                (N326)? speculative_queue_q_1__address__2_ : 
                (N325)? speculative_queue_q_2__address__2_ : 
                (N327)? speculative_queue_q_3__address__2_ : 1'b0;
  assign N382 = (N324)? speculative_queue_q_0__address__1_ : 
                (N326)? speculative_queue_q_1__address__1_ : 
                (N325)? speculative_queue_q_2__address__1_ : 
                (N327)? speculative_queue_q_3__address__1_ : 1'b0;
  assign N383 = (N324)? speculative_queue_q_0__address__0_ : 
                (N326)? speculative_queue_q_1__address__0_ : 
                (N325)? speculative_queue_q_2__address__0_ : 
                (N327)? speculative_queue_q_3__address__0_ : 1'b0;
  assign N384 = (N324)? speculative_queue_q_0__data__63_ : 
                (N326)? speculative_queue_q_1__data__63_ : 
                (N325)? speculative_queue_q_2__data__63_ : 
                (N327)? speculative_queue_q_3__data__63_ : 1'b0;
  assign N385 = (N324)? speculative_queue_q_0__data__62_ : 
                (N326)? speculative_queue_q_1__data__62_ : 
                (N325)? speculative_queue_q_2__data__62_ : 
                (N327)? speculative_queue_q_3__data__62_ : 1'b0;
  assign N386 = (N324)? speculative_queue_q_0__data__61_ : 
                (N326)? speculative_queue_q_1__data__61_ : 
                (N325)? speculative_queue_q_2__data__61_ : 
                (N327)? speculative_queue_q_3__data__61_ : 1'b0;
  assign N387 = (N324)? speculative_queue_q_0__data__60_ : 
                (N326)? speculative_queue_q_1__data__60_ : 
                (N325)? speculative_queue_q_2__data__60_ : 
                (N327)? speculative_queue_q_3__data__60_ : 1'b0;
  assign N388 = (N324)? speculative_queue_q_0__data__59_ : 
                (N326)? speculative_queue_q_1__data__59_ : 
                (N325)? speculative_queue_q_2__data__59_ : 
                (N327)? speculative_queue_q_3__data__59_ : 1'b0;
  assign N389 = (N324)? speculative_queue_q_0__data__58_ : 
                (N326)? speculative_queue_q_1__data__58_ : 
                (N325)? speculative_queue_q_2__data__58_ : 
                (N327)? speculative_queue_q_3__data__58_ : 1'b0;
  assign N390 = (N324)? speculative_queue_q_0__data__57_ : 
                (N326)? speculative_queue_q_1__data__57_ : 
                (N325)? speculative_queue_q_2__data__57_ : 
                (N327)? speculative_queue_q_3__data__57_ : 1'b0;
  assign N391 = (N324)? speculative_queue_q_0__data__56_ : 
                (N326)? speculative_queue_q_1__data__56_ : 
                (N325)? speculative_queue_q_2__data__56_ : 
                (N327)? speculative_queue_q_3__data__56_ : 1'b0;
  assign N392 = (N324)? speculative_queue_q_0__data__55_ : 
                (N326)? speculative_queue_q_1__data__55_ : 
                (N325)? speculative_queue_q_2__data__55_ : 
                (N327)? speculative_queue_q_3__data__55_ : 1'b0;
  assign N393 = (N324)? speculative_queue_q_0__data__54_ : 
                (N326)? speculative_queue_q_1__data__54_ : 
                (N325)? speculative_queue_q_2__data__54_ : 
                (N327)? speculative_queue_q_3__data__54_ : 1'b0;
  assign N394 = (N324)? speculative_queue_q_0__data__53_ : 
                (N326)? speculative_queue_q_1__data__53_ : 
                (N325)? speculative_queue_q_2__data__53_ : 
                (N327)? speculative_queue_q_3__data__53_ : 1'b0;
  assign N395 = (N324)? speculative_queue_q_0__data__52_ : 
                (N326)? speculative_queue_q_1__data__52_ : 
                (N325)? speculative_queue_q_2__data__52_ : 
                (N327)? speculative_queue_q_3__data__52_ : 1'b0;
  assign N396 = (N324)? speculative_queue_q_0__data__51_ : 
                (N326)? speculative_queue_q_1__data__51_ : 
                (N325)? speculative_queue_q_2__data__51_ : 
                (N327)? speculative_queue_q_3__data__51_ : 1'b0;
  assign N397 = (N324)? speculative_queue_q_0__data__50_ : 
                (N326)? speculative_queue_q_1__data__50_ : 
                (N325)? speculative_queue_q_2__data__50_ : 
                (N327)? speculative_queue_q_3__data__50_ : 1'b0;
  assign N398 = (N324)? speculative_queue_q_0__data__49_ : 
                (N326)? speculative_queue_q_1__data__49_ : 
                (N325)? speculative_queue_q_2__data__49_ : 
                (N327)? speculative_queue_q_3__data__49_ : 1'b0;
  assign N399 = (N324)? speculative_queue_q_0__data__48_ : 
                (N326)? speculative_queue_q_1__data__48_ : 
                (N325)? speculative_queue_q_2__data__48_ : 
                (N327)? speculative_queue_q_3__data__48_ : 1'b0;
  assign N400 = (N324)? speculative_queue_q_0__data__47_ : 
                (N326)? speculative_queue_q_1__data__47_ : 
                (N325)? speculative_queue_q_2__data__47_ : 
                (N327)? speculative_queue_q_3__data__47_ : 1'b0;
  assign N401 = (N324)? speculative_queue_q_0__data__46_ : 
                (N326)? speculative_queue_q_1__data__46_ : 
                (N325)? speculative_queue_q_2__data__46_ : 
                (N327)? speculative_queue_q_3__data__46_ : 1'b0;
  assign N402 = (N324)? speculative_queue_q_0__data__45_ : 
                (N326)? speculative_queue_q_1__data__45_ : 
                (N325)? speculative_queue_q_2__data__45_ : 
                (N327)? speculative_queue_q_3__data__45_ : 1'b0;
  assign N403 = (N324)? speculative_queue_q_0__data__44_ : 
                (N326)? speculative_queue_q_1__data__44_ : 
                (N325)? speculative_queue_q_2__data__44_ : 
                (N327)? speculative_queue_q_3__data__44_ : 1'b0;
  assign N404 = (N324)? speculative_queue_q_0__data__43_ : 
                (N326)? speculative_queue_q_1__data__43_ : 
                (N325)? speculative_queue_q_2__data__43_ : 
                (N327)? speculative_queue_q_3__data__43_ : 1'b0;
  assign N405 = (N324)? speculative_queue_q_0__data__42_ : 
                (N326)? speculative_queue_q_1__data__42_ : 
                (N325)? speculative_queue_q_2__data__42_ : 
                (N327)? speculative_queue_q_3__data__42_ : 1'b0;
  assign N406 = (N324)? speculative_queue_q_0__data__41_ : 
                (N326)? speculative_queue_q_1__data__41_ : 
                (N325)? speculative_queue_q_2__data__41_ : 
                (N327)? speculative_queue_q_3__data__41_ : 1'b0;
  assign N407 = (N324)? speculative_queue_q_0__data__40_ : 
                (N326)? speculative_queue_q_1__data__40_ : 
                (N325)? speculative_queue_q_2__data__40_ : 
                (N327)? speculative_queue_q_3__data__40_ : 1'b0;
  assign N408 = (N324)? speculative_queue_q_0__data__39_ : 
                (N326)? speculative_queue_q_1__data__39_ : 
                (N325)? speculative_queue_q_2__data__39_ : 
                (N327)? speculative_queue_q_3__data__39_ : 1'b0;
  assign N409 = (N324)? speculative_queue_q_0__data__38_ : 
                (N326)? speculative_queue_q_1__data__38_ : 
                (N325)? speculative_queue_q_2__data__38_ : 
                (N327)? speculative_queue_q_3__data__38_ : 1'b0;
  assign N410 = (N324)? speculative_queue_q_0__data__37_ : 
                (N326)? speculative_queue_q_1__data__37_ : 
                (N325)? speculative_queue_q_2__data__37_ : 
                (N327)? speculative_queue_q_3__data__37_ : 1'b0;
  assign N411 = (N324)? speculative_queue_q_0__data__36_ : 
                (N326)? speculative_queue_q_1__data__36_ : 
                (N325)? speculative_queue_q_2__data__36_ : 
                (N327)? speculative_queue_q_3__data__36_ : 1'b0;
  assign N412 = (N324)? speculative_queue_q_0__data__35_ : 
                (N326)? speculative_queue_q_1__data__35_ : 
                (N325)? speculative_queue_q_2__data__35_ : 
                (N327)? speculative_queue_q_3__data__35_ : 1'b0;
  assign N413 = (N324)? speculative_queue_q_0__data__34_ : 
                (N326)? speculative_queue_q_1__data__34_ : 
                (N325)? speculative_queue_q_2__data__34_ : 
                (N327)? speculative_queue_q_3__data__34_ : 1'b0;
  assign N414 = (N324)? speculative_queue_q_0__data__33_ : 
                (N326)? speculative_queue_q_1__data__33_ : 
                (N325)? speculative_queue_q_2__data__33_ : 
                (N327)? speculative_queue_q_3__data__33_ : 1'b0;
  assign N415 = (N324)? speculative_queue_q_0__data__32_ : 
                (N326)? speculative_queue_q_1__data__32_ : 
                (N325)? speculative_queue_q_2__data__32_ : 
                (N327)? speculative_queue_q_3__data__32_ : 1'b0;
  assign N416 = (N324)? speculative_queue_q_0__data__31_ : 
                (N326)? speculative_queue_q_1__data__31_ : 
                (N325)? speculative_queue_q_2__data__31_ : 
                (N327)? speculative_queue_q_3__data__31_ : 1'b0;
  assign N417 = (N324)? speculative_queue_q_0__data__30_ : 
                (N326)? speculative_queue_q_1__data__30_ : 
                (N325)? speculative_queue_q_2__data__30_ : 
                (N327)? speculative_queue_q_3__data__30_ : 1'b0;
  assign N418 = (N324)? speculative_queue_q_0__data__29_ : 
                (N326)? speculative_queue_q_1__data__29_ : 
                (N325)? speculative_queue_q_2__data__29_ : 
                (N327)? speculative_queue_q_3__data__29_ : 1'b0;
  assign N419 = (N324)? speculative_queue_q_0__data__28_ : 
                (N326)? speculative_queue_q_1__data__28_ : 
                (N325)? speculative_queue_q_2__data__28_ : 
                (N327)? speculative_queue_q_3__data__28_ : 1'b0;
  assign N420 = (N324)? speculative_queue_q_0__data__27_ : 
                (N326)? speculative_queue_q_1__data__27_ : 
                (N325)? speculative_queue_q_2__data__27_ : 
                (N327)? speculative_queue_q_3__data__27_ : 1'b0;
  assign N421 = (N324)? speculative_queue_q_0__data__26_ : 
                (N326)? speculative_queue_q_1__data__26_ : 
                (N325)? speculative_queue_q_2__data__26_ : 
                (N327)? speculative_queue_q_3__data__26_ : 1'b0;
  assign N422 = (N324)? speculative_queue_q_0__data__25_ : 
                (N326)? speculative_queue_q_1__data__25_ : 
                (N325)? speculative_queue_q_2__data__25_ : 
                (N327)? speculative_queue_q_3__data__25_ : 1'b0;
  assign N423 = (N324)? speculative_queue_q_0__data__24_ : 
                (N326)? speculative_queue_q_1__data__24_ : 
                (N325)? speculative_queue_q_2__data__24_ : 
                (N327)? speculative_queue_q_3__data__24_ : 1'b0;
  assign N424 = (N324)? speculative_queue_q_0__data__23_ : 
                (N326)? speculative_queue_q_1__data__23_ : 
                (N325)? speculative_queue_q_2__data__23_ : 
                (N327)? speculative_queue_q_3__data__23_ : 1'b0;
  assign N425 = (N324)? speculative_queue_q_0__data__22_ : 
                (N326)? speculative_queue_q_1__data__22_ : 
                (N325)? speculative_queue_q_2__data__22_ : 
                (N327)? speculative_queue_q_3__data__22_ : 1'b0;
  assign N426 = (N324)? speculative_queue_q_0__data__21_ : 
                (N326)? speculative_queue_q_1__data__21_ : 
                (N325)? speculative_queue_q_2__data__21_ : 
                (N327)? speculative_queue_q_3__data__21_ : 1'b0;
  assign N427 = (N324)? speculative_queue_q_0__data__20_ : 
                (N326)? speculative_queue_q_1__data__20_ : 
                (N325)? speculative_queue_q_2__data__20_ : 
                (N327)? speculative_queue_q_3__data__20_ : 1'b0;
  assign N428 = (N324)? speculative_queue_q_0__data__19_ : 
                (N326)? speculative_queue_q_1__data__19_ : 
                (N325)? speculative_queue_q_2__data__19_ : 
                (N327)? speculative_queue_q_3__data__19_ : 1'b0;
  assign N429 = (N324)? speculative_queue_q_0__data__18_ : 
                (N326)? speculative_queue_q_1__data__18_ : 
                (N325)? speculative_queue_q_2__data__18_ : 
                (N327)? speculative_queue_q_3__data__18_ : 1'b0;
  assign N430 = (N324)? speculative_queue_q_0__data__17_ : 
                (N326)? speculative_queue_q_1__data__17_ : 
                (N325)? speculative_queue_q_2__data__17_ : 
                (N327)? speculative_queue_q_3__data__17_ : 1'b0;
  assign N431 = (N324)? speculative_queue_q_0__data__16_ : 
                (N326)? speculative_queue_q_1__data__16_ : 
                (N325)? speculative_queue_q_2__data__16_ : 
                (N327)? speculative_queue_q_3__data__16_ : 1'b0;
  assign N432 = (N324)? speculative_queue_q_0__data__15_ : 
                (N326)? speculative_queue_q_1__data__15_ : 
                (N325)? speculative_queue_q_2__data__15_ : 
                (N327)? speculative_queue_q_3__data__15_ : 1'b0;
  assign N433 = (N324)? speculative_queue_q_0__data__14_ : 
                (N326)? speculative_queue_q_1__data__14_ : 
                (N325)? speculative_queue_q_2__data__14_ : 
                (N327)? speculative_queue_q_3__data__14_ : 1'b0;
  assign N434 = (N324)? speculative_queue_q_0__data__13_ : 
                (N326)? speculative_queue_q_1__data__13_ : 
                (N325)? speculative_queue_q_2__data__13_ : 
                (N327)? speculative_queue_q_3__data__13_ : 1'b0;
  assign N435 = (N324)? speculative_queue_q_0__data__12_ : 
                (N326)? speculative_queue_q_1__data__12_ : 
                (N325)? speculative_queue_q_2__data__12_ : 
                (N327)? speculative_queue_q_3__data__12_ : 1'b0;
  assign N436 = (N324)? speculative_queue_q_0__data__11_ : 
                (N326)? speculative_queue_q_1__data__11_ : 
                (N325)? speculative_queue_q_2__data__11_ : 
                (N327)? speculative_queue_q_3__data__11_ : 1'b0;
  assign N437 = (N324)? speculative_queue_q_0__data__10_ : 
                (N326)? speculative_queue_q_1__data__10_ : 
                (N325)? speculative_queue_q_2__data__10_ : 
                (N327)? speculative_queue_q_3__data__10_ : 1'b0;
  assign N438 = (N324)? speculative_queue_q_0__data__9_ : 
                (N326)? speculative_queue_q_1__data__9_ : 
                (N325)? speculative_queue_q_2__data__9_ : 
                (N327)? speculative_queue_q_3__data__9_ : 1'b0;
  assign N439 = (N324)? speculative_queue_q_0__data__8_ : 
                (N326)? speculative_queue_q_1__data__8_ : 
                (N325)? speculative_queue_q_2__data__8_ : 
                (N327)? speculative_queue_q_3__data__8_ : 1'b0;
  assign N440 = (N324)? speculative_queue_q_0__data__7_ : 
                (N326)? speculative_queue_q_1__data__7_ : 
                (N325)? speculative_queue_q_2__data__7_ : 
                (N327)? speculative_queue_q_3__data__7_ : 1'b0;
  assign N441 = (N324)? speculative_queue_q_0__data__6_ : 
                (N326)? speculative_queue_q_1__data__6_ : 
                (N325)? speculative_queue_q_2__data__6_ : 
                (N327)? speculative_queue_q_3__data__6_ : 1'b0;
  assign N442 = (N324)? speculative_queue_q_0__data__5_ : 
                (N326)? speculative_queue_q_1__data__5_ : 
                (N325)? speculative_queue_q_2__data__5_ : 
                (N327)? speculative_queue_q_3__data__5_ : 1'b0;
  assign N443 = (N324)? speculative_queue_q_0__data__4_ : 
                (N326)? speculative_queue_q_1__data__4_ : 
                (N325)? speculative_queue_q_2__data__4_ : 
                (N327)? speculative_queue_q_3__data__4_ : 1'b0;
  assign N444 = (N324)? speculative_queue_q_0__data__3_ : 
                (N326)? speculative_queue_q_1__data__3_ : 
                (N325)? speculative_queue_q_2__data__3_ : 
                (N327)? speculative_queue_q_3__data__3_ : 1'b0;
  assign N445 = (N324)? speculative_queue_q_0__data__2_ : 
                (N326)? speculative_queue_q_1__data__2_ : 
                (N325)? speculative_queue_q_2__data__2_ : 
                (N327)? speculative_queue_q_3__data__2_ : 1'b0;
  assign N446 = (N324)? speculative_queue_q_0__data__1_ : 
                (N326)? speculative_queue_q_1__data__1_ : 
                (N325)? speculative_queue_q_2__data__1_ : 
                (N327)? speculative_queue_q_3__data__1_ : 1'b0;
  assign N447 = (N324)? speculative_queue_q_0__data__0_ : 
                (N326)? speculative_queue_q_1__data__0_ : 
                (N325)? speculative_queue_q_2__data__0_ : 
                (N327)? speculative_queue_q_3__data__0_ : 1'b0;
  assign N448 = (N324)? speculative_queue_q_0__be__7_ : 
                (N326)? speculative_queue_q_1__be__7_ : 
                (N325)? speculative_queue_q_2__be__7_ : 
                (N327)? speculative_queue_q_3__be__7_ : 1'b0;
  assign N449 = (N324)? speculative_queue_q_0__be__6_ : 
                (N326)? speculative_queue_q_1__be__6_ : 
                (N325)? speculative_queue_q_2__be__6_ : 
                (N327)? speculative_queue_q_3__be__6_ : 1'b0;
  assign N450 = (N324)? speculative_queue_q_0__be__5_ : 
                (N326)? speculative_queue_q_1__be__5_ : 
                (N325)? speculative_queue_q_2__be__5_ : 
                (N327)? speculative_queue_q_3__be__5_ : 1'b0;
  assign N451 = (N324)? speculative_queue_q_0__be__4_ : 
                (N326)? speculative_queue_q_1__be__4_ : 
                (N325)? speculative_queue_q_2__be__4_ : 
                (N327)? speculative_queue_q_3__be__4_ : 1'b0;
  assign N452 = (N324)? speculative_queue_q_0__be__3_ : 
                (N326)? speculative_queue_q_1__be__3_ : 
                (N325)? speculative_queue_q_2__be__3_ : 
                (N327)? speculative_queue_q_3__be__3_ : 1'b0;
  assign N453 = (N324)? speculative_queue_q_0__be__2_ : 
                (N326)? speculative_queue_q_1__be__2_ : 
                (N325)? speculative_queue_q_2__be__2_ : 
                (N327)? speculative_queue_q_3__be__2_ : 1'b0;
  assign N454 = (N324)? speculative_queue_q_0__be__1_ : 
                (N326)? speculative_queue_q_1__be__1_ : 
                (N325)? speculative_queue_q_2__be__1_ : 
                (N327)? speculative_queue_q_3__be__1_ : 1'b0;
  assign N455 = (N324)? speculative_queue_q_0__be__0_ : 
                (N326)? speculative_queue_q_1__be__0_ : 
                (N325)? speculative_queue_q_2__be__0_ : 
                (N327)? speculative_queue_q_3__be__0_ : 1'b0;
  assign N456 = (N324)? speculative_queue_q_0__data_size__1_ : 
                (N326)? speculative_queue_q_1__data_size__1_ : 
                (N325)? speculative_queue_q_2__data_size__1_ : 
                (N327)? speculative_queue_q_3__data_size__1_ : 1'b0;
  assign N457 = (N324)? speculative_queue_q_0__data_size__0_ : 
                (N326)? speculative_queue_q_1__data_size__0_ : 
                (N325)? speculative_queue_q_2__data_size__0_ : 
                (N327)? speculative_queue_q_3__data_size__0_ : 1'b0;
  assign N458 = (N324)? speculative_queue_q_0__valid_ : 
                (N326)? speculative_queue_q_1__valid_ : 
                (N325)? speculative_queue_q_2__valid_ : 
                (N327)? speculative_queue_q_3__valid_ : 1'b0;
  assign N490 = page_offset_i[11:3] == { commit_queue_q_0__address__11_, commit_queue_q_0__address__10_, commit_queue_q_0__address__9_, commit_queue_q_0__address__8_, commit_queue_q_0__address__7_, commit_queue_q_0__address__6_, commit_queue_q_0__address__5_, commit_queue_q_0__address__4_, commit_queue_q_0__address__3_ };
  assign N496 = page_offset_i[11:3] == { commit_queue_q_1__address__11_, commit_queue_q_1__address__10_, commit_queue_q_1__address__9_, commit_queue_q_1__address__8_, commit_queue_q_1__address__7_, commit_queue_q_1__address__6_, commit_queue_q_1__address__5_, commit_queue_q_1__address__4_, commit_queue_q_1__address__3_ };
  assign N504 = page_offset_i[11:3] == { commit_queue_q_2__address__11_, commit_queue_q_2__address__10_, commit_queue_q_2__address__9_, commit_queue_q_2__address__8_, commit_queue_q_2__address__7_, commit_queue_q_2__address__6_, commit_queue_q_2__address__5_, commit_queue_q_2__address__4_, commit_queue_q_2__address__3_ };
  assign N512 = page_offset_i[11:3] == { commit_queue_q_3__address__11_, commit_queue_q_3__address__10_, commit_queue_q_3__address__9_, commit_queue_q_3__address__8_, commit_queue_q_3__address__7_, commit_queue_q_3__address__6_, commit_queue_q_3__address__5_, commit_queue_q_3__address__4_, commit_queue_q_3__address__3_ };
  assign N520 = page_offset_i[11:3] == { commit_queue_q_4__address__11_, commit_queue_q_4__address__10_, commit_queue_q_4__address__9_, commit_queue_q_4__address__8_, commit_queue_q_4__address__7_, commit_queue_q_4__address__6_, commit_queue_q_4__address__5_, commit_queue_q_4__address__4_, commit_queue_q_4__address__3_ };
  assign N528 = page_offset_i[11:3] == { commit_queue_q_5__address__11_, commit_queue_q_5__address__10_, commit_queue_q_5__address__9_, commit_queue_q_5__address__8_, commit_queue_q_5__address__7_, commit_queue_q_5__address__6_, commit_queue_q_5__address__5_, commit_queue_q_5__address__4_, commit_queue_q_5__address__3_ };
  assign N536 = page_offset_i[11:3] == { commit_queue_q_6__address__11_, commit_queue_q_6__address__10_, commit_queue_q_6__address__9_, commit_queue_q_6__address__8_, commit_queue_q_6__address__7_, commit_queue_q_6__address__6_, commit_queue_q_6__address__5_, commit_queue_q_6__address__4_, commit_queue_q_6__address__3_ };
  assign N543 = page_offset_i[11:3] == { commit_queue_q_7__address__11_, commit_queue_q_7__address__10_, commit_queue_q_7__address__9_, commit_queue_q_7__address__8_, commit_queue_q_7__address__7_, commit_queue_q_7__address__6_, commit_queue_q_7__address__5_, commit_queue_q_7__address__4_, commit_queue_q_7__address__3_ };
  assign N567 = page_offset_i[11:3] == { speculative_queue_q_0__address__11_, speculative_queue_q_0__address__10_, speculative_queue_q_0__address__9_, speculative_queue_q_0__address__8_, speculative_queue_q_0__address__7_, speculative_queue_q_0__address__6_, speculative_queue_q_0__address__5_, speculative_queue_q_0__address__4_, speculative_queue_q_0__address__3_ };
  assign N575 = page_offset_i[11:3] == { speculative_queue_q_1__address__11_, speculative_queue_q_1__address__10_, speculative_queue_q_1__address__9_, speculative_queue_q_1__address__8_, speculative_queue_q_1__address__7_, speculative_queue_q_1__address__6_, speculative_queue_q_1__address__5_, speculative_queue_q_1__address__4_, speculative_queue_q_1__address__3_ };
  assign N583 = page_offset_i[11:3] == { speculative_queue_q_2__address__11_, speculative_queue_q_2__address__10_, speculative_queue_q_2__address__9_, speculative_queue_q_2__address__8_, speculative_queue_q_2__address__7_, speculative_queue_q_2__address__6_, speculative_queue_q_2__address__5_, speculative_queue_q_2__address__4_, speculative_queue_q_2__address__3_ };
  assign N590 = page_offset_i[11:3] == { speculative_queue_q_3__address__11_, speculative_queue_q_3__address__10_, speculative_queue_q_3__address__9_, speculative_queue_q_3__address__8_, speculative_queue_q_3__address__7_, speculative_queue_q_3__address__6_, speculative_queue_q_3__address__5_, speculative_queue_q_3__address__4_, speculative_queue_q_3__address__3_ };
  assign N602 = page_offset_i[11:3] == paddr_i[11:3];

  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_write_pointer_q[1] <= 1'b0;
    end else if(N607) begin
      speculative_write_pointer_q[1] <= speculative_write_pointer_n[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_write_pointer_q[0] <= 1'b0;
    end else if(N607) begin
      speculative_write_pointer_q[0] <= speculative_write_pointer_n[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_status_cnt_q[2] <= 1'b0;
    end else if(1'b1) begin
      speculative_status_cnt_q[2] <= speculative_status_cnt_n[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_status_cnt_q[1] <= 1'b0;
    end else if(1'b1) begin
      speculative_status_cnt_q[1] <= speculative_status_cnt_n[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_status_cnt_q[0] <= 1'b0;
    end else if(1'b1) begin
      speculative_status_cnt_q[0] <= speculative_status_cnt_n[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__55_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__55_ <= paddr_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__54_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__54_ <= paddr_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__53_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__53_ <= paddr_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__52_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__52_ <= paddr_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__51_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__51_ <= paddr_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__50_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__50_ <= paddr_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__49_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__49_ <= paddr_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__48_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__48_ <= paddr_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__47_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__47_ <= paddr_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__46_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__46_ <= paddr_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__45_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__45_ <= paddr_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__44_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__44_ <= paddr_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__43_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__43_ <= paddr_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__42_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__42_ <= paddr_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__41_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__41_ <= paddr_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__40_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__40_ <= paddr_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__39_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__39_ <= paddr_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__38_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__38_ <= paddr_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__37_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__37_ <= paddr_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__36_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__36_ <= paddr_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__35_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__35_ <= paddr_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__34_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__34_ <= paddr_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__33_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__33_ <= paddr_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__32_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__32_ <= paddr_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__31_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__31_ <= paddr_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__30_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__30_ <= paddr_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__29_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__29_ <= paddr_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__28_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__28_ <= paddr_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__27_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__27_ <= paddr_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__26_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__26_ <= paddr_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__25_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__25_ <= paddr_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__24_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__24_ <= paddr_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__23_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__23_ <= paddr_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__22_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__22_ <= paddr_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__21_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__21_ <= paddr_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__20_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__20_ <= paddr_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__19_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__19_ <= paddr_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__18_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__18_ <= paddr_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__17_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__17_ <= paddr_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__16_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__16_ <= paddr_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__15_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__15_ <= paddr_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__14_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__14_ <= paddr_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__13_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__13_ <= paddr_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__12_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__12_ <= paddr_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__11_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__11_ <= paddr_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__10_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__10_ <= paddr_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__9_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__9_ <= paddr_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__8_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__8_ <= paddr_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__7_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__7_ <= paddr_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__6_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__6_ <= paddr_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__5_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__5_ <= paddr_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__4_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__4_ <= paddr_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__3_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__3_ <= paddr_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__2_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__2_ <= paddr_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__1_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__1_ <= paddr_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__address__0_ <= 1'b0;
    end else if(N610) begin
      speculative_queue_q_3__address__0_ <= paddr_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__63_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__63_ <= data_i[63];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__62_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__62_ <= data_i[62];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__61_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__61_ <= data_i[61];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__60_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__60_ <= data_i[60];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__59_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__59_ <= data_i[59];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__58_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__58_ <= data_i[58];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__57_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__57_ <= data_i[57];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__56_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__56_ <= data_i[56];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__55_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__55_ <= data_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__54_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__54_ <= data_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__53_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__53_ <= data_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__52_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__52_ <= data_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__51_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__51_ <= data_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__50_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__50_ <= data_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__49_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__49_ <= data_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__48_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__48_ <= data_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__47_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__47_ <= data_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__46_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__46_ <= data_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__45_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__45_ <= data_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__44_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__44_ <= data_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__43_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__43_ <= data_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__42_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__42_ <= data_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__41_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__41_ <= data_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__40_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__40_ <= data_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__39_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__39_ <= data_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__38_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__38_ <= data_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__37_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__37_ <= data_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__36_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__36_ <= data_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__35_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__35_ <= data_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__34_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__34_ <= data_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__33_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__33_ <= data_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__32_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__32_ <= data_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__31_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__31_ <= data_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__30_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__30_ <= data_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__29_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__29_ <= data_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__28_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__28_ <= data_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__27_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__27_ <= data_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__26_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__26_ <= data_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__25_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__25_ <= data_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__24_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__24_ <= data_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__23_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__23_ <= data_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__22_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__22_ <= data_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__21_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__21_ <= data_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__20_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__20_ <= data_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__19_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__19_ <= data_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__18_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__18_ <= data_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__17_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__17_ <= data_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__16_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__16_ <= data_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__15_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__15_ <= data_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__14_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__14_ <= data_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__13_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__13_ <= data_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__12_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__12_ <= data_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__11_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__11_ <= data_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__10_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__10_ <= data_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__9_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__9_ <= data_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__8_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__8_ <= data_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__7_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__7_ <= data_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__6_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__6_ <= data_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__5_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__5_ <= data_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__4_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__4_ <= data_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__3_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__3_ <= data_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__2_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__2_ <= data_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__1_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__1_ <= data_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data__0_ <= 1'b0;
    end else if(N613) begin
      speculative_queue_q_3__data__0_ <= data_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__7_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__7_ <= be_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__6_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__6_ <= be_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__5_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__5_ <= be_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__4_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__4_ <= be_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__3_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__3_ <= be_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__2_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__2_ <= be_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__1_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__1_ <= be_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__be__0_ <= 1'b0;
    end else if(N616) begin
      speculative_queue_q_3__be__0_ <= be_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data_size__1_ <= 1'b0;
    end else if(N619) begin
      speculative_queue_q_3__data_size__1_ <= data_size_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__data_size__0_ <= 1'b0;
    end else if(N619) begin
      speculative_queue_q_3__data_size__0_ <= data_size_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_3__valid_ <= 1'b0;
    end else if(1'b1) begin
      speculative_queue_q_3__valid_ <= speculative_queue_n_3__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__55_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__55_ <= paddr_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__54_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__54_ <= paddr_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__53_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__53_ <= paddr_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__52_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__52_ <= paddr_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__51_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__51_ <= paddr_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__50_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__50_ <= paddr_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__49_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__49_ <= paddr_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__48_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__48_ <= paddr_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__47_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__47_ <= paddr_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__46_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__46_ <= paddr_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__45_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__45_ <= paddr_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__44_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__44_ <= paddr_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__43_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__43_ <= paddr_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__42_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__42_ <= paddr_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__41_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__41_ <= paddr_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__40_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__40_ <= paddr_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__39_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__39_ <= paddr_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__38_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__38_ <= paddr_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__37_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__37_ <= paddr_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__36_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__36_ <= paddr_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__35_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__35_ <= paddr_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__34_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__34_ <= paddr_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__33_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__33_ <= paddr_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__32_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__32_ <= paddr_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__31_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__31_ <= paddr_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__30_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__30_ <= paddr_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__29_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__29_ <= paddr_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__28_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__28_ <= paddr_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__27_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__27_ <= paddr_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__26_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__26_ <= paddr_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__25_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__25_ <= paddr_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__24_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__24_ <= paddr_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__23_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__23_ <= paddr_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__22_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__22_ <= paddr_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__21_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__21_ <= paddr_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__20_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__20_ <= paddr_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__19_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__19_ <= paddr_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__18_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__18_ <= paddr_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__17_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__17_ <= paddr_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__16_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__16_ <= paddr_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__15_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__15_ <= paddr_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__14_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__14_ <= paddr_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__13_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__13_ <= paddr_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__12_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__12_ <= paddr_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__11_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__11_ <= paddr_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__10_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__10_ <= paddr_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__9_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__9_ <= paddr_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__8_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__8_ <= paddr_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__7_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__7_ <= paddr_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__6_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__6_ <= paddr_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__5_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__5_ <= paddr_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__4_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__4_ <= paddr_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__3_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__3_ <= paddr_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__2_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__2_ <= paddr_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__1_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__1_ <= paddr_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__address__0_ <= 1'b0;
    end else if(N622) begin
      speculative_queue_q_2__address__0_ <= paddr_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__63_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__63_ <= data_i[63];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__62_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__62_ <= data_i[62];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__61_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__61_ <= data_i[61];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__60_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__60_ <= data_i[60];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__59_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__59_ <= data_i[59];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__58_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__58_ <= data_i[58];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__57_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__57_ <= data_i[57];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__56_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__56_ <= data_i[56];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__55_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__55_ <= data_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__54_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__54_ <= data_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__53_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__53_ <= data_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__52_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__52_ <= data_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__51_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__51_ <= data_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__50_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__50_ <= data_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__49_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__49_ <= data_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__48_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__48_ <= data_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__47_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__47_ <= data_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__46_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__46_ <= data_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__45_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__45_ <= data_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__44_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__44_ <= data_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__43_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__43_ <= data_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__42_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__42_ <= data_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__41_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__41_ <= data_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__40_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__40_ <= data_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__39_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__39_ <= data_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__38_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__38_ <= data_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__37_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__37_ <= data_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__36_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__36_ <= data_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__35_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__35_ <= data_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__34_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__34_ <= data_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__33_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__33_ <= data_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__32_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__32_ <= data_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__31_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__31_ <= data_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__30_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__30_ <= data_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__29_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__29_ <= data_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__28_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__28_ <= data_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__27_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__27_ <= data_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__26_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__26_ <= data_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__25_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__25_ <= data_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__24_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__24_ <= data_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__23_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__23_ <= data_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__22_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__22_ <= data_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__21_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__21_ <= data_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__20_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__20_ <= data_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__19_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__19_ <= data_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__18_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__18_ <= data_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__17_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__17_ <= data_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__16_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__16_ <= data_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__15_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__15_ <= data_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__14_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__14_ <= data_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__13_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__13_ <= data_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__12_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__12_ <= data_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__11_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__11_ <= data_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__10_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__10_ <= data_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__9_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__9_ <= data_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__8_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__8_ <= data_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__7_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__7_ <= data_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__6_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__6_ <= data_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__5_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__5_ <= data_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__4_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__4_ <= data_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__3_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__3_ <= data_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__2_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__2_ <= data_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__1_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__1_ <= data_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data__0_ <= 1'b0;
    end else if(N625) begin
      speculative_queue_q_2__data__0_ <= data_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__7_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__7_ <= be_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__6_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__6_ <= be_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__5_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__5_ <= be_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__4_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__4_ <= be_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__3_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__3_ <= be_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__2_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__2_ <= be_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__1_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__1_ <= be_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__be__0_ <= 1'b0;
    end else if(N628) begin
      speculative_queue_q_2__be__0_ <= be_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data_size__1_ <= 1'b0;
    end else if(N631) begin
      speculative_queue_q_2__data_size__1_ <= data_size_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__data_size__0_ <= 1'b0;
    end else if(N631) begin
      speculative_queue_q_2__data_size__0_ <= data_size_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_2__valid_ <= 1'b0;
    end else if(1'b1) begin
      speculative_queue_q_2__valid_ <= speculative_queue_n_2__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__55_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__55_ <= paddr_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__54_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__54_ <= paddr_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__53_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__53_ <= paddr_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__52_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__52_ <= paddr_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__51_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__51_ <= paddr_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__50_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__50_ <= paddr_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__49_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__49_ <= paddr_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__48_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__48_ <= paddr_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__47_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__47_ <= paddr_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__46_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__46_ <= paddr_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__45_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__45_ <= paddr_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__44_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__44_ <= paddr_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__43_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__43_ <= paddr_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__42_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__42_ <= paddr_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__41_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__41_ <= paddr_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__40_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__40_ <= paddr_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__39_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__39_ <= paddr_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__38_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__38_ <= paddr_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__37_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__37_ <= paddr_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__36_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__36_ <= paddr_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__35_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__35_ <= paddr_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__34_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__34_ <= paddr_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__33_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__33_ <= paddr_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__32_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__32_ <= paddr_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__31_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__31_ <= paddr_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__30_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__30_ <= paddr_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__29_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__29_ <= paddr_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__28_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__28_ <= paddr_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__27_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__27_ <= paddr_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__26_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__26_ <= paddr_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__25_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__25_ <= paddr_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__24_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__24_ <= paddr_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__23_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__23_ <= paddr_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__22_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__22_ <= paddr_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__21_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__21_ <= paddr_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__20_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__20_ <= paddr_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__19_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__19_ <= paddr_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__18_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__18_ <= paddr_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__17_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__17_ <= paddr_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__16_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__16_ <= paddr_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__15_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__15_ <= paddr_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__14_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__14_ <= paddr_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__13_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__13_ <= paddr_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__12_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__12_ <= paddr_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__11_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__11_ <= paddr_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__10_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__10_ <= paddr_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__9_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__9_ <= paddr_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__8_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__8_ <= paddr_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__7_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__7_ <= paddr_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__6_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__6_ <= paddr_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__5_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__5_ <= paddr_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__4_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__4_ <= paddr_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__3_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__3_ <= paddr_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__2_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__2_ <= paddr_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__1_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__1_ <= paddr_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__address__0_ <= 1'b0;
    end else if(N634) begin
      speculative_queue_q_1__address__0_ <= paddr_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__63_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__63_ <= data_i[63];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__62_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__62_ <= data_i[62];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__61_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__61_ <= data_i[61];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__60_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__60_ <= data_i[60];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__59_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__59_ <= data_i[59];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__58_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__58_ <= data_i[58];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__57_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__57_ <= data_i[57];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__56_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__56_ <= data_i[56];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__55_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__55_ <= data_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__54_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__54_ <= data_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__53_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__53_ <= data_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__52_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__52_ <= data_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__51_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__51_ <= data_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__50_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__50_ <= data_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__49_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__49_ <= data_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__48_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__48_ <= data_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__47_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__47_ <= data_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__46_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__46_ <= data_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__45_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__45_ <= data_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__44_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__44_ <= data_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__43_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__43_ <= data_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__42_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__42_ <= data_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__41_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__41_ <= data_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__40_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__40_ <= data_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__39_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__39_ <= data_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__38_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__38_ <= data_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__37_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__37_ <= data_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__36_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__36_ <= data_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__35_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__35_ <= data_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__34_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__34_ <= data_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__33_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__33_ <= data_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__32_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__32_ <= data_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__31_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__31_ <= data_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__30_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__30_ <= data_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__29_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__29_ <= data_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__28_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__28_ <= data_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__27_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__27_ <= data_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__26_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__26_ <= data_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__25_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__25_ <= data_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__24_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__24_ <= data_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__23_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__23_ <= data_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__22_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__22_ <= data_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__21_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__21_ <= data_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__20_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__20_ <= data_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__19_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__19_ <= data_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__18_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__18_ <= data_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__17_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__17_ <= data_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__16_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__16_ <= data_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__15_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__15_ <= data_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__14_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__14_ <= data_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__13_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__13_ <= data_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__12_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__12_ <= data_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__11_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__11_ <= data_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__10_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__10_ <= data_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__9_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__9_ <= data_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__8_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__8_ <= data_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__7_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__7_ <= data_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__6_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__6_ <= data_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__5_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__5_ <= data_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__4_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__4_ <= data_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__3_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__3_ <= data_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__2_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__2_ <= data_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__1_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__1_ <= data_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data__0_ <= 1'b0;
    end else if(N637) begin
      speculative_queue_q_1__data__0_ <= data_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__7_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__7_ <= be_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__6_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__6_ <= be_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__5_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__5_ <= be_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__4_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__4_ <= be_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__3_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__3_ <= be_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__2_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__2_ <= be_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__1_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__1_ <= be_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__be__0_ <= 1'b0;
    end else if(N640) begin
      speculative_queue_q_1__be__0_ <= be_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data_size__1_ <= 1'b0;
    end else if(N643) begin
      speculative_queue_q_1__data_size__1_ <= data_size_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__data_size__0_ <= 1'b0;
    end else if(N643) begin
      speculative_queue_q_1__data_size__0_ <= data_size_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_1__valid_ <= 1'b0;
    end else if(1'b1) begin
      speculative_queue_q_1__valid_ <= speculative_queue_n_1__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__55_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__55_ <= paddr_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__54_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__54_ <= paddr_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__53_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__53_ <= paddr_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__52_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__52_ <= paddr_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__51_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__51_ <= paddr_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__50_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__50_ <= paddr_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__49_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__49_ <= paddr_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__48_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__48_ <= paddr_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__47_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__47_ <= paddr_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__46_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__46_ <= paddr_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__45_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__45_ <= paddr_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__44_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__44_ <= paddr_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__43_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__43_ <= paddr_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__42_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__42_ <= paddr_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__41_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__41_ <= paddr_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__40_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__40_ <= paddr_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__39_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__39_ <= paddr_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__38_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__38_ <= paddr_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__37_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__37_ <= paddr_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__36_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__36_ <= paddr_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__35_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__35_ <= paddr_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__34_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__34_ <= paddr_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__33_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__33_ <= paddr_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__32_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__32_ <= paddr_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__31_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__31_ <= paddr_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__30_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__30_ <= paddr_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__29_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__29_ <= paddr_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__28_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__28_ <= paddr_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__27_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__27_ <= paddr_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__26_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__26_ <= paddr_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__25_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__25_ <= paddr_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__24_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__24_ <= paddr_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__23_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__23_ <= paddr_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__22_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__22_ <= paddr_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__21_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__21_ <= paddr_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__20_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__20_ <= paddr_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__19_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__19_ <= paddr_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__18_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__18_ <= paddr_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__17_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__17_ <= paddr_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__16_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__16_ <= paddr_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__15_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__15_ <= paddr_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__14_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__14_ <= paddr_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__13_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__13_ <= paddr_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__12_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__12_ <= paddr_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__11_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__11_ <= paddr_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__10_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__10_ <= paddr_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__9_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__9_ <= paddr_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__8_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__8_ <= paddr_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__7_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__7_ <= paddr_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__6_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__6_ <= paddr_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__5_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__5_ <= paddr_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__4_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__4_ <= paddr_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__3_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__3_ <= paddr_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__2_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__2_ <= paddr_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__1_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__1_ <= paddr_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__address__0_ <= 1'b0;
    end else if(N646) begin
      speculative_queue_q_0__address__0_ <= paddr_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__63_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__63_ <= data_i[63];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__62_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__62_ <= data_i[62];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__61_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__61_ <= data_i[61];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__60_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__60_ <= data_i[60];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__59_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__59_ <= data_i[59];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__58_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__58_ <= data_i[58];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__57_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__57_ <= data_i[57];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__56_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__56_ <= data_i[56];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__55_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__55_ <= data_i[55];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__54_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__54_ <= data_i[54];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__53_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__53_ <= data_i[53];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__52_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__52_ <= data_i[52];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__51_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__51_ <= data_i[51];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__50_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__50_ <= data_i[50];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__49_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__49_ <= data_i[49];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__48_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__48_ <= data_i[48];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__47_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__47_ <= data_i[47];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__46_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__46_ <= data_i[46];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__45_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__45_ <= data_i[45];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__44_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__44_ <= data_i[44];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__43_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__43_ <= data_i[43];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__42_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__42_ <= data_i[42];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__41_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__41_ <= data_i[41];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__40_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__40_ <= data_i[40];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__39_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__39_ <= data_i[39];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__38_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__38_ <= data_i[38];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__37_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__37_ <= data_i[37];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__36_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__36_ <= data_i[36];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__35_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__35_ <= data_i[35];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__34_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__34_ <= data_i[34];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__33_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__33_ <= data_i[33];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__32_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__32_ <= data_i[32];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__31_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__31_ <= data_i[31];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__30_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__30_ <= data_i[30];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__29_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__29_ <= data_i[29];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__28_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__28_ <= data_i[28];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__27_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__27_ <= data_i[27];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__26_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__26_ <= data_i[26];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__25_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__25_ <= data_i[25];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__24_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__24_ <= data_i[24];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__23_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__23_ <= data_i[23];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__22_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__22_ <= data_i[22];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__21_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__21_ <= data_i[21];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__20_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__20_ <= data_i[20];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__19_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__19_ <= data_i[19];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__18_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__18_ <= data_i[18];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__17_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__17_ <= data_i[17];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__16_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__16_ <= data_i[16];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__15_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__15_ <= data_i[15];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__14_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__14_ <= data_i[14];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__13_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__13_ <= data_i[13];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__12_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__12_ <= data_i[12];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__11_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__11_ <= data_i[11];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__10_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__10_ <= data_i[10];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__9_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__9_ <= data_i[9];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__8_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__8_ <= data_i[8];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__7_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__7_ <= data_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__6_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__6_ <= data_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__5_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__5_ <= data_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__4_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__4_ <= data_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__3_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__3_ <= data_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__2_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__2_ <= data_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__1_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__1_ <= data_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data__0_ <= 1'b0;
    end else if(N649) begin
      speculative_queue_q_0__data__0_ <= data_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__7_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__7_ <= be_i[7];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__6_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__6_ <= be_i[6];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__5_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__5_ <= be_i[5];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__4_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__4_ <= be_i[4];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__3_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__3_ <= be_i[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__2_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__2_ <= be_i[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__1_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__1_ <= be_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__be__0_ <= 1'b0;
    end else if(N652) begin
      speculative_queue_q_0__be__0_ <= be_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data_size__1_ <= 1'b0;
    end else if(N655) begin
      speculative_queue_q_0__data_size__1_ <= data_size_i[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__data_size__0_ <= 1'b0;
    end else if(N655) begin
      speculative_queue_q_0__data_size__0_ <= data_size_i[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_queue_q_0__valid_ <= 1'b0;
    end else if(1'b1) begin
      speculative_queue_q_0__valid_ <= speculative_queue_n_0__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_read_pointer_q[1] <= 1'b0;
    end else if(commit_i) begin
      speculative_read_pointer_q[1] <= N186;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      speculative_read_pointer_q[0] <= 1'b0;
    end else if(commit_i) begin
      speculative_read_pointer_q[0] <= N185;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_write_pointer_q[2] <= 1'b0;
    end else if(commit_i) begin
      commit_write_pointer_q[2] <= N485;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_write_pointer_q[1] <= 1'b0;
    end else if(commit_i) begin
      commit_write_pointer_q[1] <= N484;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_write_pointer_q[0] <= 1'b0;
    end else if(commit_i) begin
      commit_write_pointer_q[0] <= N483;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_status_cnt_q[3] <= 1'b0;
    end else if(1'b1) begin
      commit_status_cnt_q[3] <= commit_status_cnt_n[3];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_status_cnt_q[2] <= 1'b0;
    end else if(1'b1) begin
      commit_status_cnt_q[2] <= commit_status_cnt_n[2];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_status_cnt_q[1] <= 1'b0;
    end else if(1'b1) begin
      commit_status_cnt_q[1] <= commit_status_cnt_n[1];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_status_cnt_q[0] <= 1'b0;
    end else if(1'b1) begin
      commit_status_cnt_q[0] <= commit_status_cnt_n[0];
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__55_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__54_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__53_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__52_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__51_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__50_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__49_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__48_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__47_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__46_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__45_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__44_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__43_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__42_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__41_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__40_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__39_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__38_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__37_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__36_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__35_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__34_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__33_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__32_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__31_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__30_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__29_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__28_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__27_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__26_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__25_ <= 1'b0;
    end else if(N661) begin
      commit_queue_q_7__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__24_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__23_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__22_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__21_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__20_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__19_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__18_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__17_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__16_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__15_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__14_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__13_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__12_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__11_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__10_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__9_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__8_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__7_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__6_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__5_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__4_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__3_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__2_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__1_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__address__0_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__63_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__62_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__61_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__60_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__59_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__58_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__57_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__56_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__55_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__54_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__53_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__52_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__51_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__50_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__49_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__48_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__47_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__46_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__45_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__44_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__43_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__42_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__41_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__40_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__39_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__38_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__37_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__36_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__35_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__34_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__33_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__32_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__31_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__30_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__29_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__28_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__27_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__26_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__25_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__24_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__23_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__22_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__21_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__20_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__19_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__18_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__17_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__16_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__15_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__14_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__13_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__12_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__11_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__10_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__9_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__8_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__7_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__6_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__5_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__4_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__3_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__2_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__1_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data__0_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__7_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__6_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__5_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__4_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__3_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__2_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__1_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__be__0_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data_size__1_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__data_size__0_ <= 1'b0;
    end else if(N658) begin
      commit_queue_q_7__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_7__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_7__valid_ <= commit_queue_n_7__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__55_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__54_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__53_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__52_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__51_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__50_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__49_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__48_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__47_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__46_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__45_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__44_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__43_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__42_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__41_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__40_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__39_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__38_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__37_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__36_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__35_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__34_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__33_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__32_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__31_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__30_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__29_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__28_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__27_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__26_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__25_ <= 1'b0;
    end else if(N667) begin
      commit_queue_q_6__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__24_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__23_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__22_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__21_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__20_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__19_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__18_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__17_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__16_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__15_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__14_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__13_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__12_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__11_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__10_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__9_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__8_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__7_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__6_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__5_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__4_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__3_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__2_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__1_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__address__0_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__63_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__62_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__61_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__60_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__59_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__58_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__57_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__56_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__55_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__54_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__53_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__52_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__51_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__50_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__49_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__48_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__47_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__46_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__45_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__44_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__43_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__42_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__41_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__40_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__39_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__38_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__37_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__36_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__35_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__34_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__33_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__32_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__31_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__30_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__29_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__28_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__27_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__26_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__25_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__24_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__23_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__22_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__21_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__20_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__19_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__18_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__17_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__16_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__15_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__14_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__13_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__12_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__11_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__10_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__9_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__8_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__7_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__6_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__5_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__4_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__3_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__2_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__1_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data__0_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__7_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__6_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__5_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__4_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__3_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__2_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__1_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__be__0_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data_size__1_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__data_size__0_ <= 1'b0;
    end else if(N664) begin
      commit_queue_q_6__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_6__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_6__valid_ <= commit_queue_n_6__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__55_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__54_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__53_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__52_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__51_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__50_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__49_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__48_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__47_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__46_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__45_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__44_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__43_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__42_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__41_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__40_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__39_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__38_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__37_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__36_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__35_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__34_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__33_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__32_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__31_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__30_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__29_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__28_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__27_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__26_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__25_ <= 1'b0;
    end else if(N673) begin
      commit_queue_q_5__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__24_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__23_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__22_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__21_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__20_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__19_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__18_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__17_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__16_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__15_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__14_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__13_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__12_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__11_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__10_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__9_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__8_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__7_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__6_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__5_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__4_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__3_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__2_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__1_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__address__0_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__63_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__62_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__61_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__60_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__59_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__58_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__57_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__56_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__55_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__54_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__53_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__52_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__51_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__50_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__49_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__48_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__47_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__46_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__45_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__44_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__43_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__42_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__41_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__40_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__39_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__38_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__37_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__36_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__35_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__34_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__33_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__32_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__31_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__30_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__29_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__28_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__27_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__26_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__25_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__24_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__23_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__22_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__21_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__20_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__19_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__18_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__17_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__16_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__15_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__14_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__13_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__12_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__11_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__10_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__9_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__8_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__7_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__6_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__5_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__4_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__3_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__2_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__1_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data__0_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__7_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__6_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__5_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__4_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__3_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__2_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__1_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__be__0_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data_size__1_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__data_size__0_ <= 1'b0;
    end else if(N670) begin
      commit_queue_q_5__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_5__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_5__valid_ <= commit_queue_n_5__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__55_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__54_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__53_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__52_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__51_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__50_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__49_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__48_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__47_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__46_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__45_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__44_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__43_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__42_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__41_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__40_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__39_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__38_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__37_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__36_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__35_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__34_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__33_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__32_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__31_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__30_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__29_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__28_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__27_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__26_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__25_ <= 1'b0;
    end else if(N679) begin
      commit_queue_q_4__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__24_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__23_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__22_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__21_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__20_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__19_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__18_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__17_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__16_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__15_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__14_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__13_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__12_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__11_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__10_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__9_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__8_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__7_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__6_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__5_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__4_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__3_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__2_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__1_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__address__0_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__63_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__62_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__61_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__60_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__59_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__58_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__57_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__56_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__55_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__54_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__53_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__52_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__51_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__50_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__49_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__48_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__47_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__46_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__45_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__44_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__43_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__42_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__41_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__40_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__39_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__38_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__37_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__36_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__35_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__34_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__33_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__32_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__31_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__30_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__29_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__28_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__27_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__26_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__25_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__24_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__23_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__22_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__21_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__20_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__19_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__18_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__17_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__16_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__15_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__14_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__13_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__12_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__11_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__10_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__9_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__8_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__7_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__6_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__5_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__4_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__3_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__2_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__1_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data__0_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__7_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__6_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__5_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__4_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__3_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__2_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__1_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__be__0_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data_size__1_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__data_size__0_ <= 1'b0;
    end else if(N676) begin
      commit_queue_q_4__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_4__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_4__valid_ <= commit_queue_n_4__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__55_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__54_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__53_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__52_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__51_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__50_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__49_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__48_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__47_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__46_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__45_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__44_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__43_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__42_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__41_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__40_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__39_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__38_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__37_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__36_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__35_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__34_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__33_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__32_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__31_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__30_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__29_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__28_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__27_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__26_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__25_ <= 1'b0;
    end else if(N685) begin
      commit_queue_q_3__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__24_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__23_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__22_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__21_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__20_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__19_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__18_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__17_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__16_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__15_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__14_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__13_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__12_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__11_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__10_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__9_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__8_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__7_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__6_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__5_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__4_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__3_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__2_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__1_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__address__0_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__63_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__62_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__61_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__60_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__59_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__58_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__57_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__56_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__55_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__54_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__53_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__52_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__51_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__50_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__49_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__48_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__47_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__46_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__45_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__44_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__43_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__42_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__41_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__40_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__39_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__38_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__37_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__36_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__35_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__34_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__33_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__32_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__31_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__30_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__29_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__28_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__27_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__26_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__25_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__24_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__23_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__22_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__21_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__20_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__19_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__18_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__17_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__16_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__15_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__14_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__13_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__12_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__11_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__10_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__9_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__8_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__7_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__6_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__5_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__4_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__3_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__2_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__1_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data__0_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__7_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__6_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__5_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__4_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__3_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__2_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__1_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__be__0_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data_size__1_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__data_size__0_ <= 1'b0;
    end else if(N682) begin
      commit_queue_q_3__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_3__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_3__valid_ <= commit_queue_n_3__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__55_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__54_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__53_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__52_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__51_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__50_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__49_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__48_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__47_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__46_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__45_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__44_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__43_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__42_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__41_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__40_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__39_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__38_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__37_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__36_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__35_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__34_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__33_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__32_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__31_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__30_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__29_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__28_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__27_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__26_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__25_ <= 1'b0;
    end else if(N691) begin
      commit_queue_q_2__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__24_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__23_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__22_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__21_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__20_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__19_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__18_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__17_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__16_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__15_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__14_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__13_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__12_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__11_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__10_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__9_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__8_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__7_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__6_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__5_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__4_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__3_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__2_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__1_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__address__0_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__63_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__62_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__61_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__60_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__59_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__58_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__57_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__56_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__55_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__54_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__53_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__52_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__51_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__50_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__49_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__48_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__47_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__46_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__45_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__44_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__43_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__42_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__41_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__40_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__39_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__38_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__37_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__36_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__35_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__34_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__33_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__32_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__31_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__30_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__29_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__28_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__27_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__26_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__25_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__24_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__23_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__22_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__21_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__20_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__19_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__18_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__17_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__16_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__15_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__14_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__13_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__12_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__11_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__10_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__9_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__8_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__7_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__6_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__5_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__4_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__3_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__2_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__1_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data__0_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__7_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__6_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__5_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__4_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__3_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__2_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__1_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__be__0_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data_size__1_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__data_size__0_ <= 1'b0;
    end else if(N688) begin
      commit_queue_q_2__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_2__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_2__valid_ <= commit_queue_n_2__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__55_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__54_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__53_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__52_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__51_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__50_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__49_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__48_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__47_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__46_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__45_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__44_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__43_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__42_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__41_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__40_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__39_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__38_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__37_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__36_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__35_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__34_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__33_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__32_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__31_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__30_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__29_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__28_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__27_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__26_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__25_ <= 1'b0;
    end else if(N697) begin
      commit_queue_q_1__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__24_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__23_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__22_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__21_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__20_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__19_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__18_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__17_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__16_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__15_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__14_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__13_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__12_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__11_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__10_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__9_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__8_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__7_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__6_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__5_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__4_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__3_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__2_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__1_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__address__0_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__63_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__62_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__61_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__60_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__59_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__58_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__57_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__56_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__55_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__54_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__53_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__52_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__51_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__50_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__49_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__48_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__47_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__46_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__45_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__44_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__43_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__42_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__41_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__40_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__39_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__38_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__37_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__36_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__35_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__34_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__33_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__32_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__31_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__30_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__29_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__28_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__27_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__26_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__25_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__24_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__23_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__22_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__21_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__20_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__19_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__18_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__17_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__16_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__15_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__14_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__13_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__12_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__11_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__10_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__9_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__8_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__7_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__6_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__5_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__4_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__3_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__2_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__1_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data__0_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__7_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__6_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__5_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__4_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__3_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__2_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__1_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__be__0_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data_size__1_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__data_size__0_ <= 1'b0;
    end else if(N694) begin
      commit_queue_q_1__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_1__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_1__valid_ <= commit_queue_n_1__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__55_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__55_ <= N328;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__54_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__54_ <= N329;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__53_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__53_ <= N330;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__52_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__52_ <= N331;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__51_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__51_ <= N332;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__50_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__50_ <= N333;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__49_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__49_ <= N334;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__48_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__48_ <= N335;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__47_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__47_ <= N336;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__46_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__46_ <= N337;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__45_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__45_ <= N338;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__44_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__44_ <= N339;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__43_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__43_ <= N340;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__42_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__42_ <= N341;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__41_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__41_ <= N342;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__40_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__40_ <= N343;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__39_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__39_ <= N344;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__38_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__38_ <= N345;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__37_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__37_ <= N346;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__36_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__36_ <= N347;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__35_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__35_ <= N348;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__34_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__34_ <= N349;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__33_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__33_ <= N350;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__32_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__32_ <= N351;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__31_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__31_ <= N352;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__30_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__30_ <= N353;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__29_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__29_ <= N354;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__28_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__28_ <= N355;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__27_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__27_ <= N356;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__26_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__26_ <= N357;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__25_ <= 1'b0;
    end else if(N703) begin
      commit_queue_q_0__address__25_ <= N358;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__24_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__24_ <= N359;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__23_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__23_ <= N360;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__22_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__22_ <= N361;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__21_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__21_ <= N362;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__20_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__20_ <= N363;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__19_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__19_ <= N364;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__18_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__18_ <= N365;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__17_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__17_ <= N366;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__16_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__16_ <= N367;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__15_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__15_ <= N368;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__14_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__14_ <= N369;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__13_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__13_ <= N370;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__12_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__12_ <= N371;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__11_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__11_ <= N372;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__10_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__10_ <= N373;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__9_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__9_ <= N374;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__8_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__8_ <= N375;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__7_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__7_ <= N376;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__6_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__6_ <= N377;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__5_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__5_ <= N378;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__4_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__4_ <= N379;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__3_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__3_ <= N380;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__2_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__2_ <= N381;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__1_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__1_ <= N382;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__address__0_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__address__0_ <= N383;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__63_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__63_ <= N384;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__62_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__62_ <= N385;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__61_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__61_ <= N386;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__60_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__60_ <= N387;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__59_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__59_ <= N388;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__58_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__58_ <= N389;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__57_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__57_ <= N390;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__56_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__56_ <= N391;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__55_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__55_ <= N392;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__54_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__54_ <= N393;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__53_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__53_ <= N394;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__52_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__52_ <= N395;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__51_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__51_ <= N396;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__50_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__50_ <= N397;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__49_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__49_ <= N398;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__48_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__48_ <= N399;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__47_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__47_ <= N400;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__46_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__46_ <= N401;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__45_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__45_ <= N402;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__44_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__44_ <= N403;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__43_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__43_ <= N404;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__42_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__42_ <= N405;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__41_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__41_ <= N406;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__40_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__40_ <= N407;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__39_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__39_ <= N408;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__38_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__38_ <= N409;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__37_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__37_ <= N410;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__36_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__36_ <= N411;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__35_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__35_ <= N412;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__34_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__34_ <= N413;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__33_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__33_ <= N414;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__32_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__32_ <= N415;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__31_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__31_ <= N416;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__30_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__30_ <= N417;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__29_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__29_ <= N418;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__28_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__28_ <= N419;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__27_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__27_ <= N420;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__26_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__26_ <= N421;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__25_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__25_ <= N422;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__24_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__24_ <= N423;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__23_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__23_ <= N424;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__22_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__22_ <= N425;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__21_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__21_ <= N426;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__20_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__20_ <= N427;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__19_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__19_ <= N428;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__18_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__18_ <= N429;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__17_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__17_ <= N430;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__16_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__16_ <= N431;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__15_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__15_ <= N432;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__14_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__14_ <= N433;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__13_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__13_ <= N434;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__12_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__12_ <= N435;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__11_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__11_ <= N436;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__10_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__10_ <= N437;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__9_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__9_ <= N438;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__8_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__8_ <= N439;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__7_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__7_ <= N440;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__6_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__6_ <= N441;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__5_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__5_ <= N442;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__4_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__4_ <= N443;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__3_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__3_ <= N444;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__2_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__2_ <= N445;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__1_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__1_ <= N446;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data__0_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data__0_ <= N447;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__7_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__7_ <= N448;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__6_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__6_ <= N449;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__5_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__5_ <= N450;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__4_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__4_ <= N451;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__3_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__3_ <= N452;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__2_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__2_ <= N453;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__1_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__1_ <= N454;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__be__0_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__be__0_ <= N455;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data_size__1_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data_size__1_ <= N456;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__data_size__0_ <= 1'b0;
    end else if(N700) begin
      commit_queue_q_0__data_size__0_ <= N457;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_queue_q_0__valid_ <= 1'b0;
    end else if(1'b1) begin
      commit_queue_q_0__valid_ <= commit_queue_n_0__valid_;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_read_pointer_q[2] <= 1'b0;
    end else if(N706) begin
      commit_read_pointer_q[2] <= N301;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_read_pointer_q[1] <= 1'b0;
    end else if(N706) begin
      commit_read_pointer_q[1] <= N300;
    end 
  end


  always @(posedge clk_i or posedge N605) begin
    if(N605) begin
      commit_read_pointer_q[0] <= 1'b0;
    end else if(N706) begin
      commit_read_pointer_q[0] <= N299;
    end 
  end

  assign N707 = commit_status_cnt_q[2] | commit_status_cnt_q[3];
  assign N708 = commit_status_cnt_q[1] | N707;
  assign N709 = commit_status_cnt_q[0] | N708;
  assign no_st_pending_o = ~N709;
  assign { N485, N484, N483 } = commit_write_pointer_q + 1'b1;
  assign { N186, N185 } = speculative_read_pointer_q + 1'b1;
  assign { N160, N159 } = speculative_write_pointer_q + 1'b1;
  assign { N163, N162, N161 } = speculative_status_cnt_q + 1'b1;
  assign { N193, N192, N191 } = { N170, N169, N168 } - commit_i;
  assign { N301, N300, N299 } = commit_read_pointer_q + 1'b1;
  assign { N313, N312, N311, N310 } = commit_status_cnt_q - N727;
  assign { N489, N488, N487, N486 } = { N313, N312, N311, N310 } + 1'b1;
  assign N118 = speculative_write_pointer_q[0] & speculative_write_pointer_q[1];
  assign N117 = N0 & speculative_write_pointer_q[1];
  assign N0 = ~speculative_write_pointer_q[0];
  assign N116 = speculative_write_pointer_q[0] & N1;
  assign N1 = ~speculative_write_pointer_q[1];
  assign N115 = N2 & N3;
  assign N2 = ~speculative_write_pointer_q[0];
  assign N3 = ~speculative_write_pointer_q[1];
  assign N126 = speculative_write_pointer_q[0] & speculative_write_pointer_q[1];
  assign N125 = N4 & speculative_write_pointer_q[1];
  assign N4 = ~speculative_write_pointer_q[0];
  assign N124 = speculative_write_pointer_q[0] & N5;
  assign N5 = ~speculative_write_pointer_q[1];
  assign N123 = N6 & N7;
  assign N6 = ~speculative_write_pointer_q[0];
  assign N7 = ~speculative_write_pointer_q[1];
  assign N134 = speculative_write_pointer_q[0] & speculative_write_pointer_q[1];
  assign N133 = N8 & speculative_write_pointer_q[1];
  assign N8 = ~speculative_write_pointer_q[0];
  assign N132 = speculative_write_pointer_q[0] & N9;
  assign N9 = ~speculative_write_pointer_q[1];
  assign N131 = N10 & N11;
  assign N10 = ~speculative_write_pointer_q[0];
  assign N11 = ~speculative_write_pointer_q[1];
  assign N142 = speculative_write_pointer_q[0] & speculative_write_pointer_q[1];
  assign N141 = N12 & speculative_write_pointer_q[1];
  assign N12 = ~speculative_write_pointer_q[0];
  assign N140 = speculative_write_pointer_q[0] & N13;
  assign N13 = ~speculative_write_pointer_q[1];
  assign N139 = N14 & N15;
  assign N14 = ~speculative_write_pointer_q[0];
  assign N15 = ~speculative_write_pointer_q[1];
  assign N150 = speculative_write_pointer_q[0] & speculative_write_pointer_q[1];
  assign N149 = N16 & speculative_write_pointer_q[1];
  assign N16 = ~speculative_write_pointer_q[0];
  assign N148 = speculative_write_pointer_q[0] & N17;
  assign N17 = ~speculative_write_pointer_q[1];
  assign N147 = N18 & N19;
  assign N18 = ~speculative_write_pointer_q[0];
  assign N19 = ~speculative_write_pointer_q[1];
  assign N176 = speculative_read_pointer_q[0] & speculative_read_pointer_q[1];
  assign N175 = N20 & speculative_read_pointer_q[1];
  assign N20 = ~speculative_read_pointer_q[0];
  assign N174 = speculative_read_pointer_q[0] & N21;
  assign N21 = ~speculative_read_pointer_q[1];
  assign N173 = N22 & N23;
  assign N22 = ~speculative_read_pointer_q[0];
  assign N23 = ~speculative_read_pointer_q[1];
  assign N711 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N282 = N711 & commit_read_pointer_q[2];
  assign N712 = N24 & commit_read_pointer_q[1];
  assign N24 = ~commit_read_pointer_q[0];
  assign N281 = N712 & commit_read_pointer_q[2];
  assign N713 = commit_read_pointer_q[0] & N25;
  assign N25 = ~commit_read_pointer_q[1];
  assign N280 = N713 & commit_read_pointer_q[2];
  assign N714 = N26 & N27;
  assign N26 = ~commit_read_pointer_q[0];
  assign N27 = ~commit_read_pointer_q[1];
  assign N279 = N714 & commit_read_pointer_q[2];
  assign N715 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N278 = N715 & N28;
  assign N28 = ~commit_read_pointer_q[2];
  assign N716 = N29 & commit_read_pointer_q[1];
  assign N29 = ~commit_read_pointer_q[0];
  assign N277 = N716 & N30;
  assign N30 = ~commit_read_pointer_q[2];
  assign N717 = commit_read_pointer_q[0] & N31;
  assign N31 = ~commit_read_pointer_q[1];
  assign N276 = N717 & N32;
  assign N32 = ~commit_read_pointer_q[2];
  assign N718 = N33 & N34;
  assign N33 = ~commit_read_pointer_q[0];
  assign N34 = ~commit_read_pointer_q[1];
  assign N275 = N718 & N35;
  assign N35 = ~commit_read_pointer_q[2];
  assign N719 = commit_write_pointer_q[0] & commit_write_pointer_q[1];
  assign N466 = N719 & commit_write_pointer_q[2];
  assign N720 = N36 & commit_write_pointer_q[1];
  assign N36 = ~commit_write_pointer_q[0];
  assign N465 = N720 & commit_write_pointer_q[2];
  assign N721 = commit_write_pointer_q[0] & N37;
  assign N37 = ~commit_write_pointer_q[1];
  assign N464 = N721 & commit_write_pointer_q[2];
  assign N722 = N38 & N39;
  assign N38 = ~commit_write_pointer_q[0];
  assign N39 = ~commit_write_pointer_q[1];
  assign N463 = N722 & commit_write_pointer_q[2];
  assign N723 = commit_write_pointer_q[0] & commit_write_pointer_q[1];
  assign N462 = N723 & N40;
  assign N40 = ~commit_write_pointer_q[2];
  assign N724 = N41 & commit_write_pointer_q[1];
  assign N41 = ~commit_write_pointer_q[0];
  assign N461 = N724 & N42;
  assign N42 = ~commit_write_pointer_q[2];
  assign N725 = commit_write_pointer_q[0] & N43;
  assign N43 = ~commit_write_pointer_q[1];
  assign N460 = N725 & N44;
  assign N44 = ~commit_write_pointer_q[2];
  assign N726 = N45 & N46;
  assign N45 = ~commit_write_pointer_q[0];
  assign N46 = ~commit_write_pointer_q[1];
  assign N459 = N726 & N47;
  assign N47 = ~commit_write_pointer_q[2];
  assign N152 = (N48)? 1'b1 : 
                (N151)? speculative_queue_q_0__valid_ : 1'b0;
  assign N48 = N147;
  assign N154 = (N49)? 1'b1 : 
                (N153)? speculative_queue_q_1__valid_ : 1'b0;
  assign N49 = N148;
  assign N156 = (N50)? 1'b1 : 
                (N155)? speculative_queue_q_2__valid_ : 1'b0;
  assign N50 = N149;
  assign N158 = (N51)? 1'b1 : 
                (N157)? speculative_queue_q_3__valid_ : 1'b0;
  assign N51 = N150;
  assign { N167, N166, N165, N164 } = (N52)? { N158, N156, N154, N152 } : 
                                      (N53)? { speculative_queue_q_3__valid_, speculative_queue_q_2__valid_, speculative_queue_q_1__valid_, speculative_queue_q_0__valid_ } : 1'b0;
  assign N52 = valid_i;
  assign N53 = N114;
  assign { N170, N169, N168 } = (N52)? { N163, N162, N161 } : 
                                (N53)? speculative_status_cnt_q : 1'b0;
  assign N178 = (N54)? 1'b0 : 
                (N177)? N164 : 1'b0;
  assign N54 = N173;
  assign N180 = (N55)? 1'b0 : 
                (N179)? N165 : 1'b0;
  assign N55 = N174;
  assign N182 = (N56)? 1'b0 : 
                (N181)? N166 : 1'b0;
  assign N56 = N175;
  assign N184 = (N57)? 1'b0 : 
                (N183)? N167 : 1'b0;
  assign N57 = N176;
  assign { N190, N189, N188, N187 } = (N58)? { N184, N182, N180, N178 } : 
                                      (N59)? { N167, N166, N165, N164 } : 1'b0;
  assign N58 = commit_i;
  assign N59 = N171;
  assign { speculative_queue_n_3__valid_, speculative_queue_n_2__valid_, speculative_queue_n_1__valid_, speculative_queue_n_0__valid_ } = (N60)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                          (N61)? { N190, N189, N188, N187 } : 1'b0;
  assign N60 = flush_i;
  assign N61 = N194;
  assign speculative_write_pointer_n = (N60)? speculative_read_pointer_q : 
                                       (N61)? { N160, N159 } : 1'b0;
  assign speculative_status_cnt_n = (N60)? { 1'b0, 1'b0, 1'b0 } : 
                                    (N61)? { N193, N192, N191 } : 1'b0;
  assign N284 = (N62)? 1'b0 : 
                (N283)? commit_queue_q_0__valid_ : 1'b0;
  assign N62 = N275;
  assign N286 = (N63)? 1'b0 : 
                (N285)? commit_queue_q_1__valid_ : 1'b0;
  assign N63 = N276;
  assign N288 = (N64)? 1'b0 : 
                (N287)? commit_queue_q_2__valid_ : 1'b0;
  assign N64 = N277;
  assign N290 = (N65)? 1'b0 : 
                (N289)? commit_queue_q_3__valid_ : 1'b0;
  assign N65 = N278;
  assign N292 = (N66)? 1'b0 : 
                (N291)? commit_queue_q_4__valid_ : 1'b0;
  assign N66 = N279;
  assign N294 = (N67)? 1'b0 : 
                (N293)? commit_queue_q_5__valid_ : 1'b0;
  assign N67 = N280;
  assign N296 = (N68)? 1'b0 : 
                (N295)? commit_queue_q_6__valid_ : 1'b0;
  assign N68 = N281;
  assign N298 = (N69)? 1'b0 : 
                (N297)? commit_queue_q_7__valid_ : 1'b0;
  assign N69 = N282;
  assign { N309, N308, N307, N306, N305, N304, N303, N302 } = (N70)? { N298, N296, N294, N292, N290, N288, N286, N284 } : 
                                                              (N273)? { commit_queue_q_7__valid_, commit_queue_q_6__valid_, commit_queue_q_5__valid_, commit_queue_q_4__valid_, commit_queue_q_3__valid_, commit_queue_q_2__valid_, commit_queue_q_1__valid_, commit_queue_q_0__valid_ } : 1'b0;
  assign N70 = req_port_i[65];
  assign { N321, N320, N319, N318, N317, N316, N315, N314 } = (N71)? { N309, N308, N307, N306, N305, N304, N303, N302 } : 
                                                              (N271)? { commit_queue_q_7__valid_, commit_queue_q_6__valid_, commit_queue_q_5__valid_, commit_queue_q_4__valid_, commit_queue_q_3__valid_, commit_queue_q_2__valid_, commit_queue_q_1__valid_, commit_queue_q_0__valid_ } : 1'b0;
  assign N71 = req_port_o[13];
  assign N468 = (N72)? N458 : 
                (N467)? N314 : 1'b0;
  assign N72 = N459;
  assign N470 = (N73)? N458 : 
                (N469)? N315 : 1'b0;
  assign N73 = N460;
  assign N472 = (N74)? N458 : 
                (N471)? N316 : 1'b0;
  assign N74 = N461;
  assign N474 = (N75)? N458 : 
                (N473)? N317 : 1'b0;
  assign N75 = N462;
  assign N476 = (N76)? N458 : 
                (N475)? N318 : 1'b0;
  assign N76 = N463;
  assign N478 = (N77)? N458 : 
                (N477)? N319 : 1'b0;
  assign N77 = N464;
  assign N480 = (N78)? N458 : 
                (N479)? N320 : 1'b0;
  assign N78 = N465;
  assign N482 = (N79)? N458 : 
                (N481)? N321 : 1'b0;
  assign N79 = N466;
  assign { commit_queue_n_7__valid_, commit_queue_n_6__valid_, commit_queue_n_5__valid_, commit_queue_n_4__valid_, commit_queue_n_3__valid_, commit_queue_n_2__valid_, commit_queue_n_1__valid_, commit_queue_n_0__valid_ } = (N58)? { N482, N480, N478, N476, N474, N472, N470, N468 } : 
                                                                                                                                                                                                                              (N59)? { N321, N320, N319, N318, N317, N316, N315, N314 } : 1'b0;
  assign commit_status_cnt_n = (N58)? { N489, N488, N487, N486 } : 
                               (N59)? { N313, N312, N311, N310 } : 1'b0;
  assign N492 = ~N491;
  assign N499 = (N80)? 1'b1 : 
                (N498)? N491 : 1'b0;
  assign N80 = N497;
  assign N500 = (N80)? 1'b0 : 
                (N498)? N492 : 1'b0;
  assign N507 = (N81)? 1'b1 : 
                (N506)? N499 : 1'b0;
  assign N81 = N505;
  assign N508 = (N81)? 1'b0 : 
                (N506)? N500 : 1'b0;
  assign N515 = (N82)? 1'b1 : 
                (N514)? N507 : 1'b0;
  assign N82 = N513;
  assign N516 = (N82)? 1'b0 : 
                (N514)? N508 : 1'b0;
  assign N523 = (N83)? 1'b1 : 
                (N522)? N515 : 1'b0;
  assign N83 = N521;
  assign N524 = (N83)? 1'b0 : 
                (N522)? N516 : 1'b0;
  assign N531 = (N84)? 1'b1 : 
                (N530)? N523 : 1'b0;
  assign N84 = N529;
  assign N532 = (N84)? 1'b0 : 
                (N530)? N524 : 1'b0;
  assign N539 = (N85)? 1'b1 : 
                (N538)? N531 : 1'b0;
  assign N85 = N537;
  assign N540 = (N85)? 1'b0 : 
                (N538)? N532 : 1'b0;
  assign N546 = (N86)? 1'b1 : 
                (N545)? N539 : 1'b0;
  assign N86 = N544;
  assign N548 = (N87)? N546 : 
                (N547)? N539 : 1'b0;
  assign N87 = N540;
  assign N549 = (N87)? N548 : 
                (N88)? N539 : 1'b0;
  assign N88 = N541;
  assign N551 = (N89)? N549 : 
                (N550)? N531 : 1'b0;
  assign N89 = N532;
  assign N552 = (N89)? N551 : 
                (N90)? N531 : 1'b0;
  assign N90 = N533;
  assign N554 = (N91)? N552 : 
                (N553)? N523 : 1'b0;
  assign N91 = N524;
  assign N555 = (N91)? N554 : 
                (N92)? N523 : 1'b0;
  assign N92 = N525;
  assign N557 = (N93)? N555 : 
                (N556)? N515 : 1'b0;
  assign N93 = N516;
  assign N558 = (N93)? N557 : 
                (N94)? N515 : 1'b0;
  assign N94 = N517;
  assign N560 = (N95)? N558 : 
                (N559)? N507 : 1'b0;
  assign N95 = N508;
  assign N561 = (N95)? N560 : 
                (N96)? N507 : 1'b0;
  assign N96 = N509;
  assign N563 = (N97)? N561 : 
                (N562)? N499 : 1'b0;
  assign N97 = N500;
  assign N564 = (N97)? N563 : 
                (N98)? N499 : 1'b0;
  assign N98 = N501;
  assign N565 = (N99)? N564 : 
                (N100)? N491 : 1'b0;
  assign N99 = N494;
  assign N100 = N491;
  assign N566 = (N101)? N565 : 
                (N100)? N491 : 1'b0;
  assign N101 = N492;
  assign N570 = (N102)? 1'b1 : 
                (N569)? N566 : 1'b0;
  assign N102 = N568;
  assign N571 = ~N568;
  assign N578 = (N103)? 1'b1 : 
                (N577)? N570 : 1'b0;
  assign N103 = N576;
  assign N579 = (N103)? 1'b0 : 
                (N577)? N571 : 1'b0;
  assign N586 = (N104)? 1'b1 : 
                (N585)? N578 : 1'b0;
  assign N104 = N584;
  assign N587 = (N104)? 1'b0 : 
                (N585)? N579 : 1'b0;
  assign N593 = (N105)? 1'b1 : 
                (N592)? N586 : 1'b0;
  assign N105 = N591;
  assign N595 = (N106)? N593 : 
                (N594)? N586 : 1'b0;
  assign N106 = N587;
  assign N596 = (N106)? N595 : 
                (N107)? N586 : 1'b0;
  assign N107 = N588;
  assign N598 = (N108)? N596 : 
                (N597)? N578 : 1'b0;
  assign N108 = N579;
  assign N599 = (N108)? N598 : 
                (N109)? N578 : 1'b0;
  assign N109 = N580;
  assign N600 = (N110)? N599 : 
                (N102)? N570 : 1'b0;
  assign N110 = N573;
  assign N601 = (N111)? N600 : 
                (N102)? N570 : 1'b0;
  assign N111 = N571;
  assign page_offset_matches_o = (N112)? 1'b1 : 
                                 (N604)? N601 : 1'b0;
  assign N112 = N603;
  assign ready_o = N113 | commit_i;
  assign N114 = ~valid_i;
  assign N119 = ~N115;
  assign N120 = ~N116;
  assign N121 = ~N117;
  assign N122 = ~N118;
  assign N127 = ~N123;
  assign N128 = ~N124;
  assign N129 = ~N125;
  assign N130 = ~N126;
  assign N135 = ~N131;
  assign N136 = ~N132;
  assign N137 = ~N133;
  assign N138 = ~N134;
  assign N143 = ~N139;
  assign N144 = ~N140;
  assign N145 = ~N141;
  assign N146 = ~N142;
  assign N151 = ~N147;
  assign N153 = ~N148;
  assign N155 = ~N149;
  assign N157 = ~N150;
  assign N171 = ~commit_i;
  assign N172 = commit_i;
  assign N177 = ~N173;
  assign N179 = ~N174;
  assign N181 = ~N175;
  assign N183 = ~N176;
  assign N194 = ~flush_i;
  assign N195 = ~commit_read_pointer_q[0];
  assign N196 = ~commit_read_pointer_q[1];
  assign N197 = N195 & N196;
  assign N198 = N195 & commit_read_pointer_q[1];
  assign N199 = commit_read_pointer_q[0] & N196;
  assign N200 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N201 = ~commit_read_pointer_q[2];
  assign N202 = N197 & N201;
  assign N203 = N197 & commit_read_pointer_q[2];
  assign N204 = N199 & N201;
  assign N205 = N199 & commit_read_pointer_q[2];
  assign N206 = N198 & N201;
  assign N207 = N198 & commit_read_pointer_q[2];
  assign N208 = N200 & N201;
  assign N209 = N200 & commit_read_pointer_q[2];
  assign N210 = N195 & N196;
  assign N211 = N195 & commit_read_pointer_q[1];
  assign N212 = commit_read_pointer_q[0] & N196;
  assign N213 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N214 = N210 & N201;
  assign N215 = N210 & commit_read_pointer_q[2];
  assign N216 = N212 & N201;
  assign N217 = N212 & commit_read_pointer_q[2];
  assign N218 = N211 & N201;
  assign N219 = N211 & commit_read_pointer_q[2];
  assign N220 = N213 & N201;
  assign N221 = N213 & commit_read_pointer_q[2];
  assign N222 = N195 & N196;
  assign N223 = N195 & commit_read_pointer_q[1];
  assign N224 = commit_read_pointer_q[0] & N196;
  assign N225 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N226 = N222 & N201;
  assign N227 = N222 & commit_read_pointer_q[2];
  assign N228 = N224 & N201;
  assign N229 = N224 & commit_read_pointer_q[2];
  assign N230 = N223 & N201;
  assign N231 = N223 & commit_read_pointer_q[2];
  assign N232 = N225 & N201;
  assign N233 = N225 & commit_read_pointer_q[2];
  assign N234 = N195 & N196;
  assign N235 = N195 & commit_read_pointer_q[1];
  assign N236 = commit_read_pointer_q[0] & N196;
  assign N237 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N238 = N234 & N201;
  assign N239 = N234 & commit_read_pointer_q[2];
  assign N240 = N236 & N201;
  assign N241 = N236 & commit_read_pointer_q[2];
  assign N242 = N235 & N201;
  assign N243 = N235 & commit_read_pointer_q[2];
  assign N244 = N237 & N201;
  assign N245 = N237 & commit_read_pointer_q[2];
  assign N246 = N195 & N196;
  assign N247 = N195 & commit_read_pointer_q[1];
  assign N248 = commit_read_pointer_q[0] & N196;
  assign N249 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N250 = N246 & N201;
  assign N251 = N246 & commit_read_pointer_q[2];
  assign N252 = N248 & N201;
  assign N253 = N248 & commit_read_pointer_q[2];
  assign N254 = N247 & N201;
  assign N255 = N247 & commit_read_pointer_q[2];
  assign N256 = N249 & N201;
  assign N257 = N249 & commit_read_pointer_q[2];
  assign commit_ready_o = ~commit_status_cnt_q[3];
  assign N258 = N195 & N196;
  assign N259 = N195 & commit_read_pointer_q[1];
  assign N260 = commit_read_pointer_q[0] & N196;
  assign N261 = commit_read_pointer_q[0] & commit_read_pointer_q[1];
  assign N262 = N258 & N201;
  assign N263 = N258 & commit_read_pointer_q[2];
  assign N264 = N260 & N201;
  assign N265 = N260 & commit_read_pointer_q[2];
  assign N266 = N259 & N201;
  assign N267 = N259 & commit_read_pointer_q[2];
  assign N268 = N261 & N201;
  assign N269 = N261 & commit_read_pointer_q[2];
  assign req_port_o[13] = N270;
  assign N271 = ~req_port_o[13];
  assign N272 = req_port_o[13];
  assign N273 = ~req_port_i[65];
  assign N274 = N272 & req_port_i[65];
  assign N283 = ~N275;
  assign N285 = ~N276;
  assign N287 = ~N277;
  assign N289 = ~N278;
  assign N291 = ~N279;
  assign N293 = ~N280;
  assign N295 = ~N281;
  assign N297 = ~N282;
  assign N322 = ~speculative_read_pointer_q[0];
  assign N323 = ~speculative_read_pointer_q[1];
  assign N324 = N322 & N323;
  assign N325 = N322 & speculative_read_pointer_q[1];
  assign N326 = speculative_read_pointer_q[0] & N323;
  assign N327 = speculative_read_pointer_q[0] & speculative_read_pointer_q[1];
  assign N467 = ~N459;
  assign N469 = ~N460;
  assign N471 = ~N461;
  assign N473 = ~N462;
  assign N475 = ~N463;
  assign N477 = ~N464;
  assign N479 = ~N465;
  assign N481 = ~N466;
  assign N491 = N490 & commit_queue_q_0__valid_;
  assign N493 = N492;
  assign N494 = ~N491;
  assign N495 = N493 & N494;
  assign N497 = N496 & commit_queue_q_1__valid_;
  assign N498 = ~N497;
  assign N501 = ~N500;
  assign N502 = N495 & N500;
  assign N503 = N502 & N500;
  assign N505 = N504 & commit_queue_q_2__valid_;
  assign N506 = ~N505;
  assign N509 = ~N508;
  assign N510 = N503 & N508;
  assign N511 = N510 & N508;
  assign N513 = N512 & commit_queue_q_3__valid_;
  assign N514 = ~N513;
  assign N517 = ~N516;
  assign N518 = N511 & N516;
  assign N519 = N518 & N516;
  assign N521 = N520 & commit_queue_q_4__valid_;
  assign N522 = ~N521;
  assign N525 = ~N524;
  assign N526 = N519 & N524;
  assign N527 = N526 & N524;
  assign N529 = N528 & commit_queue_q_5__valid_;
  assign N530 = ~N529;
  assign N533 = ~N532;
  assign N534 = N527 & N532;
  assign N535 = N534 & N532;
  assign N537 = N536 & commit_queue_q_6__valid_;
  assign N538 = ~N537;
  assign N541 = ~N540;
  assign N542 = N535 & N540;
  assign N544 = N543 & commit_queue_q_7__valid_;
  assign N545 = ~N544;
  assign N547 = ~N540;
  assign N550 = ~N532;
  assign N553 = ~N524;
  assign N556 = ~N516;
  assign N559 = ~N508;
  assign N562 = ~N500;
  assign N568 = N567 & speculative_queue_q_0__valid_;
  assign N569 = ~N568;
  assign N572 = N571;
  assign N573 = ~N568;
  assign N574 = N572 & N573;
  assign N576 = N575 & speculative_queue_q_1__valid_;
  assign N577 = ~N576;
  assign N580 = ~N579;
  assign N581 = N574 & N579;
  assign N582 = N581 & N579;
  assign N584 = N583 & speculative_queue_q_2__valid_;
  assign N585 = ~N584;
  assign N588 = ~N587;
  assign N589 = N582 & N587;
  assign N591 = N590 & speculative_queue_q_3__valid_;
  assign N592 = ~N591;
  assign N594 = ~N587;
  assign N597 = ~N579;
  assign N603 = N602 & valid_without_flush_i;
  assign N604 = ~N603;
  assign N605 = ~rst_ni;
  assign N606 = N114 & N194;
  assign N607 = ~N606;
  assign N608 = N122 & valid_i;
  assign N609 = N608 | N114;
  assign N610 = ~N609;
  assign N611 = N130 & valid_i;
  assign N612 = N611 | N114;
  assign N613 = ~N612;
  assign N614 = N138 & valid_i;
  assign N615 = N614 | N114;
  assign N616 = ~N615;
  assign N617 = N146 & valid_i;
  assign N618 = N617 | N114;
  assign N619 = ~N618;
  assign N620 = N121 & valid_i;
  assign N621 = N620 | N114;
  assign N622 = ~N621;
  assign N623 = N129 & valid_i;
  assign N624 = N623 | N114;
  assign N625 = ~N624;
  assign N626 = N137 & valid_i;
  assign N627 = N626 | N114;
  assign N628 = ~N627;
  assign N629 = N145 & valid_i;
  assign N630 = N629 | N114;
  assign N631 = ~N630;
  assign N632 = N120 & valid_i;
  assign N633 = N632 | N114;
  assign N634 = ~N633;
  assign N635 = N128 & valid_i;
  assign N636 = N635 | N114;
  assign N637 = ~N636;
  assign N638 = N136 & valid_i;
  assign N639 = N638 | N114;
  assign N640 = ~N639;
  assign N641 = N144 & valid_i;
  assign N642 = N641 | N114;
  assign N643 = ~N642;
  assign N644 = N119 & valid_i;
  assign N645 = N644 | N114;
  assign N646 = ~N645;
  assign N647 = N127 & valid_i;
  assign N648 = N647 | N114;
  assign N649 = ~N648;
  assign N650 = N135 & valid_i;
  assign N651 = N650 | N114;
  assign N652 = ~N651;
  assign N653 = N143 & valid_i;
  assign N654 = N653 | N114;
  assign N655 = ~N654;
  assign N656 = N481 & commit_i;
  assign N657 = N656 | N171;
  assign N658 = ~N657;
  assign N659 = N481 & commit_i;
  assign N660 = N659 | N171;
  assign N661 = ~N660;
  assign N662 = N479 & commit_i;
  assign N663 = N662 | N171;
  assign N664 = ~N663;
  assign N665 = N479 & commit_i;
  assign N666 = N665 | N171;
  assign N667 = ~N666;
  assign N668 = N477 & commit_i;
  assign N669 = N668 | N171;
  assign N670 = ~N669;
  assign N671 = N477 & commit_i;
  assign N672 = N671 | N171;
  assign N673 = ~N672;
  assign N674 = N475 & commit_i;
  assign N675 = N674 | N171;
  assign N676 = ~N675;
  assign N677 = N475 & commit_i;
  assign N678 = N677 | N171;
  assign N679 = ~N678;
  assign N680 = N473 & commit_i;
  assign N681 = N680 | N171;
  assign N682 = ~N681;
  assign N683 = N473 & commit_i;
  assign N684 = N683 | N171;
  assign N685 = ~N684;
  assign N686 = N471 & commit_i;
  assign N687 = N686 | N171;
  assign N688 = ~N687;
  assign N689 = N471 & commit_i;
  assign N690 = N689 | N171;
  assign N691 = ~N690;
  assign N692 = N469 & commit_i;
  assign N693 = N692 | N171;
  assign N694 = ~N693;
  assign N695 = N469 & commit_i;
  assign N696 = N695 | N171;
  assign N697 = ~N696;
  assign N698 = N467 & commit_i;
  assign N699 = N698 | N171;
  assign N700 = ~N699;
  assign N701 = N467 & commit_i;
  assign N702 = N701 | N171;
  assign N703 = ~N702;
  assign N704 = N273 & req_port_o[13];
  assign N705 = N704 | N271;
  assign N706 = ~N705;
  assign N727 = req_port_i[65] & req_port_o[13];
  assign N728 = N273 | N271;

endmodule