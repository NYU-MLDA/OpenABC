module DCacheModuleanon2( // @[:freechips.rocketchip.system.TinyConfig.fir@102989.2]
  input         io_in_2_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  input  [31:0] io_in_2_bits_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  input         io_in_3_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  input  [31:0] io_in_3_bits_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  output        io_in_5_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  input         io_in_5_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  output        io_in_7_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  input         io_in_7_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  input  [31:0] io_in_7_bits_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  output        io_out_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  output        io_out_bits_write, // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
  output [31:0] io_out_bits_addr // @[:freechips.rocketchip.system.TinyConfig.fir@102992.4]
);
  wire [31:0] _GEN_22; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103024.4]
  wire  _T_2; // @[Arbiter.scala 31:68:freechips.rocketchip.system.TinyConfig.fir@103058.4]
  wire  _T_9; // @[Arbiter.scala 31:78:freechips.rocketchip.system.TinyConfig.fir@103065.4]
  wire  _T_21; // @[Arbiter.scala 135:19:freechips.rocketchip.system.TinyConfig.fir@103085.4]
  assign _GEN_22 = io_in_3_valid ? io_in_3_bits_addr : io_in_7_bits_addr; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103024.4]
  assign _T_2 = io_in_2_valid | io_in_3_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.TinyConfig.fir@103058.4]
  assign _T_9 = _T_2 == 1'h0; // @[Arbiter.scala 31:78:freechips.rocketchip.system.TinyConfig.fir@103065.4]
  assign _T_21 = _T_9 == 1'h0; // @[Arbiter.scala 135:19:freechips.rocketchip.system.TinyConfig.fir@103085.4]
  assign io_in_5_ready = _T_2 == 1'h0; // @[Arbiter.scala 134:14:freechips.rocketchip.system.TinyConfig.fir@103080.4]
  assign io_in_7_ready = _T_2 == 1'h0; // @[Arbiter.scala 134:14:freechips.rocketchip.system.TinyConfig.fir@103084.4]
  assign io_out_valid = _T_21 | io_in_7_valid; // @[Arbiter.scala 135:16:freechips.rocketchip.system.TinyConfig.fir@103087.4]
  assign io_out_bits_write = io_in_2_valid ? 1'h1 : io_in_3_valid; // @[Arbiter.scala 124:15:freechips.rocketchip.system.TinyConfig.fir@102999.4 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103006.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103014.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103022.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103030.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103038.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103046.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103054.6]
  assign io_out_bits_addr = io_in_2_valid ? io_in_2_bits_addr : _GEN_22; // @[Arbiter.scala 124:15:freechips.rocketchip.system.TinyConfig.fir@102998.4 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103005.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103013.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103021.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103029.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103037.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103045.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103053.6]
endmodule