module CSRFile
(
  clk,
  reset,
  io_host_reset,
  io_host_id,
  io_host_csr_req_ready,
  io_host_csr_req_valid,
  io_host_csr_req_bits_rw,
  io_host_csr_req_bits_addr,
  io_host_csr_req_bits_data,
  io_host_csr_resp_ready,
  io_host_csr_resp_valid,
  io_host_csr_resp_bits,
  io_host_debug_stats_csr,
  io_rw_addr,
  io_rw_cmd,
  io_rw_rdata,
  io_rw_wdata,
  io_csr_stall,
  io_csr_xcpt,
  io_eret,
  io_status_sd,
  io_status_zero2,
  io_status_sd_rv32,
  io_status_zero1,
  io_status_vm,
  io_status_mprv,
  io_status_xs,
  io_status_fs,
  io_status_prv3,
  io_status_ie3,
  io_status_prv2,
  io_status_ie2,
  io_status_prv1,
  io_status_ie1,
  io_status_prv,
  io_status_ie,
  io_ptbr,
  io_evec,
  io_exception,
  io_retire,
  io_uarch_counters_15,
  io_uarch_counters_14,
  io_uarch_counters_13,
  io_uarch_counters_12,
  io_uarch_counters_11,
  io_uarch_counters_10,
  io_uarch_counters_9,
  io_uarch_counters_8,
  io_uarch_counters_7,
  io_uarch_counters_6,
  io_uarch_counters_5,
  io_uarch_counters_4,
  io_uarch_counters_3,
  io_uarch_counters_2,
  io_uarch_counters_1,
  io_uarch_counters_0,
  io_cause,
  io_pc,
  io_fatc,
  io_time,
  io_fcsr_rm,
  io_fcsr_flags_valid,
  io_fcsr_flags_bits,
  io_rocc_cmd_ready,
  io_rocc_resp_valid,
  io_rocc_resp_bits_rd,
  io_rocc_resp_bits_data,
  io_rocc_mem_req_valid,
  io_rocc_mem_req_bits_addr,
  io_rocc_mem_req_bits_tag,
  io_rocc_mem_req_bits_cmd,
  io_rocc_mem_req_bits_typ,
  io_rocc_mem_req_bits_kill,
  io_rocc_mem_req_bits_phys,
  io_rocc_mem_req_bits_data,
  io_rocc_mem_invalidate_lr,
  io_rocc_busy,
  io_rocc_interrupt,
  io_rocc_autl_acquire_valid,
  io_rocc_autl_acquire_bits_addr_block,
  io_rocc_autl_acquire_bits_client_xact_id,
  io_rocc_autl_acquire_bits_addr_beat,
  io_rocc_autl_acquire_bits_is_builtin_type,
  io_rocc_autl_acquire_bits_a_type,
  io_rocc_autl_acquire_bits_union,
  io_rocc_autl_acquire_bits_data,
  io_rocc_autl_grant_ready,
  io_rocc_fpu_req_valid,
  io_rocc_fpu_req_bits_cmd,
  io_rocc_fpu_req_bits_ldst,
  io_rocc_fpu_req_bits_wen,
  io_rocc_fpu_req_bits_ren1,
  io_rocc_fpu_req_bits_ren2,
  io_rocc_fpu_req_bits_ren3,
  io_rocc_fpu_req_bits_swap12,
  io_rocc_fpu_req_bits_swap23,
  io_rocc_fpu_req_bits_single,
  io_rocc_fpu_req_bits_fromint,
  io_rocc_fpu_req_bits_toint,
  io_rocc_fpu_req_bits_fastpipe,
  io_rocc_fpu_req_bits_fma,
  io_rocc_fpu_req_bits_div,
  io_rocc_fpu_req_bits_sqrt,
  io_rocc_fpu_req_bits_round,
  io_rocc_fpu_req_bits_wflags,
  io_rocc_fpu_req_bits_rm,
  io_rocc_fpu_req_bits_typ,
  io_rocc_fpu_req_bits_in1,
  io_rocc_fpu_req_bits_in2,
  io_rocc_fpu_req_bits_in3,
  io_rocc_fpu_resp_ready,
  io_rocc_csr_waddr,
  io_rocc_csr_wdata,
  io_rocc_csr_wen,
  io_interrupt,
  io_interrupt_cause
);

  input [11:0] io_host_csr_req_bits_addr;
  input [63:0] io_host_csr_req_bits_data;
  output [63:0] io_host_csr_resp_bits;
  input [11:0] io_rw_addr;
  input [2:0] io_rw_cmd;
  output [63:0] io_rw_rdata;
  input [63:0] io_rw_wdata;
  output [30:0] io_status_zero2;
  output [8:0] io_status_zero1;
  output [4:0] io_status_vm;
  output [1:0] io_status_xs;
  output [1:0] io_status_fs;
  output [1:0] io_status_prv3;
  output [1:0] io_status_prv2;
  output [1:0] io_status_prv1;
  output [1:0] io_status_prv;
  output [31:0] io_ptbr;
  output [39:0] io_evec;
  input [63:0] io_cause;
  input [39:0] io_pc;
  output [63:0] io_time;
  output [2:0] io_fcsr_rm;
  input [4:0] io_fcsr_flags_bits;
  input [4:0] io_rocc_resp_bits_rd;
  input [63:0] io_rocc_resp_bits_data;
  input [39:0] io_rocc_mem_req_bits_addr;
  input [9:0] io_rocc_mem_req_bits_tag;
  input [4:0] io_rocc_mem_req_bits_cmd;
  input [2:0] io_rocc_mem_req_bits_typ;
  input [63:0] io_rocc_mem_req_bits_data;
  input [25:0] io_rocc_autl_acquire_bits_addr_block;
  input [5:0] io_rocc_autl_acquire_bits_client_xact_id;
  input [1:0] io_rocc_autl_acquire_bits_addr_beat;
  input [2:0] io_rocc_autl_acquire_bits_a_type;
  input [16:0] io_rocc_autl_acquire_bits_union;
  input [127:0] io_rocc_autl_acquire_bits_data;
  input [4:0] io_rocc_fpu_req_bits_cmd;
  input [2:0] io_rocc_fpu_req_bits_rm;
  input [1:0] io_rocc_fpu_req_bits_typ;
  input [64:0] io_rocc_fpu_req_bits_in1;
  input [64:0] io_rocc_fpu_req_bits_in2;
  input [64:0] io_rocc_fpu_req_bits_in3;
  output [11:0] io_rocc_csr_waddr;
  output [63:0] io_rocc_csr_wdata;
  output [63:0] io_interrupt_cause;
  input clk;
  input reset;
  input io_host_reset;
  input io_host_id;
  input io_host_csr_req_valid;
  input io_host_csr_req_bits_rw;
  input io_host_csr_resp_ready;
  input io_exception;
  input io_retire;
  input io_uarch_counters_15;
  input io_uarch_counters_14;
  input io_uarch_counters_13;
  input io_uarch_counters_12;
  input io_uarch_counters_11;
  input io_uarch_counters_10;
  input io_uarch_counters_9;
  input io_uarch_counters_8;
  input io_uarch_counters_7;
  input io_uarch_counters_6;
  input io_uarch_counters_5;
  input io_uarch_counters_4;
  input io_uarch_counters_3;
  input io_uarch_counters_2;
  input io_uarch_counters_1;
  input io_uarch_counters_0;
  input io_fcsr_flags_valid;
  input io_rocc_cmd_ready;
  input io_rocc_resp_valid;
  input io_rocc_mem_req_valid;
  input io_rocc_mem_req_bits_kill;
  input io_rocc_mem_req_bits_phys;
  input io_rocc_mem_invalidate_lr;
  input io_rocc_busy;
  input io_rocc_interrupt;
  input io_rocc_autl_acquire_valid;
  input io_rocc_autl_acquire_bits_is_builtin_type;
  input io_rocc_autl_grant_ready;
  input io_rocc_fpu_req_valid;
  input io_rocc_fpu_req_bits_ldst;
  input io_rocc_fpu_req_bits_wen;
  input io_rocc_fpu_req_bits_ren1;
  input io_rocc_fpu_req_bits_ren2;
  input io_rocc_fpu_req_bits_ren3;
  input io_rocc_fpu_req_bits_swap12;
  input io_rocc_fpu_req_bits_swap23;
  input io_rocc_fpu_req_bits_single;
  input io_rocc_fpu_req_bits_fromint;
  input io_rocc_fpu_req_bits_toint;
  input io_rocc_fpu_req_bits_fastpipe;
  input io_rocc_fpu_req_bits_fma;
  input io_rocc_fpu_req_bits_div;
  input io_rocc_fpu_req_bits_sqrt;
  input io_rocc_fpu_req_bits_round;
  input io_rocc_fpu_req_bits_wflags;
  input io_rocc_fpu_resp_ready;
  output io_host_csr_req_ready;
  output io_host_csr_resp_valid;
  output io_host_debug_stats_csr;
  output io_csr_stall;
  output io_csr_xcpt;
  output io_eret;
  output io_status_sd;
  output io_status_sd_rv32;
  output io_status_mprv;
  output io_status_ie3;
  output io_status_ie2;
  output io_status_ie1;
  output io_status_ie;
  output io_fatc;
  output io_rocc_csr_wen;
  output io_interrupt;
  wire [63:0] io_rw_rdata,io_rocc_csr_wdata,io_interrupt_cause,T36,T48,T37,T46,T49,T442,T438,
  T447,T443,T450,T477,T451,T491,T478,T495,T492,T513,T531,T580,T593,T581,T606,T594,
  T619,T607,T632,T620,T645,T633,T658,T646,T671,T659,T684,T672,T697,T685,T710,T698,
  T723,T711,T736,T724,T749,T737,T762,T750,T775,T763,T788,T776,T806,T789,T808,T807,
  T810,T809,T821,T811,T826,T828,T830,T829,T832,T831,T837,T833,T842,T838,T846,T843,
  T856,T866,T869,T871,T870,T875,T874,T876,T878,T880,T879,T882,T881,T884,T883,T886,
  T885,T888,T887,T890,T889,T891;
  wire [1:0] io_status_xs,io_status_fs,T218;
  wire [39:0] io_evec,T364,T931,T340,T932,T343,T933,T934,T352,T935,T349;
  wire [11:0] io_rocc_csr_waddr;
  wire io_host_csr_req_ready,io_csr_xcpt,io_eret,io_status_sd,io_fatc,io_rocc_csr_wen,
  io_interrupt,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  T11,insn_break,T7,T9,T17,insn_call,T12,T15,T13,T94,T18,T19,priv_sufficient,T88,T25,
  T76,T69,T52,host_csr_req_fire,T40,T41,cpu_ren,T42,T45,T58,T53,T55,N163,T63,T61,
  cpu_wen,T64,T66,T70,T72,T78,T79,T82,T80,T83,maybe_insn_redirect_trap,T89,T91,
  T214,T95,T96,T104,T97,fp_csr,T98,T99,T101,T213,T105,addr_valid,T107,T109,T111,T113,
  T115,T117,T119,T121,T123,T124,T126,T128,T130,T132,T134,T136,T138,T140,T142,T144,
  T146,T148,T150,T152,T154,T156,T158,T160,T162,T164,T166,T168,T170,T172,T174,T176,
  T178,T180,T182,T184,T186,T188,T190,T192,T193,T195,T197,T199,T201,T203,T205,T207,
  T209,T211,T212,T312,N164,T218_63,T300,N165,T219_0,T285,N166,T220_0,T273,N167,
  T260,N168,T223,T247,T224,T246,T225,T253,T251,T259,T257,T265,T261,T264,T262,T270,
  T278,T274,T277,T275,T290,T286,T289,T287,T297,T293,T295,T301,T304,T302,T307,T311,
  T308,T309,T313,T316,T314,T322,N169,T320,N170,T331,T332,T334,T335,T369,N171,N172,
  N173,T346,N174,N175,T355,N176,N177,T362,N178,T367,T373,T402,T399,T409,T408,
  some_interrupt_pending,insn_wfi,T413,T414,T417,T415,T435,N179,T421,T433,N180,T422,T431,
  N181,T423,T429,N182,T424,T427,N183,T425,T426,T428,T430,T432,T434,T436,T439_39,
  T444_63,T452_63,T474,T465,T463,N184,T466,T468,T470,T490,T488,T486,T485,T494,T949_1,
  T950_1,T532_63,T532_31,T532_4,T532_3,T532_0,T591,T604,T617,T630,T643,T656,T669,
  T682,T695,T708,T721,T734,T747,T760,T773,T786,T798,T803,T817,T814,T815,T816,T820,
  T818,T825,T834_63,T839_63,T845,T899,N185,N186,T906,T905,T907,T910,T909,N187,N188,
  N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,
  N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,
  N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,
  N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,
  N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,
  N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,
  N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,
  N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
  N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,
  N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,
  N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,
  N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,
  N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,
  N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,
  N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,
  N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,
  N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,
  N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,
  N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,
  N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,
  N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,
  N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,
  N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,
  N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,
  N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,
  N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,
  N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,
  N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,
  N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,
  N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,
  N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,
  N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,
  N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,
  N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
  N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,
  N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,
  N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,
  N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,
  N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,
  N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,
  N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,
  N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,
  N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,
  N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,
  N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,
  N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,
  N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,
  N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,
  N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,
  N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,
  N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,
  N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,
  N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,
  N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,
  N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,
  N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,
  N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,
  N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,
  N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,
  N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,
  N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,
  N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,
  N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,
  N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,
  N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,
  N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,
  N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,
  N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,
  N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,
  N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,
  N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,
  N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,
  N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,
  N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,
  N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,
  N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,
  N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,
  N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,
  N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,
  N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,
  N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,
  N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,
  N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,
  N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,
  N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,
  N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,
  N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,
  N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,
  N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,
  N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,
  N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,
  N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,
  N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,
  N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,
  N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,
  N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,
  N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,
  N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,
  N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,
  N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,
  N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,
  N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,
  N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,
  N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,
  N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,
  N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,
  N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,
  N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,
  N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,
  N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,
  N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,
  N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,
  N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,
  N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,
  N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,
  N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,
  N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,
  N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,
  N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,
  N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,
  N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,
  N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,
  N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,
  N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,
  N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,
  N2084,N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,
  N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,
  N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,
  N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,
  N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,
  N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,
  N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,
  N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,
  N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,
  N2204,N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,
  N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,
  N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,
  N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,
  N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,
  N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,
  N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,
  N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,
  N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,
  N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,
  N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,
  N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,
  N2364,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,
  N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,
  N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,
  N2404,N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,
  N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,
  N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,
  N2444,N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,
  N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,
  N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,
  N2484,N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,
  N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,
  N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,
  N2524,N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,
  N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,
  N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,
  N2564,N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,
  N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,
  N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,
  N2604,N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,
  N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,
  N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,
  N2644,N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,
  N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,
  N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,
  N2684,N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,
  N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,
  N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,
  N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,
  N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,
  N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,
  N2764,N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,
  N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,
  N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,
  N2804,N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,
  N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,
  N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,
  N2844,N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,
  N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,
  N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,
  N2884,N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,
  N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,
  N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,
  N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,
  N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,
  N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,
  N2964,N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,
  N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,
  N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,
  N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,
  N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,
  N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,
  N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,
  N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,
  N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,
  N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,
  N3097,N3098,N3099,N3100,N3101,N3102;
  wire [0:0] T914,T216,T1003,T1005;
  wire [63:63] T219,T220,T221,T222,T439,T877;
  wire [2:0] T924,T319,T1024;
  wire [5:0] T325,T585,T598,T611,T624,T637,T650,T663,T676,T689,T702,T715,T728,T741,T754,T767,
  T780,T794;
  wire [6:6] T326,T586,T599,T612,T625,T638,T651,T664,T677,T690,T703,T716,T729,T742,T755,T768,
  T781,T795;
  wire [57:0] T329,T590,T603,T616,T629,T642,T655,T668,T681,T694,T707,T720,T733,T746,T759,T772,
  T785,T802;
  wire [39:2] T344,T350,T353;
  wire [38:0] T936,T359;
  wire [38:2] T360;
  wire [31:0] T945;
  wire [39:39] T457;
  wire [3:0] T947;
  wire [5:5] T949,T950;
  wire [16:12] T532;
  wire [7:0] T1008,T1013,T1020,T893;
  wire [30:30] T1018;
  wire [4:0] T1023,T1021,T896,T1022,T898,T902;
  reg [1:0] io_status_prv,io_status_prv1,io_status_prv2,io_status_prv3,reg_mstatus_fs,
  reg_mstatus_xs;
  reg [63:0] io_host_csr_resp_bits,read_time,reg_mtimecmp,reg_fromhost,io_time,reg_mtvec,
  reg_scause,reg_mcause,reg_sscratch,T582,T595,T608,T621,T634,T647,T660,T673,T686,
  T699,T712,T725,T738,T751,T764,T777,T790,reg_tohost,reg_mscratch;
  reg host_csr_req_valid,host_csr_bits_rw,io_status_ie,io_status_ie1,io_status_ie2,
  T515_1,T497_1,T858_7,T848_7,io_status_ie3,io_status_mprv,io_status_sd_rv32,
  io_csr_stall,io_host_debug_stats_csr,T848_0,T848_6,T858_0,T858_6,io_host_csr_resp_valid;
  reg [11:0] host_csr_bits_addr;
  reg [4:2] T858,T848;
  reg [5:5] T515,T497;
  reg [2:0] io_fcsr_rm;
  reg [40:0] T444,T839,T452,T834;
  reg [38:0] T357;
  reg [31:0] io_ptbr;
  reg [4:0] io_status_vm,T894;
  reg [8:0] io_status_zero1;
  reg [30:0] io_status_zero2;
  assign io_interrupt_cause[62] = 1'b0;
  assign io_interrupt_cause[61] = 1'b0;
  assign io_interrupt_cause[60] = 1'b0;
  assign io_interrupt_cause[59] = 1'b0;
  assign io_interrupt_cause[58] = 1'b0;
  assign io_interrupt_cause[57] = 1'b0;
  assign io_interrupt_cause[56] = 1'b0;
  assign io_interrupt_cause[55] = 1'b0;
  assign io_interrupt_cause[54] = 1'b0;
  assign io_interrupt_cause[53] = 1'b0;
  assign io_interrupt_cause[52] = 1'b0;
  assign io_interrupt_cause[51] = 1'b0;
  assign io_interrupt_cause[50] = 1'b0;
  assign io_interrupt_cause[49] = 1'b0;
  assign io_interrupt_cause[48] = 1'b0;
  assign io_interrupt_cause[47] = 1'b0;
  assign io_interrupt_cause[46] = 1'b0;
  assign io_interrupt_cause[45] = 1'b0;
  assign io_interrupt_cause[44] = 1'b0;
  assign io_interrupt_cause[43] = 1'b0;
  assign io_interrupt_cause[42] = 1'b0;
  assign io_interrupt_cause[41] = 1'b0;
  assign io_interrupt_cause[40] = 1'b0;
  assign io_interrupt_cause[39] = 1'b0;
  assign io_interrupt_cause[38] = 1'b0;
  assign io_interrupt_cause[37] = 1'b0;
  assign io_interrupt_cause[36] = 1'b0;
  assign io_interrupt_cause[35] = 1'b0;
  assign io_interrupt_cause[34] = 1'b0;
  assign io_interrupt_cause[33] = 1'b0;
  assign io_interrupt_cause[32] = 1'b0;
  assign io_interrupt_cause[31] = 1'b0;
  assign io_interrupt_cause[30] = 1'b0;
  assign io_interrupt_cause[29] = 1'b0;
  assign io_interrupt_cause[28] = 1'b0;
  assign io_interrupt_cause[27] = 1'b0;
  assign io_interrupt_cause[26] = 1'b0;
  assign io_interrupt_cause[25] = 1'b0;
  assign io_interrupt_cause[24] = 1'b0;
  assign io_interrupt_cause[23] = 1'b0;
  assign io_interrupt_cause[22] = 1'b0;
  assign io_interrupt_cause[21] = 1'b0;
  assign io_interrupt_cause[20] = 1'b0;
  assign io_interrupt_cause[19] = 1'b0;
  assign io_interrupt_cause[18] = 1'b0;
  assign io_interrupt_cause[17] = 1'b0;
  assign io_interrupt_cause[16] = 1'b0;
  assign io_interrupt_cause[15] = 1'b0;
  assign io_interrupt_cause[14] = 1'b0;
  assign io_interrupt_cause[13] = 1'b0;
  assign io_interrupt_cause[12] = 1'b0;
  assign io_interrupt_cause[11] = 1'b0;
  assign io_interrupt_cause[10] = 1'b0;
  assign io_interrupt_cause[9] = 1'b0;
  assign io_interrupt_cause[8] = 1'b0;
  assign io_interrupt_cause[7] = 1'b0;
  assign io_interrupt_cause[6] = 1'b0;
  assign io_interrupt_cause[5] = 1'b0;
  assign io_interrupt_cause[4] = 1'b0;
  assign io_interrupt_cause[3] = 1'b0;
  assign io_interrupt_cause[2] = 1'b0;
  assign io_interrupt = io_interrupt_cause[63];
  assign priv_sufficient = io_rw_addr[9:8] <= io_status_prv;
  assign T99 = io_status_fs != 1'b0;
  assign T264 = io_status_prv < { 1'b1, 1'b1 };
  assign T289 = io_status_prv < { 1'b1, 1'b1 };
  assign T293 = reg_mtimecmp <= read_time;
  assign T304 = io_status_prv < { 1'b1, 1'b1 };
  assign T316 = io_status_prv < { 1'b1, 1'b1 };
  assign T408 = io_status_xs == { 1'b1, 1'b1 };
  assign T409 = io_status_fs == { 1'b1, 1'b1 };
  assign T426 = io_status_prv <= 1'b1;
  assign T428 = io_status_prv <= { 1'b1, 1'b1 };
  assign T430 = io_status_prv <= 1'b1;
  assign T432 = io_status_prv <= { 1'b1, 1'b1 };
  assign T434 = io_status_prv <= { 1'b1, 1'b1 };
  assign T436 = io_status_prv <= { 1'b1, 1'b1 };
  assign T463 = $signed(io_rw_wdata[38:0]) < $signed(1'b0);

  always @(posedge clk) begin
    if(N192) begin
      io_status_prv[1] <= N194;
    end 
  end


  always @(posedge clk) begin
    if(N192) begin
      io_status_prv[0] <= N193;
    end 
  end


  always @(posedge clk) begin
    if(N200) begin
      io_status_prv1[1] <= N202;
    end 
  end


  always @(posedge clk) begin
    if(N200) begin
      io_status_prv1[0] <= N201;
    end 
  end


  always @(posedge clk) begin
    if(N207) begin
      io_status_prv2[1] <= N209;
    end 
  end


  always @(posedge clk) begin
    if(N207) begin
      io_status_prv2[0] <= N208;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[63] <= N276;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[62] <= N275;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[61] <= N274;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[60] <= N273;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[59] <= N272;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[58] <= N271;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[57] <= N270;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[56] <= N269;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[55] <= N268;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[54] <= N267;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[53] <= N266;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[52] <= N265;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[51] <= N264;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[50] <= N263;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[49] <= N262;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[48] <= N261;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[47] <= N260;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[46] <= N259;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[45] <= N258;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[44] <= N257;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[43] <= N256;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[42] <= N255;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[41] <= N254;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[40] <= N253;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[39] <= N252;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[38] <= N251;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[37] <= N250;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[36] <= N249;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[35] <= N248;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[34] <= N247;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[33] <= N246;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[32] <= N245;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[31] <= N244;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[30] <= N243;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[29] <= N242;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[28] <= N241;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[27] <= N240;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[26] <= N239;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[25] <= N238;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[24] <= N237;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[23] <= N236;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[22] <= N235;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[21] <= N234;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[20] <= N233;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[19] <= N232;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[18] <= N231;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[17] <= N230;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[16] <= N229;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[15] <= N228;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[14] <= N227;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[13] <= N226;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[12] <= N225;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[11] <= N224;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[10] <= N223;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[9] <= N222;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[8] <= N221;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[7] <= N220;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[6] <= N219;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[5] <= N218;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[4] <= N217;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[3] <= N216;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[2] <= N215;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[1] <= N214;
    end 
  end


  always @(posedge clk) begin
    if(N212) begin
      io_host_csr_resp_bits[0] <= N213;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      host_csr_req_valid <= N278;
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[11] <= io_host_csr_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[10] <= io_host_csr_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[9] <= io_host_csr_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[8] <= io_host_csr_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[7] <= io_host_csr_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[6] <= io_host_csr_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[5] <= io_host_csr_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[4] <= io_host_csr_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[3] <= io_host_csr_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[2] <= io_host_csr_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[1] <= io_host_csr_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_addr[0] <= io_host_csr_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(T40) begin
      host_csr_bits_rw <= io_host_csr_req_bits_rw;
    end 
  end


  always @(posedge clk) begin
    if(N284) begin
      io_status_ie <= N285;
    end 
  end


  always @(posedge clk) begin
    if(N291) begin
      io_status_ie1 <= N292;
    end 
  end


  always @(posedge clk) begin
    if(N297) begin
      io_status_ie2 <= N298;
    end 
  end


  always @(posedge clk) begin
    if(N302) begin
      T515_1 <= N303;
    end 
  end


  always @(posedge clk) begin
    if(N307) begin
      T497_1 <= N308;
    end 
  end


  always @(posedge clk) begin
    if(N312) begin
      T858[3] <= N313;
    end 
  end


  always @(posedge clk) begin
    if(N316) begin
      T848[3] <= N317;
    end 
  end


  always @(posedge clk) begin
    if(N320) begin
      T515[5] <= N321;
    end 
  end


  always @(posedge clk) begin
    if(N325) begin
      T497[5] <= N326;
    end 
  end


  always @(posedge clk) begin
    if(N330) begin
      T858_7 <= N331;
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[63] <= io_rocc_csr_wdata[63];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[62] <= io_rocc_csr_wdata[62];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[61] <= io_rocc_csr_wdata[61];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[60] <= io_rocc_csr_wdata[60];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[59] <= io_rocc_csr_wdata[59];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[58] <= io_rocc_csr_wdata[58];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[57] <= io_rocc_csr_wdata[57];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[56] <= io_rocc_csr_wdata[56];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[55] <= io_rocc_csr_wdata[55];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[54] <= io_rocc_csr_wdata[54];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[53] <= io_rocc_csr_wdata[53];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[52] <= io_rocc_csr_wdata[52];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[51] <= io_rocc_csr_wdata[51];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[50] <= io_rocc_csr_wdata[50];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[49] <= io_rocc_csr_wdata[49];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[48] <= io_rocc_csr_wdata[48];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[47] <= io_rocc_csr_wdata[47];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[46] <= io_rocc_csr_wdata[46];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[45] <= io_rocc_csr_wdata[45];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[44] <= io_rocc_csr_wdata[44];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[43] <= io_rocc_csr_wdata[43];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[42] <= io_rocc_csr_wdata[42];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[41] <= io_rocc_csr_wdata[41];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[40] <= io_rocc_csr_wdata[40];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[39] <= io_rocc_csr_wdata[39];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[38] <= io_rocc_csr_wdata[38];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[37] <= io_rocc_csr_wdata[37];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[36] <= io_rocc_csr_wdata[36];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[35] <= io_rocc_csr_wdata[35];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[34] <= io_rocc_csr_wdata[34];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[33] <= io_rocc_csr_wdata[33];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[32] <= io_rocc_csr_wdata[32];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[31] <= io_rocc_csr_wdata[31];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[30] <= io_rocc_csr_wdata[30];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[29] <= io_rocc_csr_wdata[29];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[28] <= io_rocc_csr_wdata[28];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[27] <= io_rocc_csr_wdata[27];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[26] <= io_rocc_csr_wdata[26];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[25] <= io_rocc_csr_wdata[25];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[24] <= io_rocc_csr_wdata[24];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[23] <= io_rocc_csr_wdata[23];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[22] <= io_rocc_csr_wdata[22];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[21] <= io_rocc_csr_wdata[21];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[20] <= io_rocc_csr_wdata[20];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[19] <= io_rocc_csr_wdata[19];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[18] <= io_rocc_csr_wdata[18];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[17] <= io_rocc_csr_wdata[17];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[16] <= io_rocc_csr_wdata[16];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[15] <= io_rocc_csr_wdata[15];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[14] <= io_rocc_csr_wdata[14];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[13] <= io_rocc_csr_wdata[13];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[12] <= io_rocc_csr_wdata[12];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[11] <= io_rocc_csr_wdata[11];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[10] <= io_rocc_csr_wdata[10];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[9] <= io_rocc_csr_wdata[9];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[8] <= io_rocc_csr_wdata[8];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[7] <= io_rocc_csr_wdata[7];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[6] <= io_rocc_csr_wdata[6];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[5] <= io_rocc_csr_wdata[5];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[4] <= io_rocc_csr_wdata[4];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[3] <= io_rocc_csr_wdata[3];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[2] <= io_rocc_csr_wdata[2];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[1] <= io_rocc_csr_wdata[1];
    end 
  end


  always @(posedge clk) begin
    if(T295) begin
      read_time[0] <= io_rocc_csr_wdata[0];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[63] <= io_rocc_csr_wdata[63];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[62] <= io_rocc_csr_wdata[62];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[61] <= io_rocc_csr_wdata[61];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[60] <= io_rocc_csr_wdata[60];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[59] <= io_rocc_csr_wdata[59];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[58] <= io_rocc_csr_wdata[58];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[57] <= io_rocc_csr_wdata[57];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[56] <= io_rocc_csr_wdata[56];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[55] <= io_rocc_csr_wdata[55];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[54] <= io_rocc_csr_wdata[54];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[53] <= io_rocc_csr_wdata[53];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[52] <= io_rocc_csr_wdata[52];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[51] <= io_rocc_csr_wdata[51];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[50] <= io_rocc_csr_wdata[50];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[49] <= io_rocc_csr_wdata[49];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[48] <= io_rocc_csr_wdata[48];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[47] <= io_rocc_csr_wdata[47];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[46] <= io_rocc_csr_wdata[46];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[45] <= io_rocc_csr_wdata[45];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[44] <= io_rocc_csr_wdata[44];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[43] <= io_rocc_csr_wdata[43];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[42] <= io_rocc_csr_wdata[42];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[41] <= io_rocc_csr_wdata[41];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[40] <= io_rocc_csr_wdata[40];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[39] <= io_rocc_csr_wdata[39];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[38] <= io_rocc_csr_wdata[38];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[37] <= io_rocc_csr_wdata[37];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[36] <= io_rocc_csr_wdata[36];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[35] <= io_rocc_csr_wdata[35];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[34] <= io_rocc_csr_wdata[34];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[33] <= io_rocc_csr_wdata[33];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[32] <= io_rocc_csr_wdata[32];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[31] <= io_rocc_csr_wdata[31];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[30] <= io_rocc_csr_wdata[30];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[29] <= io_rocc_csr_wdata[29];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[28] <= io_rocc_csr_wdata[28];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[27] <= io_rocc_csr_wdata[27];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[26] <= io_rocc_csr_wdata[26];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[25] <= io_rocc_csr_wdata[25];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[24] <= io_rocc_csr_wdata[24];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[23] <= io_rocc_csr_wdata[23];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[22] <= io_rocc_csr_wdata[22];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[21] <= io_rocc_csr_wdata[21];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[20] <= io_rocc_csr_wdata[20];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[19] <= io_rocc_csr_wdata[19];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[18] <= io_rocc_csr_wdata[18];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[17] <= io_rocc_csr_wdata[17];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[16] <= io_rocc_csr_wdata[16];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[15] <= io_rocc_csr_wdata[15];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[14] <= io_rocc_csr_wdata[14];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[13] <= io_rocc_csr_wdata[13];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[12] <= io_rocc_csr_wdata[12];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[11] <= io_rocc_csr_wdata[11];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[10] <= io_rocc_csr_wdata[10];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[9] <= io_rocc_csr_wdata[9];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[8] <= io_rocc_csr_wdata[8];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[7] <= io_rocc_csr_wdata[7];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[6] <= io_rocc_csr_wdata[6];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[5] <= io_rocc_csr_wdata[5];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[4] <= io_rocc_csr_wdata[4];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[3] <= io_rocc_csr_wdata[3];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[2] <= io_rocc_csr_wdata[2];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[1] <= io_rocc_csr_wdata[1];
    end 
  end


  always @(posedge clk) begin
    if(T297) begin
      reg_mtimecmp[0] <= io_rocc_csr_wdata[0];
    end 
  end


  always @(posedge clk) begin
    if(N334) begin
      T848_7 <= N335;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[63] <= N402;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[62] <= N401;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[61] <= N400;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[60] <= N399;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[59] <= N398;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[58] <= N397;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[57] <= N396;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[56] <= N395;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[55] <= N394;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[54] <= N393;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[53] <= N392;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[52] <= N391;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[51] <= N390;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[50] <= N389;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[49] <= N388;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[48] <= N387;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[47] <= N386;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[46] <= N385;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[45] <= N384;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[44] <= N383;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[43] <= N382;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[42] <= N381;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[41] <= N380;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[40] <= N379;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[39] <= N378;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[38] <= N377;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[37] <= N376;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[36] <= N375;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[35] <= N374;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[34] <= N373;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[33] <= N372;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[32] <= N371;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[31] <= N370;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[30] <= N369;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[29] <= N368;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[28] <= N367;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[27] <= N366;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[26] <= N365;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[25] <= N364;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[24] <= N363;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[23] <= N362;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[22] <= N361;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[21] <= N360;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[20] <= N359;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[19] <= N358;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[18] <= N357;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[17] <= N356;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[16] <= N355;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[15] <= N354;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[14] <= N353;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[13] <= N352;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[12] <= N351;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[11] <= N350;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[10] <= N349;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[9] <= N348;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[8] <= N347;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[7] <= N346;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[6] <= N345;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[5] <= N344;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[4] <= N343;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[3] <= N342;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[2] <= N341;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[1] <= N340;
    end 
  end


  always @(posedge clk) begin
    if(N338) begin
      reg_fromhost[0] <= N339;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_fcsr_rm[2] <= T924[2];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_fcsr_rm[1] <= T924[1];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_fcsr_rm[0] <= T924[0];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_time[5] <= N409;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_time[4] <= N408;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_time[3] <= N407;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_time[2] <= N406;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_time[1] <= N405;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      io_time[0] <= N404;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[63] <= N470;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[62] <= N469;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[61] <= N468;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[60] <= N467;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[59] <= N466;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[58] <= N465;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[57] <= N464;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[56] <= N463;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[55] <= N462;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[54] <= N461;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[53] <= N460;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[52] <= N459;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[51] <= N458;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[50] <= N457;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[49] <= N456;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[48] <= N455;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[47] <= N454;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[46] <= N453;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[45] <= N452;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[44] <= N451;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[43] <= N450;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[42] <= N449;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[41] <= N448;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[40] <= N447;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[39] <= N446;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[38] <= N445;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[37] <= N444;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[36] <= N443;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[35] <= N442;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[34] <= N441;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[33] <= N440;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[32] <= N439;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[31] <= N438;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[30] <= N437;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[29] <= N436;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[28] <= N435;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[27] <= N434;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[26] <= N433;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[25] <= N432;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[24] <= N431;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[23] <= N430;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[22] <= N429;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[21] <= N428;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[20] <= N427;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[19] <= N426;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[18] <= N425;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[17] <= N424;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[16] <= N423;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[15] <= N422;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[14] <= N421;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[13] <= N420;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[12] <= N419;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[11] <= N418;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[10] <= N417;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[9] <= N416;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[8] <= N415;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[7] <= N414;
    end 
  end


  always @(posedge clk) begin
    if(N412) begin
      io_time[6] <= N413;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[39] <= T932[39];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[38] <= T932[38];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[37] <= T932[37];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[36] <= T932[36];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[35] <= T932[35];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[34] <= T932[34];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[33] <= T932[33];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[32] <= T932[32];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[31] <= T932[31];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[30] <= T932[30];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[29] <= T932[29];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[28] <= T932[28];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[27] <= T932[27];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[26] <= T932[26];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[25] <= T932[25];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[24] <= T932[24];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[23] <= T932[23];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[22] <= T932[22];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[21] <= T932[21];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[20] <= T932[20];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[19] <= T932[19];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[18] <= T932[18];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[17] <= T932[17];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[16] <= T932[16];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[15] <= T932[15];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[14] <= T932[14];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[13] <= T932[13];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[12] <= T932[12];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[11] <= T932[11];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[10] <= T932[10];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[9] <= T932[9];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[8] <= T932[8];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[7] <= T932[7];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[6] <= T932[6];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[5] <= T932[5];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[4] <= T932[4];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[3] <= T932[3];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[2] <= T932[2];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[1] <= T932[1];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T444[0] <= T932[0];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[39] <= T934[39];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[38] <= T934[38];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[37] <= T934[37];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[36] <= T934[36];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[35] <= T934[35];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[34] <= T934[34];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[33] <= T934[33];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[32] <= T934[32];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[31] <= T934[31];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[30] <= T934[30];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[29] <= T934[29];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[28] <= T934[28];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[27] <= T934[27];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[26] <= T934[26];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[25] <= T934[25];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[24] <= T934[24];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[23] <= T934[23];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[22] <= T934[22];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[21] <= T934[21];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[20] <= T934[20];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[19] <= T934[19];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[18] <= T934[18];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[17] <= T934[17];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[16] <= T934[16];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[15] <= T934[15];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[14] <= T934[14];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[13] <= T934[13];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[12] <= T934[12];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[11] <= T934[11];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[10] <= T934[10];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[9] <= T934[9];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[8] <= T934[8];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[7] <= T934[7];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[6] <= T934[6];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[5] <= T934[5];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[4] <= T934[4];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[3] <= T934[3];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[2] <= T934[2];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[1] <= T934[1];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T839[0] <= T934[0];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[38] <= T936[38];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[37] <= T936[37];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[36] <= T936[36];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[35] <= T936[35];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[34] <= T936[34];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[33] <= T936[33];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[32] <= T936[32];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[31] <= T936[31];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[30] <= T936[30];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[29] <= T936[29];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[28] <= T936[28];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[27] <= T936[27];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[26] <= T936[26];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[25] <= T936[25];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[24] <= T936[24];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[23] <= T936[23];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[22] <= T936[22];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[21] <= T936[21];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[20] <= T936[20];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[19] <= T936[19];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[18] <= T936[18];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[17] <= T936[17];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[16] <= T936[16];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[15] <= T936[15];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[14] <= T936[14];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[13] <= T936[13];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[12] <= T936[12];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[11] <= T936[11];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[10] <= T936[10];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[9] <= T936[9];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[8] <= T936[8];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[7] <= T936[7];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[6] <= T936[6];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[5] <= T936[5];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[4] <= T936[4];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[3] <= T936[3];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[2] <= T936[2];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[1] <= T936[1];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T357[0] <= T936[0];
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[63] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[62] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[61] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[60] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[59] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[58] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[57] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[56] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[55] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[54] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[53] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[52] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[51] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[50] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[49] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[48] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[47] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[46] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[45] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[44] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[43] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[42] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[41] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[40] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[39] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[38] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[37] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[36] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[35] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[34] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[33] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[32] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[31] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[30] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[29] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[28] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[27] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[26] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[25] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[24] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[23] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[22] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[21] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[20] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[19] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[18] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[17] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[16] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[15] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[14] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[13] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[12] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[11] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[10] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[9] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[8] <= reset;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[7] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[6] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[5] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[3] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[1] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N473) begin
      reg_mtvec[0] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[31] <= io_rocc_csr_wdata[31];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[30] <= io_rocc_csr_wdata[30];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[29] <= io_rocc_csr_wdata[29];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[28] <= io_rocc_csr_wdata[28];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[27] <= io_rocc_csr_wdata[27];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[26] <= io_rocc_csr_wdata[26];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[25] <= io_rocc_csr_wdata[25];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[24] <= io_rocc_csr_wdata[24];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[23] <= io_rocc_csr_wdata[23];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[22] <= io_rocc_csr_wdata[22];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[21] <= io_rocc_csr_wdata[21];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[20] <= io_rocc_csr_wdata[20];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[19] <= io_rocc_csr_wdata[19];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[18] <= io_rocc_csr_wdata[18];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[17] <= io_rocc_csr_wdata[17];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[16] <= io_rocc_csr_wdata[16];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[15] <= io_rocc_csr_wdata[15];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[14] <= io_rocc_csr_wdata[14];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[13] <= io_rocc_csr_wdata[13];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[12] <= io_rocc_csr_wdata[12];
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[11] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[10] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[9] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[8] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[7] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[6] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[5] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[3] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[1] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(T373) begin
      io_ptbr[0] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_ie3 <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_prv3[1] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_prv3[0] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N477) begin
      reg_mstatus_fs[1] <= N479;
    end 
  end


  always @(posedge clk) begin
    if(N477) begin
      reg_mstatus_fs[0] <= N478;
    end 
  end


  always @(posedge clk) begin
    if(N483) begin
      reg_mstatus_xs[1] <= N485;
    end 
  end


  always @(posedge clk) begin
    if(N483) begin
      reg_mstatus_xs[0] <= N484;
    end 
  end


  always @(posedge clk) begin
    if(N490) begin
      io_status_mprv <= N491;
    end 
  end


  always @(posedge clk) begin
    if(N495) begin
      io_status_vm[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N495) begin
      io_status_vm[3] <= N496;
    end 
  end


  always @(posedge clk) begin
    if(N495) begin
      io_status_vm[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N495) begin
      io_status_vm[1] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N495) begin
      io_status_vm[0] <= N496;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[8] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[7] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[6] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[5] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[3] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[1] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero1[0] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_sd_rv32 <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[30] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[29] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[28] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[27] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[26] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[25] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[24] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[23] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[22] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[21] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[20] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[19] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[18] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[17] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[16] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[15] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[14] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[13] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[12] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[11] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[10] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[9] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[8] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[7] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[6] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[5] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[3] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[1] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      io_status_zero2[0] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N500) begin
      io_csr_stall <= N501;
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[39] <= T834[39];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[38] <= T834[38];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[37] <= T834[37];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[36] <= T834[36];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[35] <= T834[35];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[34] <= T834[34];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[33] <= T834[33];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[32] <= T834[32];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[31] <= T834[31];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[30] <= T834[30];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[29] <= T834[29];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[28] <= T834[28];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[27] <= T834[27];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[26] <= T834[26];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[25] <= T834[25];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[24] <= T834[24];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[23] <= T834[23];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[22] <= T834[22];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[21] <= T834[21];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[20] <= T834[20];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[19] <= T834[19];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[18] <= T834[18];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[17] <= T834[17];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[16] <= T834[16];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[15] <= T834[15];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[14] <= T834[14];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[13] <= T834[13];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[12] <= T834[12];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[11] <= T834[11];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[10] <= T834[10];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[9] <= T834[9];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[8] <= T834[8];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[7] <= T834[7];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[6] <= T834[6];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[5] <= T834[5];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[4] <= T834[4];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[3] <= T834[3];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[2] <= T834[2];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[1] <= T834[1];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      T452[0] <= T834[0];
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[39] <= N545;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[38] <= N544;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[37] <= N543;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[36] <= N542;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[35] <= N541;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[34] <= N540;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[33] <= N539;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[32] <= N538;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[31] <= N537;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[30] <= N536;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[29] <= N535;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[28] <= N534;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[27] <= N533;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[26] <= N532;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[25] <= N531;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[24] <= N530;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[23] <= N529;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[22] <= N528;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[21] <= N527;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[20] <= N526;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[19] <= N525;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[18] <= N524;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[17] <= N523;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[16] <= N522;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[15] <= N521;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[14] <= N520;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[13] <= N519;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[12] <= N518;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[11] <= N517;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[10] <= N516;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[9] <= N515;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[8] <= N514;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[7] <= N513;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[6] <= N512;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[5] <= N511;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[4] <= N510;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[3] <= N509;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[2] <= N508;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[1] <= N507;
    end 
  end


  always @(posedge clk) begin
    if(N505) begin
      T834[0] <= N506;
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[63] <= reg_mcause[63];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[62] <= reg_mcause[62];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[61] <= reg_mcause[61];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[60] <= reg_mcause[60];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[59] <= reg_mcause[59];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[58] <= reg_mcause[58];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[57] <= reg_mcause[57];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[56] <= reg_mcause[56];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[55] <= reg_mcause[55];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[54] <= reg_mcause[54];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[53] <= reg_mcause[53];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[52] <= reg_mcause[52];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[51] <= reg_mcause[51];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[50] <= reg_mcause[50];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[49] <= reg_mcause[49];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[48] <= reg_mcause[48];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[47] <= reg_mcause[47];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[46] <= reg_mcause[46];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[45] <= reg_mcause[45];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[44] <= reg_mcause[44];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[43] <= reg_mcause[43];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[42] <= reg_mcause[42];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[41] <= reg_mcause[41];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[40] <= reg_mcause[40];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[39] <= reg_mcause[39];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[38] <= reg_mcause[38];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[37] <= reg_mcause[37];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[36] <= reg_mcause[36];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[35] <= reg_mcause[35];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[34] <= reg_mcause[34];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[33] <= reg_mcause[33];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[32] <= reg_mcause[32];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[31] <= reg_mcause[31];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[30] <= reg_mcause[30];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[29] <= reg_mcause[29];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[28] <= reg_mcause[28];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[27] <= reg_mcause[27];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[26] <= reg_mcause[26];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[25] <= reg_mcause[25];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[24] <= reg_mcause[24];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[23] <= reg_mcause[23];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[22] <= reg_mcause[22];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[21] <= reg_mcause[21];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[20] <= reg_mcause[20];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[19] <= reg_mcause[19];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[18] <= reg_mcause[18];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[17] <= reg_mcause[17];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[16] <= reg_mcause[16];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[15] <= reg_mcause[15];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[14] <= reg_mcause[14];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[13] <= reg_mcause[13];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[12] <= reg_mcause[12];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[11] <= reg_mcause[11];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[10] <= reg_mcause[10];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[9] <= reg_mcause[9];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[8] <= reg_mcause[8];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[7] <= reg_mcause[7];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[6] <= reg_mcause[6];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[5] <= reg_mcause[5];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[4] <= reg_mcause[4];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[3] <= reg_mcause[3];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[2] <= reg_mcause[2];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[1] <= reg_mcause[1];
    end 
  end


  always @(posedge clk) begin
    if(T216[0]) begin
      reg_scause[0] <= reg_mcause[0];
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[63] <= N615;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[62] <= N614;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[61] <= N613;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[60] <= N612;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[59] <= N611;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[58] <= N610;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[57] <= N609;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[56] <= N608;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[55] <= N607;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[54] <= N606;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[53] <= N605;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[52] <= N604;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[51] <= N603;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[50] <= N602;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[49] <= N601;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[48] <= N600;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[47] <= N599;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[46] <= N598;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[45] <= N597;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[44] <= N596;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[43] <= N595;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[42] <= N594;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[41] <= N593;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[40] <= N592;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[39] <= N591;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[38] <= N590;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[37] <= N589;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[36] <= N588;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[35] <= N587;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[34] <= N586;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[33] <= N585;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[32] <= N584;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[31] <= N583;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[30] <= N582;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[29] <= N581;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[28] <= N580;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[27] <= N579;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[26] <= N578;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[25] <= N577;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[24] <= N576;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[23] <= N575;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[22] <= N574;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[21] <= N573;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[20] <= N572;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[19] <= N571;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[18] <= N570;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[17] <= N569;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[16] <= N568;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[15] <= N567;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[14] <= N566;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[13] <= N565;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[12] <= N564;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[11] <= N563;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[10] <= N562;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[9] <= N561;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[8] <= N560;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[7] <= N559;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[6] <= N558;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[5] <= N557;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[4] <= N556;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[3] <= N555;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[2] <= N554;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[1] <= N553;
    end 
  end


  always @(posedge clk) begin
    if(N551) begin
      reg_mcause[0] <= N552;
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[63] <= io_rocc_csr_wdata[63];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[62] <= io_rocc_csr_wdata[62];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[61] <= io_rocc_csr_wdata[61];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[60] <= io_rocc_csr_wdata[60];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[59] <= io_rocc_csr_wdata[59];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[58] <= io_rocc_csr_wdata[58];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[57] <= io_rocc_csr_wdata[57];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[56] <= io_rocc_csr_wdata[56];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[55] <= io_rocc_csr_wdata[55];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[54] <= io_rocc_csr_wdata[54];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[53] <= io_rocc_csr_wdata[53];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[52] <= io_rocc_csr_wdata[52];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[51] <= io_rocc_csr_wdata[51];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[50] <= io_rocc_csr_wdata[50];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[49] <= io_rocc_csr_wdata[49];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[48] <= io_rocc_csr_wdata[48];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[47] <= io_rocc_csr_wdata[47];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[46] <= io_rocc_csr_wdata[46];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[45] <= io_rocc_csr_wdata[45];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[44] <= io_rocc_csr_wdata[44];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[43] <= io_rocc_csr_wdata[43];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[42] <= io_rocc_csr_wdata[42];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[41] <= io_rocc_csr_wdata[41];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[40] <= io_rocc_csr_wdata[40];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[39] <= io_rocc_csr_wdata[39];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[38] <= io_rocc_csr_wdata[38];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[37] <= io_rocc_csr_wdata[37];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[36] <= io_rocc_csr_wdata[36];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[35] <= io_rocc_csr_wdata[35];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[34] <= io_rocc_csr_wdata[34];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[33] <= io_rocc_csr_wdata[33];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[32] <= io_rocc_csr_wdata[32];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[31] <= io_rocc_csr_wdata[31];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[30] <= io_rocc_csr_wdata[30];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[29] <= io_rocc_csr_wdata[29];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[28] <= io_rocc_csr_wdata[28];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[27] <= io_rocc_csr_wdata[27];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[26] <= io_rocc_csr_wdata[26];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[25] <= io_rocc_csr_wdata[25];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[24] <= io_rocc_csr_wdata[24];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[23] <= io_rocc_csr_wdata[23];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[22] <= io_rocc_csr_wdata[22];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[21] <= io_rocc_csr_wdata[21];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[20] <= io_rocc_csr_wdata[20];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[19] <= io_rocc_csr_wdata[19];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[18] <= io_rocc_csr_wdata[18];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[17] <= io_rocc_csr_wdata[17];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[16] <= io_rocc_csr_wdata[16];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[15] <= io_rocc_csr_wdata[15];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[14] <= io_rocc_csr_wdata[14];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[13] <= io_rocc_csr_wdata[13];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[12] <= io_rocc_csr_wdata[12];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[11] <= io_rocc_csr_wdata[11];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[10] <= io_rocc_csr_wdata[10];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[9] <= io_rocc_csr_wdata[9];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[8] <= io_rocc_csr_wdata[8];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[7] <= io_rocc_csr_wdata[7];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[6] <= io_rocc_csr_wdata[6];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[5] <= io_rocc_csr_wdata[5];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[4] <= io_rocc_csr_wdata[4];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[3] <= io_rocc_csr_wdata[3];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[2] <= io_rocc_csr_wdata[2];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[1] <= io_rocc_csr_wdata[1];
    end 
  end


  always @(posedge clk) begin
    if(T494) begin
      reg_sscratch[0] <= io_rocc_csr_wdata[0];
    end 
  end


  always @(posedge clk) begin
    if(N618) begin
      T582[5] <= N624;
    end 
  end


  always @(posedge clk) begin
    if(N618) begin
      T582[4] <= N623;
    end 
  end


  always @(posedge clk) begin
    if(N618) begin
      T582[3] <= N622;
    end 
  end


  always @(posedge clk) begin
    if(N618) begin
      T582[2] <= N621;
    end 
  end


  always @(posedge clk) begin
    if(N618) begin
      T582[1] <= N620;
    end 
  end


  always @(posedge clk) begin
    if(N618) begin
      T582[0] <= N619;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[63] <= N685;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[62] <= N684;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[61] <= N683;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[60] <= N682;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[59] <= N681;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[58] <= N680;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[57] <= N679;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[56] <= N678;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[55] <= N677;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[54] <= N676;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[53] <= N675;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[52] <= N674;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[51] <= N673;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[50] <= N672;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[49] <= N671;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[48] <= N670;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[47] <= N669;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[46] <= N668;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[45] <= N667;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[44] <= N666;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[43] <= N665;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[42] <= N664;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[41] <= N663;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[40] <= N662;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[39] <= N661;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[38] <= N660;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[37] <= N659;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[36] <= N658;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[35] <= N657;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[34] <= N656;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[33] <= N655;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[32] <= N654;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[31] <= N653;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[30] <= N652;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[29] <= N651;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[28] <= N650;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[27] <= N649;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[26] <= N648;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[25] <= N647;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[24] <= N646;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[23] <= N645;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[22] <= N644;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[21] <= N643;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[20] <= N642;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[19] <= N641;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[18] <= N640;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[17] <= N639;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[16] <= N638;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[15] <= N637;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[14] <= N636;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[13] <= N635;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[12] <= N634;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[11] <= N633;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[10] <= N632;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[9] <= N631;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[8] <= N630;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[7] <= N629;
    end 
  end


  always @(posedge clk) begin
    if(N627) begin
      T582[6] <= N628;
    end 
  end


  always @(posedge clk) begin
    if(N688) begin
      T595[5] <= N694;
    end 
  end


  always @(posedge clk) begin
    if(N688) begin
      T595[4] <= N693;
    end 
  end


  always @(posedge clk) begin
    if(N688) begin
      T595[3] <= N692;
    end 
  end


  always @(posedge clk) begin
    if(N688) begin
      T595[2] <= N691;
    end 
  end


  always @(posedge clk) begin
    if(N688) begin
      T595[1] <= N690;
    end 
  end


  always @(posedge clk) begin
    if(N688) begin
      T595[0] <= N689;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[63] <= N755;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[62] <= N754;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[61] <= N753;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[60] <= N752;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[59] <= N751;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[58] <= N750;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[57] <= N749;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[56] <= N748;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[55] <= N747;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[54] <= N746;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[53] <= N745;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[52] <= N744;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[51] <= N743;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[50] <= N742;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[49] <= N741;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[48] <= N740;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[47] <= N739;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[46] <= N738;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[45] <= N737;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[44] <= N736;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[43] <= N735;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[42] <= N734;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[41] <= N733;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[40] <= N732;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[39] <= N731;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[38] <= N730;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[37] <= N729;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[36] <= N728;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[35] <= N727;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[34] <= N726;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[33] <= N725;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[32] <= N724;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[31] <= N723;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[30] <= N722;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[29] <= N721;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[28] <= N720;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[27] <= N719;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[26] <= N718;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[25] <= N717;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[24] <= N716;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[23] <= N715;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[22] <= N714;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[21] <= N713;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[20] <= N712;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[19] <= N711;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[18] <= N710;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[17] <= N709;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[16] <= N708;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[15] <= N707;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[14] <= N706;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[13] <= N705;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[12] <= N704;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[11] <= N703;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[10] <= N702;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[9] <= N701;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[8] <= N700;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[7] <= N699;
    end 
  end


  always @(posedge clk) begin
    if(N697) begin
      T595[6] <= N698;
    end 
  end


  always @(posedge clk) begin
    if(N758) begin
      T608[5] <= N764;
    end 
  end


  always @(posedge clk) begin
    if(N758) begin
      T608[4] <= N763;
    end 
  end


  always @(posedge clk) begin
    if(N758) begin
      T608[3] <= N762;
    end 
  end


  always @(posedge clk) begin
    if(N758) begin
      T608[2] <= N761;
    end 
  end


  always @(posedge clk) begin
    if(N758) begin
      T608[1] <= N760;
    end 
  end


  always @(posedge clk) begin
    if(N758) begin
      T608[0] <= N759;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[63] <= N825;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[62] <= N824;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[61] <= N823;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[60] <= N822;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[59] <= N821;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[58] <= N820;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[57] <= N819;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[56] <= N818;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[55] <= N817;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[54] <= N816;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[53] <= N815;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[52] <= N814;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[51] <= N813;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[50] <= N812;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[49] <= N811;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[48] <= N810;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[47] <= N809;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[46] <= N808;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[45] <= N807;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[44] <= N806;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[43] <= N805;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[42] <= N804;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[41] <= N803;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[40] <= N802;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[39] <= N801;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[38] <= N800;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[37] <= N799;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[36] <= N798;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[35] <= N797;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[34] <= N796;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[33] <= N795;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[32] <= N794;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[31] <= N793;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[30] <= N792;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[29] <= N791;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[28] <= N790;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[27] <= N789;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[26] <= N788;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[25] <= N787;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[24] <= N786;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[23] <= N785;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[22] <= N784;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[21] <= N783;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[20] <= N782;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[19] <= N781;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[18] <= N780;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[17] <= N779;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[16] <= N778;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[15] <= N777;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[14] <= N776;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[13] <= N775;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[12] <= N774;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[11] <= N773;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[10] <= N772;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[9] <= N771;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[8] <= N770;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[7] <= N769;
    end 
  end


  always @(posedge clk) begin
    if(N767) begin
      T608[6] <= N768;
    end 
  end


  always @(posedge clk) begin
    if(N828) begin
      T621[5] <= N834;
    end 
  end


  always @(posedge clk) begin
    if(N828) begin
      T621[4] <= N833;
    end 
  end


  always @(posedge clk) begin
    if(N828) begin
      T621[3] <= N832;
    end 
  end


  always @(posedge clk) begin
    if(N828) begin
      T621[2] <= N831;
    end 
  end


  always @(posedge clk) begin
    if(N828) begin
      T621[1] <= N830;
    end 
  end


  always @(posedge clk) begin
    if(N828) begin
      T621[0] <= N829;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[63] <= N895;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[62] <= N894;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[61] <= N893;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[60] <= N892;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[59] <= N891;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[58] <= N890;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[57] <= N889;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[56] <= N888;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[55] <= N887;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[54] <= N886;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[53] <= N885;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[52] <= N884;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[51] <= N883;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[50] <= N882;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[49] <= N881;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[48] <= N880;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[47] <= N879;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[46] <= N878;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[45] <= N877;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[44] <= N876;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[43] <= N875;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[42] <= N874;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[41] <= N873;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[40] <= N872;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[39] <= N871;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[38] <= N870;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[37] <= N869;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[36] <= N868;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[35] <= N867;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[34] <= N866;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[33] <= N865;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[32] <= N864;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[31] <= N863;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[30] <= N862;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[29] <= N861;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[28] <= N860;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[27] <= N859;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[26] <= N858;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[25] <= N857;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[24] <= N856;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[23] <= N855;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[22] <= N854;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[21] <= N853;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[20] <= N852;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[19] <= N851;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[18] <= N850;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[17] <= N849;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[16] <= N848;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[15] <= N847;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[14] <= N846;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[13] <= N845;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[12] <= N844;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[11] <= N843;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[10] <= N842;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[9] <= N841;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[8] <= N840;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[7] <= N839;
    end 
  end


  always @(posedge clk) begin
    if(N837) begin
      T621[6] <= N838;
    end 
  end


  always @(posedge clk) begin
    if(N898) begin
      T634[5] <= N904;
    end 
  end


  always @(posedge clk) begin
    if(N898) begin
      T634[4] <= N903;
    end 
  end


  always @(posedge clk) begin
    if(N898) begin
      T634[3] <= N902;
    end 
  end


  always @(posedge clk) begin
    if(N898) begin
      T634[2] <= N901;
    end 
  end


  always @(posedge clk) begin
    if(N898) begin
      T634[1] <= N900;
    end 
  end


  always @(posedge clk) begin
    if(N898) begin
      T634[0] <= N899;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[63] <= N965;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[62] <= N964;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[61] <= N963;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[60] <= N962;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[59] <= N961;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[58] <= N960;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[57] <= N959;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[56] <= N958;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[55] <= N957;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[54] <= N956;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[53] <= N955;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[52] <= N954;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[51] <= N953;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[50] <= N952;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[49] <= N951;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[48] <= N950;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[47] <= N949;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[46] <= N948;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[45] <= N947;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[44] <= N946;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[43] <= N945;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[42] <= N944;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[41] <= N943;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[40] <= N942;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[39] <= N941;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[38] <= N940;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[37] <= N939;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[36] <= N938;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[35] <= N937;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[34] <= N936;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[33] <= N935;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[32] <= N934;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[31] <= N933;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[30] <= N932;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[29] <= N931;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[28] <= N930;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[27] <= N929;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[26] <= N928;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[25] <= N927;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[24] <= N926;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[23] <= N925;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[22] <= N924;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[21] <= N923;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[20] <= N922;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[19] <= N921;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[18] <= N920;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[17] <= N919;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[16] <= N918;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[15] <= N917;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[14] <= N916;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[13] <= N915;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[12] <= N914;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[11] <= N913;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[10] <= N912;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[9] <= N911;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[8] <= N910;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[7] <= N909;
    end 
  end


  always @(posedge clk) begin
    if(N907) begin
      T634[6] <= N908;
    end 
  end


  always @(posedge clk) begin
    if(N968) begin
      T647[5] <= N974;
    end 
  end


  always @(posedge clk) begin
    if(N968) begin
      T647[4] <= N973;
    end 
  end


  always @(posedge clk) begin
    if(N968) begin
      T647[3] <= N972;
    end 
  end


  always @(posedge clk) begin
    if(N968) begin
      T647[2] <= N971;
    end 
  end


  always @(posedge clk) begin
    if(N968) begin
      T647[1] <= N970;
    end 
  end


  always @(posedge clk) begin
    if(N968) begin
      T647[0] <= N969;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[63] <= N1035;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[62] <= N1034;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[61] <= N1033;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[60] <= N1032;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[59] <= N1031;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[58] <= N1030;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[57] <= N1029;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[56] <= N1028;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[55] <= N1027;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[54] <= N1026;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[53] <= N1025;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[52] <= N1024;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[51] <= N1023;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[50] <= N1022;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[49] <= N1021;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[48] <= N1020;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[47] <= N1019;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[46] <= N1018;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[45] <= N1017;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[44] <= N1016;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[43] <= N1015;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[42] <= N1014;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[41] <= N1013;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[40] <= N1012;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[39] <= N1011;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[38] <= N1010;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[37] <= N1009;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[36] <= N1008;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[35] <= N1007;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[34] <= N1006;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[33] <= N1005;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[32] <= N1004;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[31] <= N1003;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[30] <= N1002;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[29] <= N1001;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[28] <= N1000;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[27] <= N999;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[26] <= N998;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[25] <= N997;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[24] <= N996;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[23] <= N995;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[22] <= N994;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[21] <= N993;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[20] <= N992;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[19] <= N991;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[18] <= N990;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[17] <= N989;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[16] <= N988;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[15] <= N987;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[14] <= N986;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[13] <= N985;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[12] <= N984;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[11] <= N983;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[10] <= N982;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[9] <= N981;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[8] <= N980;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[7] <= N979;
    end 
  end


  always @(posedge clk) begin
    if(N977) begin
      T647[6] <= N978;
    end 
  end


  always @(posedge clk) begin
    if(N1038) begin
      T660[5] <= N1044;
    end 
  end


  always @(posedge clk) begin
    if(N1038) begin
      T660[4] <= N1043;
    end 
  end


  always @(posedge clk) begin
    if(N1038) begin
      T660[3] <= N1042;
    end 
  end


  always @(posedge clk) begin
    if(N1038) begin
      T660[2] <= N1041;
    end 
  end


  always @(posedge clk) begin
    if(N1038) begin
      T660[1] <= N1040;
    end 
  end


  always @(posedge clk) begin
    if(N1038) begin
      T660[0] <= N1039;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[63] <= N1105;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[62] <= N1104;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[61] <= N1103;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[60] <= N1102;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[59] <= N1101;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[58] <= N1100;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[57] <= N1099;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[56] <= N1098;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[55] <= N1097;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[54] <= N1096;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[53] <= N1095;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[52] <= N1094;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[51] <= N1093;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[50] <= N1092;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[49] <= N1091;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[48] <= N1090;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[47] <= N1089;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[46] <= N1088;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[45] <= N1087;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[44] <= N1086;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[43] <= N1085;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[42] <= N1084;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[41] <= N1083;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[40] <= N1082;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[39] <= N1081;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[38] <= N1080;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[37] <= N1079;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[36] <= N1078;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[35] <= N1077;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[34] <= N1076;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[33] <= N1075;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[32] <= N1074;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[31] <= N1073;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[30] <= N1072;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[29] <= N1071;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[28] <= N1070;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[27] <= N1069;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[26] <= N1068;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[25] <= N1067;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[24] <= N1066;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[23] <= N1065;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[22] <= N1064;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[21] <= N1063;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[20] <= N1062;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[19] <= N1061;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[18] <= N1060;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[17] <= N1059;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[16] <= N1058;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[15] <= N1057;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[14] <= N1056;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[13] <= N1055;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[12] <= N1054;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[11] <= N1053;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[10] <= N1052;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[9] <= N1051;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[8] <= N1050;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[7] <= N1049;
    end 
  end


  always @(posedge clk) begin
    if(N1047) begin
      T660[6] <= N1048;
    end 
  end


  always @(posedge clk) begin
    if(N1108) begin
      T673[5] <= N1114;
    end 
  end


  always @(posedge clk) begin
    if(N1108) begin
      T673[4] <= N1113;
    end 
  end


  always @(posedge clk) begin
    if(N1108) begin
      T673[3] <= N1112;
    end 
  end


  always @(posedge clk) begin
    if(N1108) begin
      T673[2] <= N1111;
    end 
  end


  always @(posedge clk) begin
    if(N1108) begin
      T673[1] <= N1110;
    end 
  end


  always @(posedge clk) begin
    if(N1108) begin
      T673[0] <= N1109;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[63] <= N1175;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[62] <= N1174;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[61] <= N1173;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[60] <= N1172;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[59] <= N1171;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[58] <= N1170;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[57] <= N1169;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[56] <= N1168;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[55] <= N1167;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[54] <= N1166;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[53] <= N1165;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[52] <= N1164;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[51] <= N1163;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[50] <= N1162;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[49] <= N1161;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[48] <= N1160;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[47] <= N1159;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[46] <= N1158;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[45] <= N1157;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[44] <= N1156;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[43] <= N1155;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[42] <= N1154;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[41] <= N1153;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[40] <= N1152;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[39] <= N1151;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[38] <= N1150;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[37] <= N1149;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[36] <= N1148;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[35] <= N1147;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[34] <= N1146;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[33] <= N1145;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[32] <= N1144;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[31] <= N1143;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[30] <= N1142;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[29] <= N1141;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[28] <= N1140;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[27] <= N1139;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[26] <= N1138;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[25] <= N1137;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[24] <= N1136;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[23] <= N1135;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[22] <= N1134;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[21] <= N1133;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[20] <= N1132;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[19] <= N1131;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[18] <= N1130;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[17] <= N1129;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[16] <= N1128;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[15] <= N1127;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[14] <= N1126;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[13] <= N1125;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[12] <= N1124;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[11] <= N1123;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[10] <= N1122;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[9] <= N1121;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[8] <= N1120;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[7] <= N1119;
    end 
  end


  always @(posedge clk) begin
    if(N1117) begin
      T673[6] <= N1118;
    end 
  end


  always @(posedge clk) begin
    if(N1178) begin
      T686[5] <= N1184;
    end 
  end


  always @(posedge clk) begin
    if(N1178) begin
      T686[4] <= N1183;
    end 
  end


  always @(posedge clk) begin
    if(N1178) begin
      T686[3] <= N1182;
    end 
  end


  always @(posedge clk) begin
    if(N1178) begin
      T686[2] <= N1181;
    end 
  end


  always @(posedge clk) begin
    if(N1178) begin
      T686[1] <= N1180;
    end 
  end


  always @(posedge clk) begin
    if(N1178) begin
      T686[0] <= N1179;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[63] <= N1245;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[62] <= N1244;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[61] <= N1243;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[60] <= N1242;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[59] <= N1241;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[58] <= N1240;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[57] <= N1239;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[56] <= N1238;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[55] <= N1237;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[54] <= N1236;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[53] <= N1235;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[52] <= N1234;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[51] <= N1233;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[50] <= N1232;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[49] <= N1231;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[48] <= N1230;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[47] <= N1229;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[46] <= N1228;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[45] <= N1227;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[44] <= N1226;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[43] <= N1225;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[42] <= N1224;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[41] <= N1223;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[40] <= N1222;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[39] <= N1221;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[38] <= N1220;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[37] <= N1219;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[36] <= N1218;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[35] <= N1217;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[34] <= N1216;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[33] <= N1215;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[32] <= N1214;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[31] <= N1213;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[30] <= N1212;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[29] <= N1211;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[28] <= N1210;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[27] <= N1209;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[26] <= N1208;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[25] <= N1207;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[24] <= N1206;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[23] <= N1205;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[22] <= N1204;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[21] <= N1203;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[20] <= N1202;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[19] <= N1201;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[18] <= N1200;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[17] <= N1199;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[16] <= N1198;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[15] <= N1197;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[14] <= N1196;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[13] <= N1195;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[12] <= N1194;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[11] <= N1193;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[10] <= N1192;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[9] <= N1191;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[8] <= N1190;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[7] <= N1189;
    end 
  end


  always @(posedge clk) begin
    if(N1187) begin
      T686[6] <= N1188;
    end 
  end


  always @(posedge clk) begin
    if(N1248) begin
      T699[5] <= N1254;
    end 
  end


  always @(posedge clk) begin
    if(N1248) begin
      T699[4] <= N1253;
    end 
  end


  always @(posedge clk) begin
    if(N1248) begin
      T699[3] <= N1252;
    end 
  end


  always @(posedge clk) begin
    if(N1248) begin
      T699[2] <= N1251;
    end 
  end


  always @(posedge clk) begin
    if(N1248) begin
      T699[1] <= N1250;
    end 
  end


  always @(posedge clk) begin
    if(N1248) begin
      T699[0] <= N1249;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[63] <= N1315;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[62] <= N1314;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[61] <= N1313;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[60] <= N1312;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[59] <= N1311;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[58] <= N1310;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[57] <= N1309;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[56] <= N1308;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[55] <= N1307;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[54] <= N1306;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[53] <= N1305;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[52] <= N1304;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[51] <= N1303;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[50] <= N1302;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[49] <= N1301;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[48] <= N1300;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[47] <= N1299;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[46] <= N1298;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[45] <= N1297;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[44] <= N1296;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[43] <= N1295;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[42] <= N1294;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[41] <= N1293;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[40] <= N1292;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[39] <= N1291;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[38] <= N1290;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[37] <= N1289;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[36] <= N1288;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[35] <= N1287;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[34] <= N1286;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[33] <= N1285;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[32] <= N1284;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[31] <= N1283;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[30] <= N1282;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[29] <= N1281;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[28] <= N1280;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[27] <= N1279;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[26] <= N1278;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[25] <= N1277;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[24] <= N1276;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[23] <= N1275;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[22] <= N1274;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[21] <= N1273;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[20] <= N1272;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[19] <= N1271;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[18] <= N1270;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[17] <= N1269;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[16] <= N1268;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[15] <= N1267;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[14] <= N1266;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[13] <= N1265;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[12] <= N1264;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[11] <= N1263;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[10] <= N1262;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[9] <= N1261;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[8] <= N1260;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[7] <= N1259;
    end 
  end


  always @(posedge clk) begin
    if(N1257) begin
      T699[6] <= N1258;
    end 
  end


  always @(posedge clk) begin
    if(N1318) begin
      T712[5] <= N1324;
    end 
  end


  always @(posedge clk) begin
    if(N1318) begin
      T712[4] <= N1323;
    end 
  end


  always @(posedge clk) begin
    if(N1318) begin
      T712[3] <= N1322;
    end 
  end


  always @(posedge clk) begin
    if(N1318) begin
      T712[2] <= N1321;
    end 
  end


  always @(posedge clk) begin
    if(N1318) begin
      T712[1] <= N1320;
    end 
  end


  always @(posedge clk) begin
    if(N1318) begin
      T712[0] <= N1319;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[63] <= N1385;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[62] <= N1384;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[61] <= N1383;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[60] <= N1382;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[59] <= N1381;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[58] <= N1380;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[57] <= N1379;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[56] <= N1378;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[55] <= N1377;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[54] <= N1376;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[53] <= N1375;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[52] <= N1374;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[51] <= N1373;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[50] <= N1372;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[49] <= N1371;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[48] <= N1370;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[47] <= N1369;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[46] <= N1368;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[45] <= N1367;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[44] <= N1366;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[43] <= N1365;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[42] <= N1364;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[41] <= N1363;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[40] <= N1362;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[39] <= N1361;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[38] <= N1360;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[37] <= N1359;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[36] <= N1358;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[35] <= N1357;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[34] <= N1356;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[33] <= N1355;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[32] <= N1354;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[31] <= N1353;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[30] <= N1352;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[29] <= N1351;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[28] <= N1350;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[27] <= N1349;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[26] <= N1348;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[25] <= N1347;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[24] <= N1346;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[23] <= N1345;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[22] <= N1344;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[21] <= N1343;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[20] <= N1342;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[19] <= N1341;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[18] <= N1340;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[17] <= N1339;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[16] <= N1338;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[15] <= N1337;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[14] <= N1336;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[13] <= N1335;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[12] <= N1334;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[11] <= N1333;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[10] <= N1332;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[9] <= N1331;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[8] <= N1330;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[7] <= N1329;
    end 
  end


  always @(posedge clk) begin
    if(N1327) begin
      T712[6] <= N1328;
    end 
  end


  always @(posedge clk) begin
    if(N1388) begin
      T725[5] <= N1394;
    end 
  end


  always @(posedge clk) begin
    if(N1388) begin
      T725[4] <= N1393;
    end 
  end


  always @(posedge clk) begin
    if(N1388) begin
      T725[3] <= N1392;
    end 
  end


  always @(posedge clk) begin
    if(N1388) begin
      T725[2] <= N1391;
    end 
  end


  always @(posedge clk) begin
    if(N1388) begin
      T725[1] <= N1390;
    end 
  end


  always @(posedge clk) begin
    if(N1388) begin
      T725[0] <= N1389;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[63] <= N1455;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[62] <= N1454;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[61] <= N1453;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[60] <= N1452;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[59] <= N1451;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[58] <= N1450;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[57] <= N1449;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[56] <= N1448;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[55] <= N1447;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[54] <= N1446;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[53] <= N1445;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[52] <= N1444;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[51] <= N1443;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[50] <= N1442;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[49] <= N1441;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[48] <= N1440;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[47] <= N1439;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[46] <= N1438;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[45] <= N1437;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[44] <= N1436;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[43] <= N1435;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[42] <= N1434;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[41] <= N1433;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[40] <= N1432;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[39] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[38] <= N1430;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[37] <= N1429;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[36] <= N1428;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[35] <= N1427;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[34] <= N1426;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[33] <= N1425;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[32] <= N1424;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[31] <= N1423;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[30] <= N1422;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[29] <= N1421;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[28] <= N1420;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[27] <= N1419;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[26] <= N1418;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[25] <= N1417;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[24] <= N1416;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[23] <= N1415;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[22] <= N1414;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[21] <= N1413;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[20] <= N1412;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[19] <= N1411;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[18] <= N1410;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[17] <= N1409;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[16] <= N1408;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[15] <= N1407;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[14] <= N1406;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[13] <= N1405;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[12] <= N1404;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[11] <= N1403;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[10] <= N1402;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[9] <= N1401;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[8] <= N1400;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[7] <= N1399;
    end 
  end


  always @(posedge clk) begin
    if(N1397) begin
      T725[6] <= N1398;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T738[5] <= N1464;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T738[4] <= N1463;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T738[3] <= N1462;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T738[2] <= N1461;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T738[1] <= N1460;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T738[0] <= N1459;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[63] <= N1525;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[62] <= N1524;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[61] <= N1523;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[60] <= N1522;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[59] <= N1521;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[58] <= N1520;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[57] <= N1519;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[56] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[55] <= N1517;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[54] <= N1516;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[53] <= N1515;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[52] <= N1514;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[51] <= N1513;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[50] <= N1512;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[49] <= N1511;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[48] <= N1510;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[47] <= N1509;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[46] <= N1508;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[45] <= N1507;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[44] <= N1506;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[43] <= N1505;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[42] <= N1504;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[41] <= N1503;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[40] <= N1502;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[39] <= N1501;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[38] <= N1500;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[37] <= N1499;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[36] <= N1498;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[35] <= N1497;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[34] <= N1496;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[33] <= N1495;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[32] <= N1494;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[31] <= N1493;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[30] <= N1492;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[29] <= N1491;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[28] <= N1490;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[27] <= N1489;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[26] <= N1488;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[25] <= N1487;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[24] <= N1486;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[23] <= N1485;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[22] <= N1484;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[21] <= N1483;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[20] <= N1482;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[19] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[18] <= N1480;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[17] <= N1479;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[16] <= N1478;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[15] <= N1477;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[14] <= N1476;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[13] <= N1475;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[12] <= N1474;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[11] <= N1473;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[10] <= N1472;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[9] <= N1471;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[8] <= N1470;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[7] <= N1469;
    end 
  end


  always @(posedge clk) begin
    if(N1467) begin
      T738[6] <= N1468;
    end 
  end


  always @(posedge clk) begin
    if(N1528) begin
      T751[5] <= N1534;
    end 
  end


  always @(posedge clk) begin
    if(N1528) begin
      T751[4] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1528) begin
      T751[3] <= N1532;
    end 
  end


  always @(posedge clk) begin
    if(N1528) begin
      T751[2] <= N1531;
    end 
  end


  always @(posedge clk) begin
    if(N1528) begin
      T751[1] <= N1530;
    end 
  end


  always @(posedge clk) begin
    if(N1528) begin
      T751[0] <= N1529;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[63] <= N1595;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[62] <= N1594;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[61] <= N1593;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[60] <= N1592;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[59] <= N1591;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[58] <= N1590;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[57] <= N1589;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[56] <= N1588;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[55] <= N1587;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[54] <= N1586;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[53] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[52] <= N1584;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[51] <= N1583;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[50] <= N1582;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[49] <= N1581;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[48] <= N1580;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[47] <= N1579;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[46] <= N1578;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[45] <= N1577;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[44] <= N1576;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[43] <= N1575;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[42] <= N1574;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[41] <= N1573;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[40] <= N1572;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[39] <= N1571;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[38] <= N1570;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[37] <= N1569;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[36] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[35] <= N1567;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[34] <= N1566;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[33] <= N1565;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[32] <= N1564;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[31] <= N1563;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[30] <= N1562;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[29] <= N1561;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[28] <= N1560;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[27] <= N1559;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[26] <= N1558;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[25] <= N1557;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[24] <= N1556;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[23] <= N1555;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[22] <= N1554;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[21] <= N1553;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[20] <= N1552;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[19] <= N1551;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[18] <= N1550;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[17] <= N1549;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[16] <= N1548;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[15] <= N1547;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[14] <= N1546;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[13] <= N1545;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[12] <= N1544;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[11] <= N1543;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[10] <= N1542;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[9] <= N1541;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[8] <= N1540;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[7] <= N1539;
    end 
  end


  always @(posedge clk) begin
    if(N1537) begin
      T751[6] <= N1538;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T764[5] <= N1604;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T764[4] <= N1603;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T764[3] <= N1602;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T764[2] <= N1601;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T764[1] <= N1600;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T764[0] <= N1599;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[63] <= N1665;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[62] <= N1664;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[61] <= N1663;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[60] <= N1662;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[59] <= N1661;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[58] <= N1660;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[57] <= N1659;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[56] <= N1658;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[55] <= N1657;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[54] <= N1656;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[53] <= N1655;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[52] <= N1654;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[51] <= N1653;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[50] <= N1652;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[49] <= N1651;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[48] <= N1650;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[47] <= N1649;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[46] <= N1648;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[45] <= N1647;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[44] <= N1646;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[43] <= N1645;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[42] <= N1644;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[41] <= N1643;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[40] <= N1642;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[39] <= N1641;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[38] <= N1640;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[37] <= N1639;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[36] <= N1638;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[35] <= N1637;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[34] <= N1636;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[33] <= N1635;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[32] <= N1634;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[31] <= N1633;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[30] <= N1632;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[29] <= N1631;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[28] <= N1630;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[27] <= N1629;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[26] <= N1628;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[25] <= N1627;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[24] <= N1626;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[23] <= N1625;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[22] <= N1624;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[21] <= N1623;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[20] <= N1622;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[19] <= N1621;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[18] <= N1620;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[17] <= N1619;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[16] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[15] <= N1617;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[14] <= N1616;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[13] <= N1615;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[12] <= N1614;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[11] <= N1613;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[10] <= N1612;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[9] <= N1611;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[8] <= N1610;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[7] <= N1609;
    end 
  end


  always @(posedge clk) begin
    if(N1607) begin
      T764[6] <= N1608;
    end 
  end


  always @(posedge clk) begin
    if(N1668) begin
      T777[5] <= N1674;
    end 
  end


  always @(posedge clk) begin
    if(N1668) begin
      T777[4] <= N1673;
    end 
  end


  always @(posedge clk) begin
    if(N1668) begin
      T777[3] <= N1672;
    end 
  end


  always @(posedge clk) begin
    if(N1668) begin
      T777[2] <= N1671;
    end 
  end


  always @(posedge clk) begin
    if(N1668) begin
      T777[1] <= N1670;
    end 
  end


  always @(posedge clk) begin
    if(N1668) begin
      T777[0] <= N1669;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[63] <= N1735;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[62] <= N1734;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[61] <= N1733;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[60] <= N1732;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[59] <= N1731;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[58] <= N1730;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[57] <= N1729;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[56] <= N1728;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[55] <= N1727;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[54] <= N1726;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[53] <= N1725;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[52] <= N1724;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[51] <= N1723;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[50] <= N1722;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[49] <= N1721;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[48] <= N1720;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[47] <= N1719;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[46] <= N1718;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[45] <= N1717;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[44] <= N1716;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[43] <= N1715;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[42] <= N1714;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[41] <= N1713;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[40] <= N1712;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[39] <= N1711;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[38] <= N1710;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[37] <= N1709;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[36] <= N1708;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[35] <= N1707;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[34] <= N1706;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[33] <= N1705;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[32] <= N1704;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[31] <= N1703;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[30] <= N1702;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[29] <= N1701;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[28] <= N1700;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[27] <= N1699;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[26] <= N1698;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[25] <= N1697;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[24] <= N1696;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[23] <= N1695;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[22] <= N1694;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[21] <= N1693;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[20] <= N1692;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[19] <= N1691;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[18] <= N1690;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[17] <= N1689;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[16] <= N1688;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[15] <= N1687;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[14] <= N1686;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[13] <= N1685;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[12] <= N1684;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[11] <= N1683;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[10] <= N1682;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[9] <= N1681;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[8] <= N1680;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[7] <= N1679;
    end 
  end


  always @(posedge clk) begin
    if(N1677) begin
      T777[6] <= N1678;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T790[5] <= N1745;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T790[4] <= N1744;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T790[3] <= N1743;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T790[2] <= N1742;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T790[1] <= N1741;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T790[0] <= N1740;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[63] <= N1807;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[62] <= N1806;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[61] <= N1805;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[60] <= N1804;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[59] <= N1803;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[58] <= N1802;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[57] <= N1801;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[56] <= N1800;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[55] <= N1799;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[54] <= N1798;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[53] <= N1797;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[52] <= N1796;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[51] <= N1795;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[50] <= N1794;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[49] <= N1793;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[48] <= N1792;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[47] <= N1791;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[46] <= N1790;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[45] <= N1789;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[44] <= N1788;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[43] <= N1787;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[42] <= N1786;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[41] <= N1785;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[40] <= N1784;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[39] <= N1783;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[38] <= N1782;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[37] <= N1781;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[36] <= N1780;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[35] <= N1779;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[34] <= N1778;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[33] <= N1777;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[32] <= N1776;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[31] <= N1775;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[30] <= N1774;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[29] <= N1773;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[28] <= N1772;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[27] <= N1771;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[26] <= N1770;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[25] <= N1769;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[24] <= N1768;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[23] <= N1767;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[22] <= N1766;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[21] <= N1765;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[20] <= N1764;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[19] <= N1763;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[18] <= N1762;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[17] <= N1761;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[16] <= N1760;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[15] <= N1759;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[14] <= N1758;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[13] <= N1757;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[12] <= N1756;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[11] <= N1755;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[10] <= N1754;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[9] <= N1753;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[8] <= N1752;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[7] <= N1751;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T790[6] <= N1750;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[63] <= N1875;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[62] <= N1874;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[61] <= N1873;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[60] <= N1872;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[59] <= N1871;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[58] <= N1870;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[57] <= N1869;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[56] <= N1868;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[55] <= N1867;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[54] <= N1866;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[53] <= N1865;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[52] <= N1864;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[51] <= N1863;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[50] <= N1862;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[49] <= N1861;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[48] <= N1860;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[47] <= N1859;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[46] <= N1858;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[45] <= N1857;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[44] <= N1856;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[43] <= N1855;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[42] <= N1854;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[41] <= N1853;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[40] <= N1852;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[39] <= N1851;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[38] <= N1850;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[37] <= N1849;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[36] <= N1848;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[35] <= N1847;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[34] <= N1846;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[33] <= N1845;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[32] <= N1844;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[31] <= N1843;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[30] <= N1842;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[29] <= N1841;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[28] <= N1840;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[27] <= N1839;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[26] <= N1838;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[25] <= N1837;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[24] <= N1836;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[23] <= N1835;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[22] <= N1834;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[21] <= N1833;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[20] <= N1832;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[19] <= N1831;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[18] <= N1830;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[17] <= N1829;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[16] <= N1828;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[15] <= N1827;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[14] <= N1826;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[13] <= N1825;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[12] <= N1824;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[11] <= N1823;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[10] <= N1822;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[9] <= N1821;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[8] <= N1820;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[7] <= N1819;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[6] <= N1818;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[5] <= N1817;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[4] <= N1816;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[3] <= N1815;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[2] <= N1814;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[1] <= N1813;
    end 
  end


  always @(posedge clk) begin
    if(N1811) begin
      reg_tohost[0] <= N1812;
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      io_host_debug_stats_csr <= N1879;
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[63] <= io_rocc_csr_wdata[63];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[62] <= io_rocc_csr_wdata[62];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[61] <= io_rocc_csr_wdata[61];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[60] <= io_rocc_csr_wdata[60];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[59] <= io_rocc_csr_wdata[59];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[58] <= io_rocc_csr_wdata[58];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[57] <= io_rocc_csr_wdata[57];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[56] <= io_rocc_csr_wdata[56];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[55] <= io_rocc_csr_wdata[55];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[54] <= io_rocc_csr_wdata[54];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[53] <= io_rocc_csr_wdata[53];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[52] <= io_rocc_csr_wdata[52];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[51] <= io_rocc_csr_wdata[51];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[50] <= io_rocc_csr_wdata[50];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[49] <= io_rocc_csr_wdata[49];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[48] <= io_rocc_csr_wdata[48];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[47] <= io_rocc_csr_wdata[47];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[46] <= io_rocc_csr_wdata[46];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[45] <= io_rocc_csr_wdata[45];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[44] <= io_rocc_csr_wdata[44];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[43] <= io_rocc_csr_wdata[43];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[42] <= io_rocc_csr_wdata[42];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[41] <= io_rocc_csr_wdata[41];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[40] <= io_rocc_csr_wdata[40];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[39] <= io_rocc_csr_wdata[39];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[38] <= io_rocc_csr_wdata[38];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[37] <= io_rocc_csr_wdata[37];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[36] <= io_rocc_csr_wdata[36];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[35] <= io_rocc_csr_wdata[35];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[34] <= io_rocc_csr_wdata[34];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[33] <= io_rocc_csr_wdata[33];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[32] <= io_rocc_csr_wdata[32];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[31] <= io_rocc_csr_wdata[31];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[30] <= io_rocc_csr_wdata[30];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[29] <= io_rocc_csr_wdata[29];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[28] <= io_rocc_csr_wdata[28];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[27] <= io_rocc_csr_wdata[27];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[26] <= io_rocc_csr_wdata[26];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[25] <= io_rocc_csr_wdata[25];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[24] <= io_rocc_csr_wdata[24];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[23] <= io_rocc_csr_wdata[23];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[22] <= io_rocc_csr_wdata[22];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[21] <= io_rocc_csr_wdata[21];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[20] <= io_rocc_csr_wdata[20];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[19] <= io_rocc_csr_wdata[19];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[18] <= io_rocc_csr_wdata[18];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[17] <= io_rocc_csr_wdata[17];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[16] <= io_rocc_csr_wdata[16];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[15] <= io_rocc_csr_wdata[15];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[14] <= io_rocc_csr_wdata[14];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[13] <= io_rocc_csr_wdata[13];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[12] <= io_rocc_csr_wdata[12];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[11] <= io_rocc_csr_wdata[11];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[10] <= io_rocc_csr_wdata[10];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[9] <= io_rocc_csr_wdata[9];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[8] <= io_rocc_csr_wdata[8];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[7] <= io_rocc_csr_wdata[7];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[6] <= io_rocc_csr_wdata[6];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[5] <= io_rocc_csr_wdata[5];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[4] <= io_rocc_csr_wdata[4];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[3] <= io_rocc_csr_wdata[3];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[2] <= io_rocc_csr_wdata[2];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[1] <= io_rocc_csr_wdata[1];
    end 
  end


  always @(posedge clk) begin
    if(T845) begin
      reg_mscratch[0] <= io_rocc_csr_wdata[0];
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T848_0 <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T848[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T848[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T848_6 <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T858_0 <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T858[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T858[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(reset) begin
      T858_6 <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T894[4] <= T1021[4];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T894[3] <= T1021[3];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T894[2] <= T1021[2];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T894[1] <= T1021[1];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      T894[0] <= T1021[0];
    end 
  end


  always @(posedge clk) begin
    if(T906) begin
      io_host_csr_resp_valid <= 1'b0;
    end else if(1'b1) begin
      io_host_csr_resp_valid <= N1881;
    end 
  end

  assign N2034 = io_rw_wdata[62] & io_rw_wdata[63];
  assign N2035 = io_rw_wdata[61] & N2034;
  assign N2036 = io_rw_wdata[60] & N2035;
  assign N2037 = io_rw_wdata[59] & N2036;
  assign N2038 = io_rw_wdata[58] & N2037;
  assign N2039 = io_rw_wdata[57] & N2038;
  assign N2040 = io_rw_wdata[56] & N2039;
  assign N2041 = io_rw_wdata[55] & N2040;
  assign N2042 = io_rw_wdata[54] & N2041;
  assign N2043 = io_rw_wdata[53] & N2042;
  assign N2044 = io_rw_wdata[52] & N2043;
  assign N2045 = io_rw_wdata[51] & N2044;
  assign N2046 = io_rw_wdata[50] & N2045;
  assign N2047 = io_rw_wdata[49] & N2046;
  assign N2048 = io_rw_wdata[48] & N2047;
  assign N2049 = io_rw_wdata[47] & N2048;
  assign N2050 = io_rw_wdata[46] & N2049;
  assign N2051 = io_rw_wdata[45] & N2050;
  assign N2052 = io_rw_wdata[44] & N2051;
  assign N2053 = io_rw_wdata[43] & N2052;
  assign N2054 = io_rw_wdata[42] & N2053;
  assign N2055 = io_rw_wdata[41] & N2054;
  assign N2056 = io_rw_wdata[40] & N2055;
  assign N2057 = io_rw_wdata[39] & N2056;
  assign N2058 = io_rw_wdata[62] | io_rw_wdata[63];
  assign N2059 = io_rw_wdata[61] | N2058;
  assign N2060 = io_rw_wdata[60] | N2059;
  assign N2061 = io_rw_wdata[59] | N2060;
  assign N2062 = io_rw_wdata[58] | N2061;
  assign N2063 = io_rw_wdata[57] | N2062;
  assign N2064 = io_rw_wdata[56] | N2063;
  assign N2065 = io_rw_wdata[55] | N2064;
  assign N2066 = io_rw_wdata[54] | N2065;
  assign N2067 = io_rw_wdata[53] | N2066;
  assign N2068 = io_rw_wdata[52] | N2067;
  assign N2069 = io_rw_wdata[51] | N2068;
  assign N2070 = io_rw_wdata[50] | N2069;
  assign N2071 = io_rw_wdata[49] | N2070;
  assign N2072 = io_rw_wdata[48] | N2071;
  assign N2073 = io_rw_wdata[47] | N2072;
  assign N2074 = io_rw_wdata[46] | N2073;
  assign N2075 = io_rw_wdata[45] | N2074;
  assign N2076 = io_rw_wdata[44] | N2075;
  assign N2077 = io_rw_wdata[43] | N2076;
  assign N2078 = io_rw_wdata[42] | N2077;
  assign N2079 = io_rw_wdata[41] | N2078;
  assign N2080 = io_rw_wdata[40] | N2079;
  assign N2081 = io_rw_wdata[39] | N2080;
  assign N2082 = io_status_prv[0] & io_status_prv[1];
  assign N2083 = io_rocc_csr_wdata[20] | io_rocc_csr_wdata[21];
  assign N2084 = io_rocc_csr_wdata[19] | N2083;
  assign N2085 = io_rocc_csr_wdata[18] | N2084;
  assign N2086 = io_rocc_csr_wdata[17] | N2085;
  assign N2087 = ~N2086;
  assign N2088 = io_status_prv[0] & io_status_prv[1];
  assign N2089 = reg_fromhost[62] | reg_fromhost[63];
  assign N2090 = reg_fromhost[61] | N2089;
  assign N2091 = reg_fromhost[60] | N2090;
  assign N2092 = reg_fromhost[59] | N2091;
  assign N2093 = reg_fromhost[58] | N2092;
  assign N2094 = reg_fromhost[57] | N2093;
  assign N2095 = reg_fromhost[56] | N2094;
  assign N2096 = reg_fromhost[55] | N2095;
  assign N2097 = reg_fromhost[54] | N2096;
  assign N2098 = reg_fromhost[53] | N2097;
  assign N2099 = reg_fromhost[52] | N2098;
  assign N2100 = reg_fromhost[51] | N2099;
  assign N2101 = reg_fromhost[50] | N2100;
  assign N2102 = reg_fromhost[49] | N2101;
  assign N2103 = reg_fromhost[48] | N2102;
  assign N2104 = reg_fromhost[47] | N2103;
  assign N2105 = reg_fromhost[46] | N2104;
  assign N2106 = reg_fromhost[45] | N2105;
  assign N2107 = reg_fromhost[44] | N2106;
  assign N2108 = reg_fromhost[43] | N2107;
  assign N2109 = reg_fromhost[42] | N2108;
  assign N2110 = reg_fromhost[41] | N2109;
  assign N2111 = reg_fromhost[40] | N2110;
  assign N2112 = reg_fromhost[39] | N2111;
  assign N2113 = reg_fromhost[38] | N2112;
  assign N2114 = reg_fromhost[37] | N2113;
  assign N2115 = reg_fromhost[36] | N2114;
  assign N2116 = reg_fromhost[35] | N2115;
  assign N2117 = reg_fromhost[34] | N2116;
  assign N2118 = reg_fromhost[33] | N2117;
  assign N2119 = reg_fromhost[32] | N2118;
  assign N2120 = reg_fromhost[31] | N2119;
  assign N2121 = reg_fromhost[30] | N2120;
  assign N2122 = reg_fromhost[29] | N2121;
  assign N2123 = reg_fromhost[28] | N2122;
  assign N2124 = reg_fromhost[27] | N2123;
  assign N2125 = reg_fromhost[26] | N2124;
  assign N2126 = reg_fromhost[25] | N2125;
  assign N2127 = reg_fromhost[24] | N2126;
  assign N2128 = reg_fromhost[23] | N2127;
  assign N2129 = reg_fromhost[22] | N2128;
  assign N2130 = reg_fromhost[21] | N2129;
  assign N2131 = reg_fromhost[20] | N2130;
  assign N2132 = reg_fromhost[19] | N2131;
  assign N2133 = reg_fromhost[18] | N2132;
  assign N2134 = reg_fromhost[17] | N2133;
  assign N2135 = reg_fromhost[16] | N2134;
  assign N2136 = reg_fromhost[15] | N2135;
  assign N2137 = reg_fromhost[14] | N2136;
  assign N2138 = reg_fromhost[13] | N2137;
  assign N2139 = reg_fromhost[12] | N2138;
  assign N2140 = reg_fromhost[11] | N2139;
  assign N2141 = reg_fromhost[10] | N2140;
  assign N2142 = reg_fromhost[9] | N2141;
  assign N2143 = reg_fromhost[8] | N2142;
  assign N2144 = reg_fromhost[7] | N2143;
  assign N2145 = reg_fromhost[6] | N2144;
  assign N2146 = reg_fromhost[5] | N2145;
  assign N2147 = reg_fromhost[4] | N2146;
  assign N2148 = reg_fromhost[3] | N2147;
  assign N2149 = reg_fromhost[2] | N2148;
  assign N2150 = reg_fromhost[1] | N2149;
  assign N2151 = reg_fromhost[0] | N2150;
  assign N2152 = ~N2151;
  assign N2153 = ~io_rocc_csr_wdata[20];
  assign N2154 = ~io_rocc_csr_wdata[17];
  assign N2155 = N2153 | io_rocc_csr_wdata[21];
  assign N2156 = io_rocc_csr_wdata[19] | N2155;
  assign N2157 = io_rocc_csr_wdata[18] | N2156;
  assign N2158 = N2154 | N2157;
  assign N2159 = ~N2158;
  assign N2160 = io_status_prv[0] & io_status_prv[1];
  assign N2161 = ~io_cause[2];
  assign N2162 = ~io_cause[1];
  assign N2163 = io_cause[62] | io_cause[63];
  assign N2164 = io_cause[61] | N2163;
  assign N2165 = io_cause[60] | N2164;
  assign N2166 = io_cause[59] | N2165;
  assign N2167 = io_cause[58] | N2166;
  assign N2168 = io_cause[57] | N2167;
  assign N2169 = io_cause[56] | N2168;
  assign N2170 = io_cause[55] | N2169;
  assign N2171 = io_cause[54] | N2170;
  assign N2172 = io_cause[53] | N2171;
  assign N2173 = io_cause[52] | N2172;
  assign N2174 = io_cause[51] | N2173;
  assign N2175 = io_cause[50] | N2174;
  assign N2176 = io_cause[49] | N2175;
  assign N2177 = io_cause[48] | N2176;
  assign N2178 = io_cause[47] | N2177;
  assign N2179 = io_cause[46] | N2178;
  assign N2180 = io_cause[45] | N2179;
  assign N2181 = io_cause[44] | N2180;
  assign N2182 = io_cause[43] | N2181;
  assign N2183 = io_cause[42] | N2182;
  assign N2184 = io_cause[41] | N2183;
  assign N2185 = io_cause[40] | N2184;
  assign N2186 = io_cause[39] | N2185;
  assign N2187 = io_cause[38] | N2186;
  assign N2188 = io_cause[37] | N2187;
  assign N2189 = io_cause[36] | N2188;
  assign N2190 = io_cause[35] | N2189;
  assign N2191 = io_cause[34] | N2190;
  assign N2192 = io_cause[33] | N2191;
  assign N2193 = io_cause[32] | N2192;
  assign N2194 = io_cause[31] | N2193;
  assign N2195 = io_cause[30] | N2194;
  assign N2196 = io_cause[29] | N2195;
  assign N2197 = io_cause[28] | N2196;
  assign N2198 = io_cause[27] | N2197;
  assign N2199 = io_cause[26] | N2198;
  assign N2200 = io_cause[25] | N2199;
  assign N2201 = io_cause[24] | N2200;
  assign N2202 = io_cause[23] | N2201;
  assign N2203 = io_cause[22] | N2202;
  assign N2204 = io_cause[21] | N2203;
  assign N2205 = io_cause[20] | N2204;
  assign N2206 = io_cause[19] | N2205;
  assign N2207 = io_cause[18] | N2206;
  assign N2208 = io_cause[17] | N2207;
  assign N2209 = io_cause[16] | N2208;
  assign N2210 = io_cause[15] | N2209;
  assign N2211 = io_cause[14] | N2210;
  assign N2212 = io_cause[13] | N2211;
  assign N2213 = io_cause[12] | N2212;
  assign N2214 = io_cause[11] | N2213;
  assign N2215 = io_cause[10] | N2214;
  assign N2216 = io_cause[9] | N2215;
  assign N2217 = io_cause[8] | N2216;
  assign N2218 = io_cause[7] | N2217;
  assign N2219 = io_cause[6] | N2218;
  assign N2220 = io_cause[5] | N2219;
  assign N2221 = io_cause[4] | N2220;
  assign N2222 = io_cause[3] | N2221;
  assign N2223 = N2161 | N2222;
  assign N2224 = N2162 | N2223;
  assign N2225 = io_cause[0] | N2224;
  assign N2226 = ~N2225;
  assign N2227 = reg_tohost[62] | reg_tohost[63];
  assign N2228 = reg_tohost[61] | N2227;
  assign N2229 = reg_tohost[60] | N2228;
  assign N2230 = reg_tohost[59] | N2229;
  assign N2231 = reg_tohost[58] | N2230;
  assign N2232 = reg_tohost[57] | N2231;
  assign N2233 = reg_tohost[56] | N2232;
  assign N2234 = reg_tohost[55] | N2233;
  assign N2235 = reg_tohost[54] | N2234;
  assign N2236 = reg_tohost[53] | N2235;
  assign N2237 = reg_tohost[52] | N2236;
  assign N2238 = reg_tohost[51] | N2237;
  assign N2239 = reg_tohost[50] | N2238;
  assign N2240 = reg_tohost[49] | N2239;
  assign N2241 = reg_tohost[48] | N2240;
  assign N2242 = reg_tohost[47] | N2241;
  assign N2243 = reg_tohost[46] | N2242;
  assign N2244 = reg_tohost[45] | N2243;
  assign N2245 = reg_tohost[44] | N2244;
  assign N2246 = reg_tohost[43] | N2245;
  assign N2247 = reg_tohost[42] | N2246;
  assign N2248 = reg_tohost[41] | N2247;
  assign N2249 = reg_tohost[40] | N2248;
  assign N2250 = reg_tohost[39] | N2249;
  assign N2251 = reg_tohost[38] | N2250;
  assign N2252 = reg_tohost[37] | N2251;
  assign N2253 = reg_tohost[36] | N2252;
  assign N2254 = reg_tohost[35] | N2253;
  assign N2255 = reg_tohost[34] | N2254;
  assign N2256 = reg_tohost[33] | N2255;
  assign N2257 = reg_tohost[32] | N2256;
  assign N2258 = reg_tohost[31] | N2257;
  assign N2259 = reg_tohost[30] | N2258;
  assign N2260 = reg_tohost[29] | N2259;
  assign N2261 = reg_tohost[28] | N2260;
  assign N2262 = reg_tohost[27] | N2261;
  assign N2263 = reg_tohost[26] | N2262;
  assign N2264 = reg_tohost[25] | N2263;
  assign N2265 = reg_tohost[24] | N2264;
  assign N2266 = reg_tohost[23] | N2265;
  assign N2267 = reg_tohost[22] | N2266;
  assign N2268 = reg_tohost[21] | N2267;
  assign N2269 = reg_tohost[20] | N2268;
  assign N2270 = reg_tohost[19] | N2269;
  assign N2271 = reg_tohost[18] | N2270;
  assign N2272 = reg_tohost[17] | N2271;
  assign N2273 = reg_tohost[16] | N2272;
  assign N2274 = reg_tohost[15] | N2273;
  assign N2275 = reg_tohost[14] | N2274;
  assign N2276 = reg_tohost[13] | N2275;
  assign N2277 = reg_tohost[12] | N2276;
  assign N2278 = reg_tohost[11] | N2277;
  assign N2279 = reg_tohost[10] | N2278;
  assign N2280 = reg_tohost[9] | N2279;
  assign N2281 = reg_tohost[8] | N2280;
  assign N2282 = reg_tohost[7] | N2281;
  assign N2283 = reg_tohost[6] | N2282;
  assign N2284 = reg_tohost[5] | N2283;
  assign N2285 = reg_tohost[4] | N2284;
  assign N2286 = reg_tohost[3] | N2285;
  assign N2287 = reg_tohost[2] | N2286;
  assign N2288 = reg_tohost[1] | N2287;
  assign N2289 = reg_tohost[0] | N2288;
  assign N2290 = ~N2289;
  assign N2291 = ~io_status_prv[0];
  assign N2292 = N2291 | io_status_prv[1];
  assign N2293 = ~N2292;
  assign N2294 = ~io_rocc_csr_wdata[4];
  assign N2295 = N2294 | io_rocc_csr_wdata[5];
  assign N2296 = ~N2295;
  assign N2297 = ~io_rocc_csr_wdata[7];
  assign N2298 = N2297 | io_rocc_csr_wdata[8];
  assign N2299 = ~N2298;
  assign N2300 = ~io_cause[0];
  assign N2301 = N2300 | N2224;
  assign N2302 = ~N2301;
  assign N2303 = io_status_prv[0] & io_status_prv[1];
  assign N2304 = ~io_rocc_csr_wdata[1];
  assign N2305 = N2304 | io_rocc_csr_wdata[2];
  assign N2306 = ~N2305;
  assign N2307 = io_rocc_csr_wdata[4] & io_rocc_csr_wdata[5];
  assign N2308 = io_rocc_csr_wdata[4] | io_rocc_csr_wdata[5];
  assign N2309 = ~N2308;
  assign N2310 = io_rocc_csr_wdata[7] & io_rocc_csr_wdata[8];
  assign N2311 = io_rocc_csr_wdata[7] | io_rocc_csr_wdata[8];
  assign N2312 = ~N2311;
  assign N2313 = io_cause[1] | N2223;
  assign N2314 = N2300 | N2313;
  assign N2315 = ~N2314;
  assign N2316 = io_cause[0] | N2313;
  assign N2317 = ~N2316;
  assign N2318 = N2291 | io_status_prv[1];
  assign N2319 = ~N2318;
  assign N2320 = io_rocc_csr_wdata[1] & io_rocc_csr_wdata[2];
  assign N2321 = io_rocc_csr_wdata[1] | io_rocc_csr_wdata[2];
  assign N2322 = ~N2321;
  assign N2323 = reg_fromhost[62] | reg_fromhost[63];
  assign N2324 = reg_fromhost[61] | N2323;
  assign N2325 = reg_fromhost[60] | N2324;
  assign N2326 = reg_fromhost[59] | N2325;
  assign N2327 = reg_fromhost[58] | N2326;
  assign N2328 = reg_fromhost[57] | N2327;
  assign N2329 = reg_fromhost[56] | N2328;
  assign N2330 = reg_fromhost[55] | N2329;
  assign N2331 = reg_fromhost[54] | N2330;
  assign N2332 = reg_fromhost[53] | N2331;
  assign N2333 = reg_fromhost[52] | N2332;
  assign N2334 = reg_fromhost[51] | N2333;
  assign N2335 = reg_fromhost[50] | N2334;
  assign N2336 = reg_fromhost[49] | N2335;
  assign N2337 = reg_fromhost[48] | N2336;
  assign N2338 = reg_fromhost[47] | N2337;
  assign N2339 = reg_fromhost[46] | N2338;
  assign N2340 = reg_fromhost[45] | N2339;
  assign N2341 = reg_fromhost[44] | N2340;
  assign N2342 = reg_fromhost[43] | N2341;
  assign N2343 = reg_fromhost[42] | N2342;
  assign N2344 = reg_fromhost[41] | N2343;
  assign N2345 = reg_fromhost[40] | N2344;
  assign N2346 = reg_fromhost[39] | N2345;
  assign N2347 = reg_fromhost[38] | N2346;
  assign N2348 = reg_fromhost[37] | N2347;
  assign N2349 = reg_fromhost[36] | N2348;
  assign N2350 = reg_fromhost[35] | N2349;
  assign N2351 = reg_fromhost[34] | N2350;
  assign N2352 = reg_fromhost[33] | N2351;
  assign N2353 = reg_fromhost[32] | N2352;
  assign N2354 = reg_fromhost[31] | N2353;
  assign N2355 = reg_fromhost[30] | N2354;
  assign N2356 = reg_fromhost[29] | N2355;
  assign N2357 = reg_fromhost[28] | N2356;
  assign N2358 = reg_fromhost[27] | N2357;
  assign N2359 = reg_fromhost[26] | N2358;
  assign N2360 = reg_fromhost[25] | N2359;
  assign N2361 = reg_fromhost[24] | N2360;
  assign N2362 = reg_fromhost[23] | N2361;
  assign N2363 = reg_fromhost[22] | N2362;
  assign N2364 = reg_fromhost[21] | N2363;
  assign N2365 = reg_fromhost[20] | N2364;
  assign N2366 = reg_fromhost[19] | N2365;
  assign N2367 = reg_fromhost[18] | N2366;
  assign N2368 = reg_fromhost[17] | N2367;
  assign N2369 = reg_fromhost[16] | N2368;
  assign N2370 = reg_fromhost[15] | N2369;
  assign N2371 = reg_fromhost[14] | N2370;
  assign N2372 = reg_fromhost[13] | N2371;
  assign N2373 = reg_fromhost[12] | N2372;
  assign N2374 = reg_fromhost[11] | N2373;
  assign N2375 = reg_fromhost[10] | N2374;
  assign N2376 = reg_fromhost[9] | N2375;
  assign N2377 = reg_fromhost[8] | N2376;
  assign N2378 = reg_fromhost[7] | N2377;
  assign N2379 = reg_fromhost[6] | N2378;
  assign N2380 = reg_fromhost[5] | N2379;
  assign N2381 = reg_fromhost[4] | N2380;
  assign N2382 = reg_fromhost[3] | N2381;
  assign N2383 = reg_fromhost[2] | N2382;
  assign N2384 = reg_fromhost[1] | N2383;
  assign N2385 = reg_fromhost[0] | N2384;
  assign N2386 = ~io_rw_cmd[0];
  assign N2387 = io_rw_cmd[1] | io_rw_cmd[2];
  assign N2388 = N2386 | N2387;
  assign N2389 = ~N2388;
  assign N2390 = ~io_rw_cmd[1];
  assign N2391 = N2390 | io_rw_cmd[2];
  assign N2392 = N2386 | N2391;
  assign N2393 = ~N2392;
  assign N2394 = io_rw_addr[10] & io_rw_addr[11];
  assign N2395 = io_rw_cmd[0] | N2391;
  assign N2396 = ~N2395;
  assign N2397 = ~io_rw_cmd[2];
  assign N2398 = io_rw_cmd[1] | N2397;
  assign N2399 = N2386 | N2398;
  assign N2400 = ~io_rocc_csr_waddr[8];
  assign N2401 = ~io_rocc_csr_waddr[0];
  assign N2402 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2403 = io_rocc_csr_waddr[9] | N2402;
  assign N2404 = N2400 | N2403;
  assign N2405 = io_rocc_csr_waddr[7] | N2404;
  assign N2406 = io_rocc_csr_waddr[6] | N2405;
  assign N2407 = io_rocc_csr_waddr[5] | N2406;
  assign N2408 = io_rocc_csr_waddr[4] | N2407;
  assign N2409 = io_rocc_csr_waddr[3] | N2408;
  assign N2410 = io_rocc_csr_waddr[2] | N2409;
  assign N2411 = io_rocc_csr_waddr[1] | N2410;
  assign N2412 = N2401 | N2411;
  assign N2413 = ~N2412;
  assign N2414 = ~io_rocc_csr_waddr[6];
  assign N2415 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2416 = io_rocc_csr_waddr[9] | N2415;
  assign N2417 = N2400 | N2416;
  assign N2418 = io_rocc_csr_waddr[7] | N2417;
  assign N2419 = N2414 | N2418;
  assign N2420 = io_rocc_csr_waddr[5] | N2419;
  assign N2421 = io_rocc_csr_waddr[4] | N2420;
  assign N2422 = io_rocc_csr_waddr[3] | N2421;
  assign N2423 = io_rocc_csr_waddr[2] | N2422;
  assign N2424 = io_rocc_csr_waddr[1] | N2423;
  assign N2425 = N2401 | N2424;
  assign N2426 = ~N2425;
  assign N2427 = ~io_rocc_csr_waddr[7];
  assign N2428 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2429 = io_rocc_csr_waddr[9] | N2428;
  assign N2430 = N2400 | N2429;
  assign N2431 = N2427 | N2430;
  assign N2432 = io_rocc_csr_waddr[6] | N2431;
  assign N2433 = io_rocc_csr_waddr[5] | N2432;
  assign N2434 = io_rocc_csr_waddr[4] | N2433;
  assign N2435 = io_rocc_csr_waddr[3] | N2434;
  assign N2436 = io_rocc_csr_waddr[2] | N2435;
  assign N2437 = io_rocc_csr_waddr[1] | N2436;
  assign N2438 = N2401 | N2437;
  assign N2439 = ~N2438;
  assign N2440 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2441 = io_rocc_csr_waddr[9] | N2440;
  assign N2442 = N2400 | N2441;
  assign N2443 = N2427 | N2442;
  assign N2444 = io_rocc_csr_waddr[6] | N2443;
  assign N2445 = io_rocc_csr_waddr[5] | N2444;
  assign N2446 = io_rocc_csr_waddr[4] | N2445;
  assign N2447 = io_rocc_csr_waddr[3] | N2446;
  assign N2448 = io_rocc_csr_waddr[2] | N2447;
  assign N2449 = io_rocc_csr_waddr[1] | N2448;
  assign N2450 = io_rocc_csr_waddr[0] | N2449;
  assign N2451 = ~N2450;
  assign N2452 = ~io_rocc_csr_waddr[11];
  assign N2453 = ~io_rocc_csr_waddr[10];
  assign N2454 = ~io_rocc_csr_waddr[1];
  assign N2455 = N2453 | N2452;
  assign N2456 = io_rocc_csr_waddr[9] | N2455;
  assign N2457 = N2400 | N2456;
  assign N2458 = io_rocc_csr_waddr[7] | N2457;
  assign N2459 = N2414 | N2458;
  assign N2460 = io_rocc_csr_waddr[5] | N2459;
  assign N2461 = io_rocc_csr_waddr[4] | N2460;
  assign N2462 = io_rocc_csr_waddr[3] | N2461;
  assign N2463 = io_rocc_csr_waddr[2] | N2462;
  assign N2464 = N2454 | N2463;
  assign N2465 = N2401 | N2464;
  assign N2466 = ~N2465;
  assign N2467 = N2453 | N2452;
  assign N2468 = io_rocc_csr_waddr[9] | N2467;
  assign N2469 = N2400 | N2468;
  assign N2470 = io_rocc_csr_waddr[7] | N2469;
  assign N2471 = N2414 | N2470;
  assign N2472 = io_rocc_csr_waddr[5] | N2471;
  assign N2473 = io_rocc_csr_waddr[4] | N2472;
  assign N2474 = io_rocc_csr_waddr[3] | N2473;
  assign N2475 = io_rocc_csr_waddr[2] | N2474;
  assign N2476 = N2454 | N2475;
  assign N2477 = io_rocc_csr_waddr[0] | N2476;
  assign N2478 = ~N2477;
  assign N2479 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2480 = io_rocc_csr_waddr[9] | N2479;
  assign N2481 = N2400 | N2480;
  assign N2482 = io_rocc_csr_waddr[7] | N2481;
  assign N2483 = N2414 | N2482;
  assign N2484 = io_rocc_csr_waddr[5] | N2483;
  assign N2485 = io_rocc_csr_waddr[4] | N2484;
  assign N2486 = io_rocc_csr_waddr[3] | N2485;
  assign N2487 = io_rocc_csr_waddr[2] | N2486;
  assign N2488 = io_rocc_csr_waddr[1] | N2487;
  assign N2489 = io_rocc_csr_waddr[0] | N2488;
  assign N2490 = ~N2489;
  assign N2491 = ~io_rocc_csr_waddr[2];
  assign N2492 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2493 = io_rocc_csr_waddr[9] | N2492;
  assign N2494 = N2400 | N2493;
  assign N2495 = io_rocc_csr_waddr[7] | N2494;
  assign N2496 = io_rocc_csr_waddr[6] | N2495;
  assign N2497 = io_rocc_csr_waddr[5] | N2496;
  assign N2498 = io_rocc_csr_waddr[4] | N2497;
  assign N2499 = io_rocc_csr_waddr[3] | N2498;
  assign N2500 = N2491 | N2499;
  assign N2501 = io_rocc_csr_waddr[1] | N2500;
  assign N2502 = io_rocc_csr_waddr[0] | N2501;
  assign N2503 = ~N2502;
  assign N2504 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2505 = io_rocc_csr_waddr[9] | N2504;
  assign N2506 = N2400 | N2505;
  assign N2507 = io_rocc_csr_waddr[7] | N2506;
  assign N2508 = N2414 | N2507;
  assign N2509 = io_rocc_csr_waddr[5] | N2508;
  assign N2510 = io_rocc_csr_waddr[4] | N2509;
  assign N2511 = io_rocc_csr_waddr[3] | N2510;
  assign N2512 = N2491 | N2511;
  assign N2513 = io_rocc_csr_waddr[1] | N2512;
  assign N2514 = io_rocc_csr_waddr[0] | N2513;
  assign N2515 = ~N2514;
  assign N2516 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2517 = io_rocc_csr_waddr[9] | N2516;
  assign N2518 = N2400 | N2517;
  assign N2519 = io_rocc_csr_waddr[7] | N2518;
  assign N2520 = io_rocc_csr_waddr[6] | N2519;
  assign N2521 = io_rocc_csr_waddr[5] | N2520;
  assign N2522 = io_rocc_csr_waddr[4] | N2521;
  assign N2523 = io_rocc_csr_waddr[3] | N2522;
  assign N2524 = io_rocc_csr_waddr[2] | N2523;
  assign N2525 = io_rocc_csr_waddr[1] | N2524;
  assign N2526 = io_rocc_csr_waddr[0] | N2525;
  assign N2527 = ~N2526;
  assign N2528 = ~io_rocc_csr_waddr[3];
  assign N2529 = N2453 | N2452;
  assign N2530 = io_rocc_csr_waddr[9] | N2529;
  assign N2531 = io_rocc_csr_waddr[8] | N2530;
  assign N2532 = N2427 | N2531;
  assign N2533 = N2414 | N2532;
  assign N2534 = io_rocc_csr_waddr[5] | N2533;
  assign N2535 = io_rocc_csr_waddr[4] | N2534;
  assign N2536 = N2528 | N2535;
  assign N2537 = N2491 | N2536;
  assign N2538 = N2454 | N2537;
  assign N2539 = N2401 | N2538;
  assign N2540 = ~N2539;
  assign N2541 = N2453 | N2452;
  assign N2542 = io_rocc_csr_waddr[9] | N2541;
  assign N2543 = io_rocc_csr_waddr[8] | N2542;
  assign N2544 = N2427 | N2543;
  assign N2545 = N2414 | N2544;
  assign N2546 = io_rocc_csr_waddr[5] | N2545;
  assign N2547 = io_rocc_csr_waddr[4] | N2546;
  assign N2548 = N2528 | N2547;
  assign N2549 = N2491 | N2548;
  assign N2550 = N2454 | N2549;
  assign N2551 = io_rocc_csr_waddr[0] | N2550;
  assign N2552 = ~N2551;
  assign N2553 = N2453 | N2452;
  assign N2554 = io_rocc_csr_waddr[9] | N2553;
  assign N2555 = io_rocc_csr_waddr[8] | N2554;
  assign N2556 = N2427 | N2555;
  assign N2557 = N2414 | N2556;
  assign N2558 = io_rocc_csr_waddr[5] | N2557;
  assign N2559 = io_rocc_csr_waddr[4] | N2558;
  assign N2560 = N2528 | N2559;
  assign N2561 = N2491 | N2560;
  assign N2562 = io_rocc_csr_waddr[1] | N2561;
  assign N2563 = N2401 | N2562;
  assign N2564 = ~N2563;
  assign N2565 = N2453 | N2452;
  assign N2566 = io_rocc_csr_waddr[9] | N2565;
  assign N2567 = io_rocc_csr_waddr[8] | N2566;
  assign N2568 = N2427 | N2567;
  assign N2569 = N2414 | N2568;
  assign N2570 = io_rocc_csr_waddr[5] | N2569;
  assign N2571 = io_rocc_csr_waddr[4] | N2570;
  assign N2572 = N2528 | N2571;
  assign N2573 = N2491 | N2572;
  assign N2574 = io_rocc_csr_waddr[1] | N2573;
  assign N2575 = io_rocc_csr_waddr[0] | N2574;
  assign N2576 = ~N2575;
  assign N2577 = N2453 | N2452;
  assign N2578 = io_rocc_csr_waddr[9] | N2577;
  assign N2579 = io_rocc_csr_waddr[8] | N2578;
  assign N2580 = N2427 | N2579;
  assign N2581 = N2414 | N2580;
  assign N2582 = io_rocc_csr_waddr[5] | N2581;
  assign N2583 = io_rocc_csr_waddr[4] | N2582;
  assign N2584 = N2528 | N2583;
  assign N2585 = io_rocc_csr_waddr[2] | N2584;
  assign N2586 = N2454 | N2585;
  assign N2587 = N2401 | N2586;
  assign N2588 = ~N2587;
  assign N2589 = N2453 | N2452;
  assign N2590 = io_rocc_csr_waddr[9] | N2589;
  assign N2591 = io_rocc_csr_waddr[8] | N2590;
  assign N2592 = N2427 | N2591;
  assign N2593 = N2414 | N2592;
  assign N2594 = io_rocc_csr_waddr[5] | N2593;
  assign N2595 = io_rocc_csr_waddr[4] | N2594;
  assign N2596 = N2528 | N2595;
  assign N2597 = io_rocc_csr_waddr[2] | N2596;
  assign N2598 = N2454 | N2597;
  assign N2599 = io_rocc_csr_waddr[0] | N2598;
  assign N2600 = ~N2599;
  assign N2601 = N2453 | N2452;
  assign N2602 = io_rocc_csr_waddr[9] | N2601;
  assign N2603 = io_rocc_csr_waddr[8] | N2602;
  assign N2604 = N2427 | N2603;
  assign N2605 = N2414 | N2604;
  assign N2606 = io_rocc_csr_waddr[5] | N2605;
  assign N2607 = io_rocc_csr_waddr[4] | N2606;
  assign N2608 = N2528 | N2607;
  assign N2609 = io_rocc_csr_waddr[2] | N2608;
  assign N2610 = io_rocc_csr_waddr[1] | N2609;
  assign N2611 = N2401 | N2610;
  assign N2612 = ~N2611;
  assign N2613 = N2453 | N2452;
  assign N2614 = io_rocc_csr_waddr[9] | N2613;
  assign N2615 = io_rocc_csr_waddr[8] | N2614;
  assign N2616 = N2427 | N2615;
  assign N2617 = N2414 | N2616;
  assign N2618 = io_rocc_csr_waddr[5] | N2617;
  assign N2619 = io_rocc_csr_waddr[4] | N2618;
  assign N2620 = N2528 | N2619;
  assign N2621 = io_rocc_csr_waddr[2] | N2620;
  assign N2622 = io_rocc_csr_waddr[1] | N2621;
  assign N2623 = io_rocc_csr_waddr[0] | N2622;
  assign N2624 = ~N2623;
  assign N2625 = N2453 | N2452;
  assign N2626 = io_rocc_csr_waddr[9] | N2625;
  assign N2627 = io_rocc_csr_waddr[8] | N2626;
  assign N2628 = N2427 | N2627;
  assign N2629 = N2414 | N2628;
  assign N2630 = io_rocc_csr_waddr[5] | N2629;
  assign N2631 = io_rocc_csr_waddr[4] | N2630;
  assign N2632 = io_rocc_csr_waddr[3] | N2631;
  assign N2633 = N2491 | N2632;
  assign N2634 = N2454 | N2633;
  assign N2635 = N2401 | N2634;
  assign N2636 = ~N2635;
  assign N2637 = N2453 | N2452;
  assign N2638 = io_rocc_csr_waddr[9] | N2637;
  assign N2639 = io_rocc_csr_waddr[8] | N2638;
  assign N2640 = N2427 | N2639;
  assign N2641 = N2414 | N2640;
  assign N2642 = io_rocc_csr_waddr[5] | N2641;
  assign N2643 = io_rocc_csr_waddr[4] | N2642;
  assign N2644 = io_rocc_csr_waddr[3] | N2643;
  assign N2645 = N2491 | N2644;
  assign N2646 = N2454 | N2645;
  assign N2647 = io_rocc_csr_waddr[0] | N2646;
  assign N2648 = ~N2647;
  assign N2649 = N2453 | N2452;
  assign N2650 = io_rocc_csr_waddr[9] | N2649;
  assign N2651 = io_rocc_csr_waddr[8] | N2650;
  assign N2652 = N2427 | N2651;
  assign N2653 = N2414 | N2652;
  assign N2654 = io_rocc_csr_waddr[5] | N2653;
  assign N2655 = io_rocc_csr_waddr[4] | N2654;
  assign N2656 = io_rocc_csr_waddr[3] | N2655;
  assign N2657 = N2491 | N2656;
  assign N2658 = io_rocc_csr_waddr[1] | N2657;
  assign N2659 = N2401 | N2658;
  assign N2660 = ~N2659;
  assign N2661 = N2453 | N2452;
  assign N2662 = io_rocc_csr_waddr[9] | N2661;
  assign N2663 = io_rocc_csr_waddr[8] | N2662;
  assign N2664 = N2427 | N2663;
  assign N2665 = N2414 | N2664;
  assign N2666 = io_rocc_csr_waddr[5] | N2665;
  assign N2667 = io_rocc_csr_waddr[4] | N2666;
  assign N2668 = io_rocc_csr_waddr[3] | N2667;
  assign N2669 = N2491 | N2668;
  assign N2670 = io_rocc_csr_waddr[1] | N2669;
  assign N2671 = io_rocc_csr_waddr[0] | N2670;
  assign N2672 = ~N2671;
  assign N2673 = N2453 | N2452;
  assign N2674 = io_rocc_csr_waddr[9] | N2673;
  assign N2675 = io_rocc_csr_waddr[8] | N2674;
  assign N2676 = N2427 | N2675;
  assign N2677 = N2414 | N2676;
  assign N2678 = io_rocc_csr_waddr[5] | N2677;
  assign N2679 = io_rocc_csr_waddr[4] | N2678;
  assign N2680 = io_rocc_csr_waddr[3] | N2679;
  assign N2681 = io_rocc_csr_waddr[2] | N2680;
  assign N2682 = N2454 | N2681;
  assign N2683 = N2401 | N2682;
  assign N2684 = ~N2683;
  assign N2685 = N2453 | N2452;
  assign N2686 = io_rocc_csr_waddr[9] | N2685;
  assign N2687 = io_rocc_csr_waddr[8] | N2686;
  assign N2688 = N2427 | N2687;
  assign N2689 = N2414 | N2688;
  assign N2690 = io_rocc_csr_waddr[5] | N2689;
  assign N2691 = io_rocc_csr_waddr[4] | N2690;
  assign N2692 = io_rocc_csr_waddr[3] | N2691;
  assign N2693 = io_rocc_csr_waddr[2] | N2692;
  assign N2694 = N2454 | N2693;
  assign N2695 = io_rocc_csr_waddr[0] | N2694;
  assign N2696 = ~N2695;
  assign N2697 = N2453 | N2452;
  assign N2698 = io_rocc_csr_waddr[9] | N2697;
  assign N2699 = io_rocc_csr_waddr[8] | N2698;
  assign N2700 = N2427 | N2699;
  assign N2701 = N2414 | N2700;
  assign N2702 = io_rocc_csr_waddr[5] | N2701;
  assign N2703 = io_rocc_csr_waddr[4] | N2702;
  assign N2704 = io_rocc_csr_waddr[3] | N2703;
  assign N2705 = io_rocc_csr_waddr[2] | N2704;
  assign N2706 = io_rocc_csr_waddr[1] | N2705;
  assign N2707 = N2401 | N2706;
  assign N2708 = ~N2707;
  assign N2709 = N2453 | N2452;
  assign N2710 = io_rocc_csr_waddr[9] | N2709;
  assign N2711 = io_rocc_csr_waddr[8] | N2710;
  assign N2712 = N2427 | N2711;
  assign N2713 = N2414 | N2712;
  assign N2714 = io_rocc_csr_waddr[5] | N2713;
  assign N2715 = io_rocc_csr_waddr[4] | N2714;
  assign N2716 = io_rocc_csr_waddr[3] | N2715;
  assign N2717 = io_rocc_csr_waddr[2] | N2716;
  assign N2718 = io_rocc_csr_waddr[1] | N2717;
  assign N2719 = io_rocc_csr_waddr[0] | N2718;
  assign N2720 = ~N2719;
  assign N2721 = io_rocc_csr_waddr[10] | N2452;
  assign N2722 = io_rocc_csr_waddr[9] | N2721;
  assign N2723 = N2400 | N2722;
  assign N2724 = io_rocc_csr_waddr[7] | N2723;
  assign N2725 = io_rocc_csr_waddr[6] | N2724;
  assign N2726 = io_rocc_csr_waddr[5] | N2725;
  assign N2727 = io_rocc_csr_waddr[4] | N2726;
  assign N2728 = io_rocc_csr_waddr[3] | N2727;
  assign N2729 = io_rocc_csr_waddr[2] | N2728;
  assign N2730 = N2454 | N2729;
  assign N2731 = io_rocc_csr_waddr[0] | N2730;
  assign N2732 = ~N2731;
  assign N2733 = N2453 | N2452;
  assign N2734 = io_rocc_csr_waddr[9] | N2733;
  assign N2735 = io_rocc_csr_waddr[8] | N2734;
  assign N2736 = io_rocc_csr_waddr[7] | N2735;
  assign N2737 = io_rocc_csr_waddr[6] | N2736;
  assign N2738 = io_rocc_csr_waddr[5] | N2737;
  assign N2739 = io_rocc_csr_waddr[4] | N2738;
  assign N2740 = io_rocc_csr_waddr[3] | N2739;
  assign N2741 = io_rocc_csr_waddr[2] | N2740;
  assign N2742 = N2454 | N2741;
  assign N2743 = io_rocc_csr_waddr[0] | N2742;
  assign N2744 = ~N2743;
  assign N2745 = ~io_rocc_csr_waddr[9];
  assign N2746 = N2453 | io_rocc_csr_waddr[11];
  assign N2747 = N2745 | N2746;
  assign N2748 = N2400 | N2747;
  assign N2749 = N2427 | N2748;
  assign N2750 = io_rocc_csr_waddr[6] | N2749;
  assign N2751 = io_rocc_csr_waddr[5] | N2750;
  assign N2752 = io_rocc_csr_waddr[4] | N2751;
  assign N2753 = io_rocc_csr_waddr[3] | N2752;
  assign N2754 = io_rocc_csr_waddr[2] | N2753;
  assign N2755 = io_rocc_csr_waddr[1] | N2754;
  assign N2756 = N2401 | N2755;
  assign N2757 = ~N2756;
  assign N2758 = N2453 | io_rocc_csr_waddr[11];
  assign N2759 = N2745 | N2758;
  assign N2760 = N2400 | N2759;
  assign N2761 = N2427 | N2760;
  assign N2762 = io_rocc_csr_waddr[6] | N2761;
  assign N2763 = io_rocc_csr_waddr[5] | N2762;
  assign N2764 = io_rocc_csr_waddr[4] | N2763;
  assign N2765 = io_rocc_csr_waddr[3] | N2764;
  assign N2766 = io_rocc_csr_waddr[2] | N2765;
  assign N2767 = io_rocc_csr_waddr[1] | N2766;
  assign N2768 = io_rocc_csr_waddr[0] | N2767;
  assign N2769 = ~N2768;
  assign N2770 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2771 = io_rocc_csr_waddr[9] | N2770;
  assign N2772 = io_rocc_csr_waddr[8] | N2771;
  assign N2773 = N2427 | N2772;
  assign N2774 = N2414 | N2773;
  assign N2775 = io_rocc_csr_waddr[5] | N2774;
  assign N2776 = io_rocc_csr_waddr[4] | N2775;
  assign N2777 = io_rocc_csr_waddr[3] | N2776;
  assign N2778 = io_rocc_csr_waddr[2] | N2777;
  assign N2779 = io_rocc_csr_waddr[1] | N2778;
  assign N2780 = io_rocc_csr_waddr[0] | N2779;
  assign N2781 = ~N2780;
  assign N2782 = ~io_rocc_csr_waddr[4];
  assign N2783 = N2453 | N2452;
  assign N2784 = N2745 | N2783;
  assign N2785 = N2400 | N2784;
  assign N2786 = io_rocc_csr_waddr[7] | N2785;
  assign N2787 = io_rocc_csr_waddr[6] | N2786;
  assign N2788 = io_rocc_csr_waddr[5] | N2787;
  assign N2789 = N2782 | N2788;
  assign N2790 = io_rocc_csr_waddr[3] | N2789;
  assign N2791 = io_rocc_csr_waddr[2] | N2790;
  assign N2792 = io_rocc_csr_waddr[1] | N2791;
  assign N2793 = io_rocc_csr_waddr[0] | N2792;
  assign N2794 = ~N2793;
  assign N2795 = reg_mstatus_fs[0] | reg_mstatus_fs[1];
  assign N2796 = reg_mstatus_xs[0] | reg_mstatus_xs[1];
  assign N2797 = ~io_rocc_csr_waddr[5];
  assign N2798 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2799 = N2745 | N2798;
  assign N2800 = N2400 | N2799;
  assign N2801 = io_rocc_csr_waddr[7] | N2800;
  assign N2802 = io_rocc_csr_waddr[6] | N2801;
  assign N2803 = N2797 | N2802;
  assign N2804 = io_rocc_csr_waddr[4] | N2803;
  assign N2805 = io_rocc_csr_waddr[3] | N2804;
  assign N2806 = io_rocc_csr_waddr[2] | N2805;
  assign N2807 = io_rocc_csr_waddr[1] | N2806;
  assign N2808 = N2401 | N2807;
  assign N2809 = ~N2808;
  assign N2810 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2811 = N2745 | N2810;
  assign N2812 = N2400 | N2811;
  assign N2813 = io_rocc_csr_waddr[7] | N2812;
  assign N2814 = N2414 | N2813;
  assign N2815 = io_rocc_csr_waddr[5] | N2814;
  assign N2816 = io_rocc_csr_waddr[4] | N2815;
  assign N2817 = io_rocc_csr_waddr[3] | N2816;
  assign N2818 = io_rocc_csr_waddr[2] | N2817;
  assign N2819 = N2454 | N2818;
  assign N2820 = io_rocc_csr_waddr[0] | N2819;
  assign N2821 = ~N2820;
  assign N2822 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2823 = N2745 | N2822;
  assign N2824 = N2400 | N2823;
  assign N2825 = io_rocc_csr_waddr[7] | N2824;
  assign N2826 = N2414 | N2825;
  assign N2827 = io_rocc_csr_waddr[5] | N2826;
  assign N2828 = io_rocc_csr_waddr[4] | N2827;
  assign N2829 = io_rocc_csr_waddr[3] | N2828;
  assign N2830 = io_rocc_csr_waddr[2] | N2829;
  assign N2831 = N2454 | N2830;
  assign N2832 = N2401 | N2831;
  assign N2833 = ~N2832;
  assign N2834 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2835 = N2745 | N2834;
  assign N2836 = N2400 | N2835;
  assign N2837 = io_rocc_csr_waddr[7] | N2836;
  assign N2838 = N2414 | N2837;
  assign N2839 = io_rocc_csr_waddr[5] | N2838;
  assign N2840 = io_rocc_csr_waddr[4] | N2839;
  assign N2841 = io_rocc_csr_waddr[3] | N2840;
  assign N2842 = io_rocc_csr_waddr[2] | N2841;
  assign N2843 = io_rocc_csr_waddr[1] | N2842;
  assign N2844 = N2401 | N2843;
  assign N2845 = ~N2844;
  assign N2846 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2847 = N2745 | N2846;
  assign N2848 = N2400 | N2847;
  assign N2849 = io_rocc_csr_waddr[7] | N2848;
  assign N2850 = N2414 | N2849;
  assign N2851 = io_rocc_csr_waddr[5] | N2850;
  assign N2852 = io_rocc_csr_waddr[4] | N2851;
  assign N2853 = io_rocc_csr_waddr[3] | N2852;
  assign N2854 = io_rocc_csr_waddr[2] | N2853;
  assign N2855 = io_rocc_csr_waddr[1] | N2854;
  assign N2856 = io_rocc_csr_waddr[0] | N2855;
  assign N2857 = ~N2856;
  assign N2858 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2859 = N2745 | N2858;
  assign N2860 = N2400 | N2859;
  assign N2861 = io_rocc_csr_waddr[7] | N2860;
  assign N2862 = io_rocc_csr_waddr[6] | N2861;
  assign N2863 = io_rocc_csr_waddr[5] | N2862;
  assign N2864 = io_rocc_csr_waddr[4] | N2863;
  assign N2865 = io_rocc_csr_waddr[3] | N2864;
  assign N2866 = N2491 | N2865;
  assign N2867 = io_rocc_csr_waddr[1] | N2866;
  assign N2868 = io_rocc_csr_waddr[0] | N2867;
  assign N2869 = ~N2868;
  assign N2870 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2871 = N2745 | N2870;
  assign N2872 = N2400 | N2871;
  assign N2873 = io_rocc_csr_waddr[7] | N2872;
  assign N2874 = N2414 | N2873;
  assign N2875 = io_rocc_csr_waddr[5] | N2874;
  assign N2876 = io_rocc_csr_waddr[4] | N2875;
  assign N2877 = io_rocc_csr_waddr[3] | N2876;
  assign N2878 = N2491 | N2877;
  assign N2879 = io_rocc_csr_waddr[1] | N2878;
  assign N2880 = io_rocc_csr_waddr[0] | N2879;
  assign N2881 = ~N2880;
  assign N2882 = N2453 | io_rocc_csr_waddr[11];
  assign N2883 = N2745 | N2882;
  assign N2884 = N2400 | N2883;
  assign N2885 = N2427 | N2884;
  assign N2886 = io_rocc_csr_waddr[6] | N2885;
  assign N2887 = io_rocc_csr_waddr[5] | N2886;
  assign N2888 = io_rocc_csr_waddr[4] | N2887;
  assign N2889 = io_rocc_csr_waddr[3] | N2888;
  assign N2890 = io_rocc_csr_waddr[2] | N2889;
  assign N2891 = N2454 | N2890;
  assign N2892 = N2401 | N2891;
  assign N2893 = ~N2892;
  assign N2894 = N2453 | io_rocc_csr_waddr[11];
  assign N2895 = N2745 | N2894;
  assign N2896 = N2400 | N2895;
  assign N2897 = N2427 | N2896;
  assign N2898 = io_rocc_csr_waddr[6] | N2897;
  assign N2899 = io_rocc_csr_waddr[5] | N2898;
  assign N2900 = io_rocc_csr_waddr[4] | N2899;
  assign N2901 = io_rocc_csr_waddr[3] | N2900;
  assign N2902 = N2491 | N2901;
  assign N2903 = io_rocc_csr_waddr[1] | N2902;
  assign N2904 = io_rocc_csr_waddr[0] | N2903;
  assign N2905 = ~N2904;
  assign N2906 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2907 = N2745 | N2906;
  assign N2908 = N2400 | N2907;
  assign N2909 = io_rocc_csr_waddr[7] | N2908;
  assign N2910 = io_rocc_csr_waddr[6] | N2909;
  assign N2911 = io_rocc_csr_waddr[5] | N2910;
  assign N2912 = io_rocc_csr_waddr[4] | N2911;
  assign N2913 = io_rocc_csr_waddr[3] | N2912;
  assign N2914 = io_rocc_csr_waddr[2] | N2913;
  assign N2915 = io_rocc_csr_waddr[1] | N2914;
  assign N2916 = N2401 | N2915;
  assign N2917 = ~N2916;
  assign N2918 = N2453 | io_rocc_csr_waddr[11];
  assign N2919 = N2745 | N2918;
  assign N2920 = N2400 | N2919;
  assign N2921 = N2427 | N2920;
  assign N2922 = io_rocc_csr_waddr[6] | N2921;
  assign N2923 = io_rocc_csr_waddr[5] | N2922;
  assign N2924 = io_rocc_csr_waddr[4] | N2923;
  assign N2925 = io_rocc_csr_waddr[3] | N2924;
  assign N2926 = io_rocc_csr_waddr[2] | N2925;
  assign N2927 = N2454 | N2926;
  assign N2928 = io_rocc_csr_waddr[0] | N2927;
  assign N2929 = ~N2928;
  assign N2930 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2931 = N2745 | N2930;
  assign N2932 = N2400 | N2931;
  assign N2933 = io_rocc_csr_waddr[7] | N2932;
  assign N2934 = io_rocc_csr_waddr[6] | N2933;
  assign N2935 = io_rocc_csr_waddr[5] | N2934;
  assign N2936 = io_rocc_csr_waddr[4] | N2935;
  assign N2937 = io_rocc_csr_waddr[3] | N2936;
  assign N2938 = io_rocc_csr_waddr[2] | N2937;
  assign N2939 = N2454 | N2938;
  assign N2940 = io_rocc_csr_waddr[0] | N2939;
  assign N2941 = ~N2940;
  assign N2942 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N2943 = N2745 | N2942;
  assign N2944 = N2400 | N2943;
  assign N2945 = io_rocc_csr_waddr[7] | N2944;
  assign N2946 = io_rocc_csr_waddr[6] | N2945;
  assign N2947 = io_rocc_csr_waddr[5] | N2946;
  assign N2948 = io_rocc_csr_waddr[4] | N2947;
  assign N2949 = io_rocc_csr_waddr[3] | N2948;
  assign N2950 = io_rocc_csr_waddr[2] | N2949;
  assign N2951 = io_rocc_csr_waddr[1] | N2950;
  assign N2952 = io_rocc_csr_waddr[0] | N2951;
  assign N2953 = ~N2952;
  assign N2954 = N2453 | N2452;
  assign N2955 = N2745 | N2954;
  assign N2956 = N2400 | N2955;
  assign N2957 = io_rocc_csr_waddr[7] | N2956;
  assign N2958 = io_rocc_csr_waddr[6] | N2957;
  assign N2959 = io_rocc_csr_waddr[5] | N2958;
  assign N2960 = io_rocc_csr_waddr[4] | N2959;
  assign N2961 = io_rocc_csr_waddr[3] | N2960;
  assign N2962 = io_rocc_csr_waddr[2] | N2961;
  assign N2963 = io_rocc_csr_waddr[1] | N2962;
  assign N2964 = N2401 | N2963;
  assign N2965 = ~N2964;
  assign N2966 = N2453 | N2452;
  assign N2967 = N2745 | N2966;
  assign N2968 = N2400 | N2967;
  assign N2969 = io_rocc_csr_waddr[7] | N2968;
  assign N2970 = io_rocc_csr_waddr[6] | N2969;
  assign N2971 = io_rocc_csr_waddr[5] | N2970;
  assign N2972 = io_rocc_csr_waddr[4] | N2971;
  assign N2973 = io_rocc_csr_waddr[3] | N2972;
  assign N2974 = io_rocc_csr_waddr[2] | N2973;
  assign N2975 = io_rocc_csr_waddr[1] | N2974;
  assign N2976 = io_rocc_csr_waddr[0] | N2975;
  assign N2977 = ~N2976;
  assign N2978 = N2453 | io_rocc_csr_waddr[11];
  assign N2979 = N2745 | N2978;
  assign N2980 = N2400 | N2979;
  assign N2981 = io_rocc_csr_waddr[7] | N2980;
  assign N2982 = io_rocc_csr_waddr[6] | N2981;
  assign N2983 = io_rocc_csr_waddr[5] | N2982;
  assign N2984 = io_rocc_csr_waddr[4] | N2983;
  assign N2985 = io_rocc_csr_waddr[3] | N2984;
  assign N2986 = io_rocc_csr_waddr[2] | N2985;
  assign N2987 = io_rocc_csr_waddr[1] | N2986;
  assign N2988 = N2401 | N2987;
  assign N2989 = ~N2988;
  assign N2990 = io_rocc_csr_waddr[10] | N2452;
  assign N2991 = N2745 | N2990;
  assign N2992 = io_rocc_csr_waddr[8] | N2991;
  assign N2993 = io_rocc_csr_waddr[7] | N2992;
  assign N2994 = io_rocc_csr_waddr[6] | N2993;
  assign N2995 = io_rocc_csr_waddr[5] | N2994;
  assign N2996 = io_rocc_csr_waddr[4] | N2995;
  assign N2997 = io_rocc_csr_waddr[3] | N2996;
  assign N2998 = io_rocc_csr_waddr[2] | N2997;
  assign N2999 = io_rocc_csr_waddr[1] | N2998;
  assign N3000 = N2401 | N2999;
  assign N3001 = ~N3000;
  assign N3002 = N2453 | N2452;
  assign N3003 = io_rocc_csr_waddr[9] | N3002;
  assign N3004 = N2400 | N3003;
  assign N3005 = io_rocc_csr_waddr[7] | N3004;
  assign N3006 = io_rocc_csr_waddr[6] | N3005;
  assign N3007 = io_rocc_csr_waddr[5] | N3006;
  assign N3008 = io_rocc_csr_waddr[4] | N3007;
  assign N3009 = io_rocc_csr_waddr[3] | N3008;
  assign N3010 = io_rocc_csr_waddr[2] | N3009;
  assign N3011 = io_rocc_csr_waddr[1] | N3010;
  assign N3012 = N2401 | N3011;
  assign N3013 = ~N3012;
  assign N3014 = io_rocc_csr_waddr[10] | N2452;
  assign N3015 = io_rocc_csr_waddr[9] | N3014;
  assign N3016 = N2400 | N3015;
  assign N3017 = io_rocc_csr_waddr[7] | N3016;
  assign N3018 = io_rocc_csr_waddr[6] | N3017;
  assign N3019 = io_rocc_csr_waddr[5] | N3018;
  assign N3020 = io_rocc_csr_waddr[4] | N3019;
  assign N3021 = io_rocc_csr_waddr[3] | N3020;
  assign N3022 = io_rocc_csr_waddr[2] | N3021;
  assign N3023 = io_rocc_csr_waddr[1] | N3022;
  assign N3024 = N2401 | N3023;
  assign N3025 = ~N3024;
  assign N3026 = N2453 | N2452;
  assign N3027 = io_rocc_csr_waddr[9] | N3026;
  assign N3028 = io_rocc_csr_waddr[8] | N3027;
  assign N3029 = io_rocc_csr_waddr[7] | N3028;
  assign N3030 = io_rocc_csr_waddr[6] | N3029;
  assign N3031 = io_rocc_csr_waddr[5] | N3030;
  assign N3032 = io_rocc_csr_waddr[4] | N3031;
  assign N3033 = io_rocc_csr_waddr[3] | N3032;
  assign N3034 = io_rocc_csr_waddr[2] | N3033;
  assign N3035 = io_rocc_csr_waddr[1] | N3034;
  assign N3036 = N2401 | N3035;
  assign N3037 = ~N3036;
  assign N3038 = io_rocc_csr_waddr[10] | N2452;
  assign N3039 = io_rocc_csr_waddr[9] | N3038;
  assign N3040 = N2400 | N3039;
  assign N3041 = io_rocc_csr_waddr[7] | N3040;
  assign N3042 = io_rocc_csr_waddr[6] | N3041;
  assign N3043 = io_rocc_csr_waddr[5] | N3042;
  assign N3044 = io_rocc_csr_waddr[4] | N3043;
  assign N3045 = io_rocc_csr_waddr[3] | N3044;
  assign N3046 = io_rocc_csr_waddr[2] | N3045;
  assign N3047 = io_rocc_csr_waddr[1] | N3046;
  assign N3048 = io_rocc_csr_waddr[0] | N3047;
  assign N3049 = ~N3048;
  assign N3050 = N2453 | N2452;
  assign N3051 = io_rocc_csr_waddr[9] | N3050;
  assign N3052 = io_rocc_csr_waddr[8] | N3051;
  assign N3053 = io_rocc_csr_waddr[7] | N3052;
  assign N3054 = io_rocc_csr_waddr[6] | N3053;
  assign N3055 = io_rocc_csr_waddr[5] | N3054;
  assign N3056 = io_rocc_csr_waddr[4] | N3055;
  assign N3057 = io_rocc_csr_waddr[3] | N3056;
  assign N3058 = io_rocc_csr_waddr[2] | N3057;
  assign N3059 = io_rocc_csr_waddr[1] | N3058;
  assign N3060 = io_rocc_csr_waddr[0] | N3059;
  assign N3061 = ~N3060;
  assign N3062 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N3063 = io_rocc_csr_waddr[9] | N3062;
  assign N3064 = io_rocc_csr_waddr[8] | N3063;
  assign N3065 = io_rocc_csr_waddr[7] | N3064;
  assign N3066 = io_rocc_csr_waddr[6] | N3065;
  assign N3067 = io_rocc_csr_waddr[5] | N3066;
  assign N3068 = io_rocc_csr_waddr[4] | N3067;
  assign N3069 = io_rocc_csr_waddr[3] | N3068;
  assign N3070 = io_rocc_csr_waddr[2] | N3069;
  assign N3071 = N2454 | N3070;
  assign N3072 = N2401 | N3071;
  assign N3073 = ~N3072;
  assign N3074 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N3075 = io_rocc_csr_waddr[9] | N3074;
  assign N3076 = io_rocc_csr_waddr[8] | N3075;
  assign N3077 = io_rocc_csr_waddr[7] | N3076;
  assign N3078 = io_rocc_csr_waddr[6] | N3077;
  assign N3079 = io_rocc_csr_waddr[5] | N3078;
  assign N3080 = io_rocc_csr_waddr[4] | N3079;
  assign N3081 = io_rocc_csr_waddr[3] | N3080;
  assign N3082 = io_rocc_csr_waddr[2] | N3081;
  assign N3083 = io_rocc_csr_waddr[1] | N3082;
  assign N3084 = N2401 | N3083;
  assign N3085 = ~N3084;
  assign N3086 = io_rocc_csr_waddr[10] | io_rocc_csr_waddr[11];
  assign N3087 = io_rocc_csr_waddr[9] | N3086;
  assign N3088 = io_rocc_csr_waddr[8] | N3087;
  assign N3089 = io_rocc_csr_waddr[7] | N3088;
  assign N3090 = io_rocc_csr_waddr[6] | N3089;
  assign N3091 = io_rocc_csr_waddr[5] | N3090;
  assign N3092 = io_rocc_csr_waddr[4] | N3091;
  assign N3093 = io_rocc_csr_waddr[3] | N3092;
  assign N3094 = io_rocc_csr_waddr[2] | N3093;
  assign N3095 = N2454 | N3094;
  assign N3096 = io_rocc_csr_waddr[0] | N3095;
  assign N3097 = ~N3096;
  assign N3098 = io_rw_cmd[0] | N2387;
  assign N3099 = io_rw_cmd[0] | N2398;
  assign N3100 = ~N3099;
  assign T947 = io_status_prv + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign { T326[6:6], T325 } = io_time[5:0] + 1'b1;
  assign T329 = io_time[63:6] + 1'b1;
  assign { T444_63, T444[40:40] } = 1'b0 - T444[39];
  assign { T839_63, T839[40:40] } = 1'b0 - T839[39];
  assign { T439[63:63], T439_39 } = 1'b0 - T357[38];
  assign T364 = { io_status_prv, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } + reg_mtvec[39:0];
  assign { T452_63, T452[40:40] } = 1'b0 - T452[39];
  assign { T834_63, T834[40:40] } = 1'b0 - T834[39];
  assign { T586[6:6], T585 } = T582[5:0] + 1'b1;
  assign T590 = T582[63:6] + 1'b1;
  assign { T599[6:6], T598 } = T595[5:0] + 1'b1;
  assign T603 = T595[63:6] + 1'b1;
  assign { T612[6:6], T611 } = T608[5:0] + 1'b1;
  assign T616 = T608[63:6] + 1'b1;
  assign { T625[6:6], T624 } = T621[5:0] + 1'b1;
  assign T629 = T621[63:6] + 1'b1;
  assign { T638[6:6], T637 } = T634[5:0] + 1'b1;
  assign T642 = T634[63:6] + 1'b1;
  assign { T651[6:6], T650 } = T647[5:0] + 1'b1;
  assign T655 = T647[63:6] + 1'b1;
  assign { T664[6:6], T663 } = T660[5:0] + 1'b1;
  assign T668 = T660[63:6] + 1'b1;
  assign { T677[6:6], T676 } = T673[5:0] + 1'b1;
  assign T681 = T673[63:6] + 1'b1;
  assign { T690[6:6], T689 } = T686[5:0] + 1'b1;
  assign T694 = T686[63:6] + 1'b1;
  assign { T703[6:6], T702 } = T699[5:0] + 1'b1;
  assign T707 = T699[63:6] + 1'b1;
  assign { T716[6:6], T715 } = T712[5:0] + 1'b1;
  assign T720 = T712[63:6] + 1'b1;
  assign { T729[6:6], T728 } = T725[5:0] + 1'b1;
  assign T733 = T725[63:6] + 1'b1;
  assign { T742[6:6], T741 } = T738[5:0] + 1'b1;
  assign T746 = T738[63:6] + 1'b1;
  assign { T755[6:6], T754 } = T751[5:0] + 1'b1;
  assign T759 = T751[63:6] + 1'b1;
  assign { T768[6:6], T767 } = T764[5:0] + 1'b1;
  assign T772 = T764[63:6] + 1'b1;
  assign { T781[6:6], T780 } = T777[5:0] + 1'b1;
  assign T785 = T777[63:6] + 1'b1;
  assign { T795[6:6], T794 } = T790[5:0] + 1'b1;
  assign T802 = T790[63:6] + 1'b1;
  assign io_status_fs = 1'b0 - N2795;
  assign io_status_xs = 1'b0 - N2796;
  assign io_rocc_csr_wdata = (N0)? io_rw_wdata : 
                             (N1)? T36 : 1'b0;
  assign N0 = N2389;
  assign N1 = N2388;
  assign T36 = (N2)? T48 : 
               (N3)? T37 : 1'b0;
  assign N2 = N2393;
  assign N3 = N2392;
  assign T37 = (N4)? T46 : 
               (N5)? io_host_csr_resp_bits : 1'b0;
  assign N4 = N2396;
  assign N5 = N2395;
  assign io_rocc_csr_waddr = (N6)? io_rw_addr : 
                             (N7)? host_csr_bits_addr : 1'b0;
  assign N6 = cpu_ren;
  assign N7 = N163;
  assign { io_interrupt_cause[63:63], io_interrupt_cause[1:0] } = (N8)? { 1'b1, 1'b1, 1'b1 } : 
                                                                  (N9)? { T218_63, T218 } : 1'b0;
  assign N8 = T312;
  assign N9 = N164;
  assign { T218_63, T218[0:0] } = (N10)? { 1'b1, 1'b0 } : 
                                  (N11)? { T219[63:63], T219_0 } : 1'b0;
  assign N10 = T218[1];
  assign N11 = N165;
  assign { T219[63:63], T219_0 } = (N12)? { 1'b1, 1'b1 } : 
                                   (N13)? { T220[63:63], T220_0 } : 1'b0;
  assign N12 = T285;
  assign N13 = N166;
  assign T220[63] = (N14)? 1'b1 : 
                    (N15)? T221[63] : 1'b0;
  assign N14 = T220_0;
  assign N15 = N167;
  assign T221[63] = (N16)? 1'b1 : 
                    (N17)? T222[63] : 1'b0;
  assign N16 = T260;
  assign N17 = N168;
  assign T924 = (N18)? io_rocc_csr_wdata[7:5] : 
                (N19)? T319 : 1'b0;
  assign N18 = T322;
  assign N19 = N169;
  assign T319 = (N20)? io_rocc_csr_wdata[2:0] : 
                (N21)? io_fcsr_rm : 1'b0;
  assign N20 = T320;
  assign N21 = N170;
  assign io_evec = (N22)? T364 : 
                   (N23)? T931 : 1'b0;
  assign N22 = T369;
  assign N23 = N171;
  assign T931 = (N24)? { T357[38:38], T357 } : 
                (N25)? T340 : 1'b0;
  assign N24 = maybe_insn_redirect_trap;
  assign N25 = N172;
  assign T340 = (N26)? T839[39:0] : 
                (N27)? T444[39:0] : 1'b0;
  assign N26 = io_status_prv[1];
  assign N27 = N173;
  assign T932 = (N28)? T343 : 
                (N29)? T933 : 1'b0;
  assign N28 = T346;
  assign N29 = N174;
  assign T933 = (N30)? T839[39:0] : 
                (N31)? T444[39:0] : 1'b0;
  assign N30 = T216[0];
  assign N31 = N175;
  assign T934 = (N32)? T352 : 
                (N33)? T935 : 1'b0;
  assign N32 = T355;
  assign N33 = N176;
  assign T935 = (N34)? T349 : 
                (N35)? T839[39:0] : 1'b0;
  assign N34 = T25;
  assign N35 = N177;
  assign T936 = (N36)? T359 : 
                (N37)? T357 : 1'b0;
  assign N36 = T362;
  assign N37 = N178;
  assign some_interrupt_pending = (N38)? 1'b1 : 
                                  (N39)? T421 : 1'b0;
  assign N38 = T435;
  assign N39 = N179;
  assign T421 = (N40)? 1'b1 : 
                (N41)? T422 : 1'b0;
  assign N40 = T433;
  assign N41 = N180;
  assign T422 = (N42)? 1'b1 : 
                (N43)? T423 : 1'b0;
  assign N42 = T431;
  assign N43 = N181;
  assign T423 = (N44)? 1'b1 : 
                (N45)? T424 : 1'b0;
  assign N44 = T429;
  assign N45 = N182;
  assign T424 = (N46)? 1'b1 : 
                (N47)? T425 : 1'b0;
  assign N46 = T427;
  assign N47 = N183;
  assign T438 = (N48)? { T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439[63:63], T439_39, T357 } : 
                (N49)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = N2413;
  assign N49 = N2412;
  assign T443 = (N50)? { T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444_63, T444 } : 
                (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N50 = N2426;
  assign N51 = N2425;
  assign T945 = (N52)? io_ptbr : 
                (N53)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = N2451;
  assign N53 = N2450;
  assign T451 = (N54)? { T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452_63, T452 } : 
                (N55)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N54 = N2466;
  assign N55 = N2465;
  assign T457[39] = (N56)? N2057 : 
                    (N57)? N2081 : 1'b0;
  assign N56 = T463;
  assign N57 = N184;
  assign T478 = (N58)? reg_scause : 
                (N59)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N58 = N2478;
  assign N59 = N2477;
  assign T492 = (N60)? reg_sscratch : 
                (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = N2490;
  assign N61 = N2489;
  assign { T949[5:5], T949_1 } = (N62)? { T497[5:5], T497_1 } : 
                                 (N63)? { 1'b0, 1'b0 } : 1'b0;
  assign N62 = N2503;
  assign N63 = N2502;
  assign { T950[5:5], T950_1 } = (N64)? { T515[5:5], T515_1 } : 
                                 (N65)? { 1'b0, 1'b0 } : 1'b0;
  assign N64 = N2515;
  assign N65 = N2514;
  assign { T532_63, T532_31, T532, T532_4, T532_3, T532_0 } = (N66)? { io_status_sd, io_status_sd_rv32, io_status_mprv, io_status_xs, io_status_fs, io_status_prv1[0:0], io_status_ie1, io_status_ie } : 
                                                              (N67)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N66 = N2527;
  assign N67 = N2526;
  assign T581 = (N68)? T582 : 
                (N69)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N68 = N2540;
  assign N69 = N2539;
  assign T594 = (N70)? T595 : 
                (N71)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N70 = N2552;
  assign N71 = N2551;
  assign T607 = (N72)? T608 : 
                (N73)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N72 = N2564;
  assign N73 = N2563;
  assign T620 = (N74)? T621 : 
                (N75)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N74 = N2576;
  assign N75 = N2575;
  assign T633 = (N76)? T634 : 
                (N77)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N76 = N2588;
  assign N77 = N2587;
  assign T646 = (N78)? T647 : 
                (N79)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N78 = N2600;
  assign N79 = N2599;
  assign T659 = (N80)? T660 : 
                (N81)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N80 = N2612;
  assign N81 = N2611;
  assign T672 = (N82)? T673 : 
                (N83)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N82 = N2624;
  assign N83 = N2623;
  assign T685 = (N84)? T686 : 
                (N85)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N84 = N2636;
  assign N85 = N2635;
  assign T698 = (N86)? T699 : 
                (N87)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N86 = N2648;
  assign N87 = N2647;
  assign T711 = (N88)? T712 : 
                (N89)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N88 = N2660;
  assign N89 = N2659;
  assign T724 = (N90)? T725 : 
                (N91)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N90 = N2672;
  assign N91 = N2671;
  assign T737 = (N92)? T738 : 
                (N93)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N92 = N2684;
  assign N93 = N2683;
  assign T750 = (N94)? T751 : 
                (N95)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N94 = N2696;
  assign N95 = N2695;
  assign T763 = (N96)? T764 : 
                (N97)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N96 = N2708;
  assign N97 = N2707;
  assign T776 = (N98)? T777 : 
                (N99)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N98 = N2720;
  assign N99 = N2719;
  assign T789 = (N100)? T790 : 
                (N101)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N100 = N2732;
  assign N101 = N2731;
  assign T807 = (N102)? T790 : 
                (N103)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N102 = N2744;
  assign N103 = N2743;
  assign T809 = (N104)? reg_fromhost : 
                (N105)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N104 = N2757;
  assign N105 = N2756;
  assign T811 = (N106)? reg_tohost : 
                (N107)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N106 = N2769;
  assign N107 = N2768;
  assign T1003[0] = (N108)? io_host_debug_stats_csr : 
                    (N109)? 1'b0 : 1'b0;
  assign N108 = N2781;
  assign N109 = N2780;
  assign T1005[0] = (N110)? io_host_id : 
                    (N111)? 1'b0 : 1'b0;
  assign N110 = N2794;
  assign N111 = N2793;
  assign T829 = (N112)? reg_mtimecmp : 
                (N113)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N112 = N2809;
  assign N113 = N2808;
  assign T831 = (N114)? reg_mcause : 
                (N115)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N114 = N2821;
  assign N115 = N2820;
  assign T833 = (N116)? { T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834_63, T834 } : 
                (N117)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N116 = N2833;
  assign N117 = N2832;
  assign T838 = (N118)? { T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839_63, T839 } : 
                (N119)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N118 = N2845;
  assign N119 = N2844;
  assign T843 = (N120)? reg_mscratch : 
                (N121)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N120 = N2857;
  assign N121 = N2856;
  assign T1008 = (N122)? { T848_7, T848_6, T497[5:5], T848, T497_1, T848_0 } : 
                 (N123)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N122 = N2869;
  assign N123 = N2868;
  assign T1013 = (N124)? { T858_7, T858_6, T515[5:5], T858, T515_1, T858_0 } : 
                 (N125)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N124 = N2881;
  assign N125 = N2880;
  assign T870 = (N126)? reg_mtvec : 
                (N127)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N126 = N2917;
  assign N127 = N2916;
  assign T874 = (N128)? { io_status_sd, io_status_zero2, io_status_sd_rv32, io_status_zero1, io_status_vm, io_status_mprv, io_status_xs, io_status_fs, io_status_prv3, io_status_ie3, io_status_prv2, io_status_ie2, io_status_prv1, io_status_ie1, io_status_prv, io_status_ie } : 
                (N129)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N128 = N2953;
  assign N129 = N2952;
  assign T879 = (N130)? read_time : 
                (N131)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N130 = N2989;
  assign N131 = N2988;
  assign T881 = (N132)? read_time : 
                (N133)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N132 = N3001;
  assign N133 = N3000;
  assign T883 = (N134)? read_time : 
                (N135)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N134 = N3013;
  assign N135 = N3012;
  assign T885 = (N136)? read_time : 
                (N137)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N136 = N3025;
  assign N137 = N3024;
  assign T887 = (N138)? read_time : 
                (N139)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N138 = N3037;
  assign N139 = N3036;
  assign T889 = (N140)? io_time : 
                (N141)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N140 = N3049;
  assign N141 = N3048;
  assign T891 = (N142)? io_time : 
                (N143)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N142 = N3061;
  assign N143 = N3060;
  assign T893 = (N144)? { io_fcsr_rm, T894 } : 
                (N145)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N144 = N3073;
  assign N145 = N3072;
  assign T1021 = (N18)? io_rocc_csr_wdata[4:0] : 
                 (N19)? T896 : 1'b0;
  assign T896 = (N146)? io_rocc_csr_wdata[4:0] : 
                (N147)? T1022 : 1'b0;
  assign N146 = T899;
  assign N147 = N185;
  assign T1022 = (N148)? T898 : 
                 (N149)? T894 : 1'b0;
  assign N148 = io_fcsr_flags_valid;
  assign N149 = N186;
  assign T1024 = (N150)? io_fcsr_rm : 
                 (N151)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N150 = N3097;
  assign N151 = N3096;
  assign T902 = (N152)? T894 : 
                (N153)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N152 = N3085;
  assign N153 = N3084;
  assign N192 = (N154)? 1'b1 : 
                (N1882)? 1'b1 : 
                (N1885)? 1'b1 : 
                (N1888)? 1'b1 : 
                (N1891)? 1'b1 : 
                (N191)? 1'b0 : 1'b0;
  assign N154 = reset;
  assign { N194, N193 } = (N154)? { 1'b1, 1'b1 } : 
                          (N1882)? io_rocc_csr_wdata[2:1] : 
                          (N1885)? { 1'b0, 1'b1 } : 
                          (N1888)? io_status_prv1 : 
                          (N1891)? { 1'b1, 1'b1 } : 1'b0;
  assign N200 = (N154)? 1'b1 : 
                (N1892)? 1'b1 : 
                (N1895)? 1'b1 : 
                (N1898)? 1'b1 : 
                (N1900)? 1'b1 : 
                (N199)? 1'b0 : 1'b0;
  assign { N202, N201 } = (N154)? { 1'b1, 1'b1 } : 
                          (N1892)? { 1'b0, io_rocc_csr_wdata[4:4] } : 
                          (N1895)? io_rocc_csr_wdata[5:4] : 
                          (N1898)? io_status_prv2 : 
                          (N1900)? io_status_prv : 1'b0;
  assign N207 = (N154)? 1'b1 : 
                (N1902)? 1'b1 : 
                (N1905)? 1'b1 : 
                (N1907)? 1'b1 : 
                (N206)? 1'b0 : 1'b0;
  assign { N209, N208 } = (N154)? { 1'b0, 1'b0 } : 
                          (N1902)? io_rocc_csr_wdata[8:7] : 
                          (N1905)? { 1'b0, 1'b0 } : 
                          (N1907)? io_status_prv1 : 1'b0;
  assign N212 = (N155)? 1'b1 : 
                (N1909)? 1'b1 : 
                (N211)? 1'b0 : 1'b0;
  assign N155 = host_csr_req_fire;
  assign { N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213 } = (N155)? io_rw_rdata : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1909)? io_host_csr_req_bits_data : 1'b0;
  assign N278 = (N156)? cpu_ren : 
                (N157)? T45 : 1'b0;
  assign N156 = host_csr_req_valid;
  assign N157 = N277;
  assign N284 = (N154)? 1'b1 : 
                (N1910)? 1'b1 : 
                (N1912)? 1'b1 : 
                (N1915)? 1'b1 : 
                (N1917)? 1'b1 : 
                (N283)? 1'b0 : 1'b0;
  assign N285 = (N154)? 1'b0 : 
                (N1910)? io_rocc_csr_wdata[0] : 
                (N1912)? io_rocc_csr_wdata[0] : 
                (N1915)? io_status_ie1 : 
                (N1917)? 1'b0 : 1'b0;
  assign N291 = (N154)? 1'b1 : 
                (N1918)? 1'b1 : 
                (N1920)? 1'b1 : 
                (N1922)? 1'b1 : 
                (N1924)? 1'b1 : 
                (N290)? 1'b0 : 1'b0;
  assign N292 = (N154)? 1'b0 : 
                (N1918)? io_rocc_csr_wdata[3] : 
                (N1920)? io_rocc_csr_wdata[3] : 
                (N1922)? io_status_ie2 : 
                (N1924)? io_status_ie : 1'b0;
  assign N297 = (N154)? 1'b1 : 
                (N1925)? 1'b1 : 
                (N1927)? 1'b1 : 
                (N1929)? 1'b1 : 
                (N296)? 1'b0 : 1'b0;
  assign N298 = (N154)? 1'b0 : 
                (N1925)? io_rocc_csr_wdata[6] : 
                (N1927)? 1'b1 : 
                (N1929)? io_status_ie1 : 1'b0;
  assign N302 = (N154)? 1'b1 : 
                (N1930)? 1'b1 : 
                (N1933)? 1'b1 : 
                (N301)? 1'b0 : 1'b0;
  assign N303 = (N154)? 1'b0 : 
                (N1930)? io_rocc_csr_wdata[1] : 
                (N1933)? io_rocc_csr_wdata[1] : 1'b0;
  assign N307 = (N154)? 1'b1 : 
                (N1934)? 1'b1 : 
                (N1937)? 1'b1 : 
                (N306)? 1'b0 : 1'b0;
  assign N308 = (N154)? 1'b0 : 
                (N1934)? io_rocc_csr_wdata[1] : 
                (N1937)? io_rocc_csr_wdata[1] : 1'b0;
  assign N312 = (N154)? 1'b1 : 
                (N1938)? 1'b1 : 
                (N1941)? 1'b1 : 
                (N311)? 1'b0 : 1'b0;
  assign N313 = (N154)? 1'b0 : 
                (N1938)? io_rocc_csr_wdata[0] : 
                (N1941)? io_rocc_csr_wdata[3] : 1'b0;
  assign N316 = (N154)? 1'b1 : 
                (N1942)? 1'b1 : 
                (N315)? 1'b0 : 1'b0;
  assign N317 = (N154)? 1'b0 : 
                (N1942)? io_rocc_csr_wdata[3] : 1'b0;
  assign N320 = (N154)? 1'b1 : 
                (N1943)? 1'b1 : 
                (N319)? 1'b0 : 1'b0;
  assign N321 = (N154)? 1'b0 : 
                (N1943)? io_rocc_csr_wdata[5] : 1'b0;
  assign N325 = (N154)? 1'b1 : 
                (N1944)? 1'b1 : 
                (N1946)? 1'b1 : 
                (N324)? 1'b0 : 1'b0;
  assign N326 = (N154)? 1'b0 : 
                (N1944)? io_rocc_csr_wdata[5] : 
                (N1946)? io_rocc_csr_wdata[5] : 1'b0;
  assign N330 = (N154)? 1'b1 : 
                (N1947)? 1'b1 : 
                (N1950)? 1'b1 : 
                (N329)? 1'b0 : 1'b0;
  assign N331 = (N154)? 1'b0 : 
                (N1947)? 1'b0 : 
                (N1950)? 1'b1 : 1'b0;
  assign N334 = (N154)? 1'b1 : 
                (N1951)? 1'b1 : 
                (N333)? 1'b0 : 1'b0;
  assign N335 = (N154)? 1'b0 : 
                (N1951)? io_rocc_csr_wdata[7] : 1'b0;
  assign N338 = (N154)? 1'b1 : 
                (N1952)? 1'b1 : 
                (N337)? 1'b0 : 1'b0;
  assign { N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1952)? io_rocc_csr_wdata : 1'b0;
  assign { N409, N408, N407, N406, N405, N404 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N158)? T325 : 1'b0;
  assign N158 = N403;
  assign N412 = (N154)? 1'b1 : 
                (N1953)? 1'b1 : 
                (N411)? 1'b0 : 1'b0;
  assign { N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                          (N1953)? T329 : 1'b0;
  assign N473 = (N154)? 1'b1 : 
                (N1954)? 1'b1 : 
                (N472)? 1'b0 : 1'b0;
  assign N477 = (N154)? 1'b1 : 
                (N1955)? 1'b1 : 
                (N1957)? 1'b1 : 
                (N476)? 1'b0 : 1'b0;
  assign { N479, N478 } = (N154)? { 1'b0, 1'b0 } : 
                          (N1955)? io_rocc_csr_wdata[13:12] : 
                          (N1957)? io_rocc_csr_wdata[13:12] : 1'b0;
  assign N483 = (N154)? 1'b1 : 
                (N1958)? 1'b1 : 
                (N1960)? 1'b1 : 
                (N482)? 1'b0 : 1'b0;
  assign { N485, N484 } = (N154)? { 1'b0, 1'b0 } : 
                          (N1958)? io_rocc_csr_wdata[15:14] : 
                          (N1960)? io_rocc_csr_wdata[15:14] : 1'b0;
  assign N490 = (N154)? 1'b1 : 
                (N1961)? 1'b1 : 
                (N1963)? 1'b1 : 
                (N1965)? 1'b1 : 
                (N489)? 1'b0 : 1'b0;
  assign N491 = (N154)? 1'b0 : 
                (N1961)? io_rocc_csr_wdata[16] : 
                (N1963)? io_rocc_csr_wdata[16] : 
                (N1965)? 1'b0 : 1'b0;
  assign N495 = (N154)? 1'b1 : 
                (N1966)? 1'b1 : 
                (N1969)? 1'b1 : 
                (N494)? 1'b0 : 1'b0;
  assign N496 = (N154)? 1'b0 : 
                (N1966)? 1'b1 : 
                (N1969)? 1'b0 : 1'b0;
  assign N500 = (N154)? 1'b1 : 
                (N1970)? 1'b1 : 
                (N1973)? 1'b1 : 
                (N499)? 1'b0 : 1'b0;
  assign N501 = (N154)? 1'b0 : 
                (N1970)? 1'b0 : 
                (N1973)? 1'b1 : 1'b0;
  assign N505 = (N159)? 1'b1 : 
                (N1975)? 1'b1 : 
                (N1978)? 1'b1 : 
                (N504)? 1'b0 : 1'b0;
  assign N159 = T474;
  assign { N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506 } = (N159)? io_rocc_csr_wdata[39:0] : 
                                                                                                                                                                                                                                                              (N1975)? { T457[39:39], io_rw_wdata[38:0] } : 
                                                                                                                                                                                                                                                              (N1978)? io_pc : 1'b0;
  assign N551 = (N160)? 1'b1 : 
                (N1980)? 1'b1 : 
                (N1983)? 1'b1 : 
                (N1986)? 1'b1 : 
                (N1989)? 1'b1 : 
                (N550)? 1'b0 : 1'b0;
  assign N160 = T490;
  assign { N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552 } = (N160)? { io_rocc_csr_wdata[63:63], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, io_rocc_csr_wdata[4:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1980)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T947 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1983)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1986)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N1989)? io_cause : 1'b0;
  assign N618 = (N154)? 1'b1 : 
                (N1990)? 1'b1 : 
                (N617)? 1'b0 : 1'b0;
  assign { N624, N623, N622, N621, N620, N619 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N1990)? T585 : 1'b0;
  assign N627 = (N154)? 1'b1 : 
                (N1991)? 1'b1 : 
                (N626)? 1'b0 : 1'b0;
  assign { N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                          (N1991)? T590 : 1'b0;
  assign N688 = (N154)? 1'b1 : 
                (N1992)? 1'b1 : 
                (N687)? 1'b0 : 1'b0;
  assign { N694, N693, N692, N691, N690, N689 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N1992)? T598 : 1'b0;
  assign N697 = (N154)? 1'b1 : 
                (N1993)? 1'b1 : 
                (N696)? 1'b0 : 1'b0;
  assign { N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                          (N1993)? T603 : 1'b0;
  assign N758 = (N154)? 1'b1 : 
                (N1994)? 1'b1 : 
                (N757)? 1'b0 : 1'b0;
  assign { N764, N763, N762, N761, N760, N759 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N1994)? T611 : 1'b0;
  assign N767 = (N154)? 1'b1 : 
                (N1995)? 1'b1 : 
                (N766)? 1'b0 : 1'b0;
  assign { N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                          (N1995)? T616 : 1'b0;
  assign N828 = (N154)? 1'b1 : 
                (N1996)? 1'b1 : 
                (N827)? 1'b0 : 1'b0;
  assign { N834, N833, N832, N831, N830, N829 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N1996)? T624 : 1'b0;
  assign N837 = (N154)? 1'b1 : 
                (N1997)? 1'b1 : 
                (N836)? 1'b0 : 1'b0;
  assign { N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                          (N1997)? T629 : 1'b0;
  assign N898 = (N154)? 1'b1 : 
                (N1998)? 1'b1 : 
                (N897)? 1'b0 : 1'b0;
  assign { N904, N903, N902, N901, N900, N899 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N1998)? T637 : 1'b0;
  assign N907 = (N154)? 1'b1 : 
                (N1999)? 1'b1 : 
                (N906)? 1'b0 : 1'b0;
  assign { N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                          (N1999)? T642 : 1'b0;
  assign N968 = (N154)? 1'b1 : 
                (N2000)? 1'b1 : 
                (N967)? 1'b0 : 1'b0;
  assign { N974, N973, N972, N971, N970, N969 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N2000)? T650 : 1'b0;
  assign N977 = (N154)? 1'b1 : 
                (N2001)? 1'b1 : 
                (N976)? 1'b0 : 1'b0;
  assign { N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N2001)? T655 : 1'b0;
  assign N1038 = (N154)? 1'b1 : 
                 (N2002)? 1'b1 : 
                 (N1037)? 1'b0 : 1'b0;
  assign { N1044, N1043, N1042, N1041, N1040, N1039 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2002)? T663 : 1'b0;
  assign N1047 = (N154)? 1'b1 : 
                 (N2003)? 1'b1 : 
                 (N1046)? 1'b0 : 1'b0;
  assign { N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2003)? T668 : 1'b0;
  assign N1108 = (N154)? 1'b1 : 
                 (N2004)? 1'b1 : 
                 (N1107)? 1'b0 : 1'b0;
  assign { N1114, N1113, N1112, N1111, N1110, N1109 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2004)? T676 : 1'b0;
  assign N1117 = (N154)? 1'b1 : 
                 (N2005)? 1'b1 : 
                 (N1116)? 1'b0 : 1'b0;
  assign { N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2005)? T681 : 1'b0;
  assign N1178 = (N154)? 1'b1 : 
                 (N2006)? 1'b1 : 
                 (N1177)? 1'b0 : 1'b0;
  assign { N1184, N1183, N1182, N1181, N1180, N1179 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2006)? T689 : 1'b0;
  assign N1187 = (N154)? 1'b1 : 
                 (N2007)? 1'b1 : 
                 (N1186)? 1'b0 : 1'b0;
  assign { N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2007)? T694 : 1'b0;
  assign N1248 = (N154)? 1'b1 : 
                 (N2008)? 1'b1 : 
                 (N1247)? 1'b0 : 1'b0;
  assign { N1254, N1253, N1252, N1251, N1250, N1249 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2008)? T702 : 1'b0;
  assign N1257 = (N154)? 1'b1 : 
                 (N2009)? 1'b1 : 
                 (N1256)? 1'b0 : 1'b0;
  assign { N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2009)? T707 : 1'b0;
  assign N1318 = (N154)? 1'b1 : 
                 (N2010)? 1'b1 : 
                 (N1317)? 1'b0 : 1'b0;
  assign { N1324, N1323, N1322, N1321, N1320, N1319 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2010)? T715 : 1'b0;
  assign N1327 = (N154)? 1'b1 : 
                 (N2011)? 1'b1 : 
                 (N1326)? 1'b0 : 1'b0;
  assign { N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2011)? T720 : 1'b0;
  assign N1388 = (N154)? 1'b1 : 
                 (N2012)? 1'b1 : 
                 (N1387)? 1'b0 : 1'b0;
  assign { N1394, N1393, N1392, N1391, N1390, N1389 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2012)? T728 : 1'b0;
  assign N1397 = (N154)? 1'b1 : 
                 (N2013)? 1'b1 : 
                 (N1396)? 1'b0 : 1'b0;
  assign { N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2013)? T733 : 1'b0;
  assign N1458 = (N154)? 1'b1 : 
                 (N2014)? 1'b1 : 
                 (N1457)? 1'b0 : 1'b0;
  assign { N1464, N1463, N1462, N1461, N1460, N1459 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2014)? T741 : 1'b0;
  assign N1467 = (N154)? 1'b1 : 
                 (N2015)? 1'b1 : 
                 (N1466)? 1'b0 : 1'b0;
  assign { N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2015)? T746 : 1'b0;
  assign N1528 = (N154)? 1'b1 : 
                 (N2016)? 1'b1 : 
                 (N1527)? 1'b0 : 1'b0;
  assign { N1534, N1533, N1532, N1531, N1530, N1529 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2016)? T754 : 1'b0;
  assign N1537 = (N154)? 1'b1 : 
                 (N2017)? 1'b1 : 
                 (N1536)? 1'b0 : 1'b0;
  assign { N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2017)? T759 : 1'b0;
  assign N1598 = (N154)? 1'b1 : 
                 (N2018)? 1'b1 : 
                 (N1597)? 1'b0 : 1'b0;
  assign { N1604, N1603, N1602, N1601, N1600, N1599 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2018)? T767 : 1'b0;
  assign N1607 = (N154)? 1'b1 : 
                 (N2019)? 1'b1 : 
                 (N1606)? 1'b0 : 1'b0;
  assign { N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2019)? T772 : 1'b0;
  assign N1668 = (N154)? 1'b1 : 
                 (N2020)? 1'b1 : 
                 (N1667)? 1'b0 : 1'b0;
  assign { N1674, N1673, N1672, N1671, N1670, N1669 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2020)? T780 : 1'b0;
  assign N1677 = (N154)? 1'b1 : 
                 (N2021)? 1'b1 : 
                 (N1676)? 1'b0 : 1'b0;
  assign { N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2021)? T785 : 1'b0;
  assign N1739 = (N154)? 1'b1 : 
                 (N2022)? 1'b1 : 
                 (N2025)? 1'b1 : 
                 (N1738)? 1'b0 : 1'b0;
  assign { N1745, N1744, N1743, N1742, N1741, N1740 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2022)? io_rocc_csr_wdata[5:0] : 
                                                        (N2025)? T794 : 1'b0;
  assign N1749 = (N154)? 1'b1 : 
                 (N2026)? 1'b1 : 
                 (N2028)? 1'b1 : 
                 (N1748)? 1'b0 : 1'b0;
  assign { N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2026)? io_rocc_csr_wdata[63:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N2028)? T802 : 1'b0;
  assign N1811 = (N154)? 1'b1 : 
                 (N2029)? 1'b1 : 
                 (N2032)? 1'b1 : 
                 (N1810)? 1'b0 : 1'b0;
  assign { N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812 } = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2029)? io_rocc_csr_wdata : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2032)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1878 = (N154)? 1'b1 : 
                 (N2033)? 1'b1 : 
                 (N1877)? 1'b0 : 1'b0;
  assign N1879 = (N154)? 1'b0 : 
                 (N2033)? io_rocc_csr_wdata[0] : 1'b0;
  assign N1881 = (N161)? T905 : 
                 (N162)? host_csr_req_fire : 1'b0;
  assign N161 = io_host_csr_resp_valid;
  assign N162 = N1880;
  assign io_csr_xcpt = T11 | insn_break;
  assign insn_break = T7 & N3100;
  assign T7 = T9 & io_rw_addr[0];
  assign T9 = ~io_rw_addr[8];
  assign T11 = T17 | insn_call;
  assign insn_call = T12 & N3100;
  assign T12 = T15 & T13;
  assign T13 = ~io_rw_addr[0];
  assign T15 = ~io_rw_addr[8];
  assign T17 = T94 | T18;
  assign T18 = N3100 & T19;
  assign T19 = ~priv_sufficient;
  assign T25 = io_exception | io_csr_xcpt;
  assign T40 = io_host_csr_req_ready & io_host_csr_req_valid;
  assign host_csr_req_fire = host_csr_req_valid & T41;
  assign T41 = ~cpu_ren;
  assign cpu_ren = N3098 & T42;
  assign T42 = ~N3100;
  assign T45 = io_host_csr_req_ready & io_host_csr_req_valid;
  assign T46[63] = io_rw_rdata[63] | io_rw_wdata[63];
  assign T46[62] = io_rw_rdata[62] | io_rw_wdata[62];
  assign T46[61] = io_rw_rdata[61] | io_rw_wdata[61];
  assign T46[60] = io_rw_rdata[60] | io_rw_wdata[60];
  assign T46[59] = io_rw_rdata[59] | io_rw_wdata[59];
  assign T46[58] = io_rw_rdata[58] | io_rw_wdata[58];
  assign T46[57] = io_rw_rdata[57] | io_rw_wdata[57];
  assign T46[56] = io_rw_rdata[56] | io_rw_wdata[56];
  assign T46[55] = io_rw_rdata[55] | io_rw_wdata[55];
  assign T46[54] = io_rw_rdata[54] | io_rw_wdata[54];
  assign T46[53] = io_rw_rdata[53] | io_rw_wdata[53];
  assign T46[52] = io_rw_rdata[52] | io_rw_wdata[52];
  assign T46[51] = io_rw_rdata[51] | io_rw_wdata[51];
  assign T46[50] = io_rw_rdata[50] | io_rw_wdata[50];
  assign T46[49] = io_rw_rdata[49] | io_rw_wdata[49];
  assign T46[48] = io_rw_rdata[48] | io_rw_wdata[48];
  assign T46[47] = io_rw_rdata[47] | io_rw_wdata[47];
  assign T46[46] = io_rw_rdata[46] | io_rw_wdata[46];
  assign T46[45] = io_rw_rdata[45] | io_rw_wdata[45];
  assign T46[44] = io_rw_rdata[44] | io_rw_wdata[44];
  assign T46[43] = io_rw_rdata[43] | io_rw_wdata[43];
  assign T46[42] = io_rw_rdata[42] | io_rw_wdata[42];
  assign T46[41] = io_rw_rdata[41] | io_rw_wdata[41];
  assign T46[40] = io_rw_rdata[40] | io_rw_wdata[40];
  assign T46[39] = io_rw_rdata[39] | io_rw_wdata[39];
  assign T46[38] = io_rw_rdata[38] | io_rw_wdata[38];
  assign T46[37] = io_rw_rdata[37] | io_rw_wdata[37];
  assign T46[36] = io_rw_rdata[36] | io_rw_wdata[36];
  assign T46[35] = io_rw_rdata[35] | io_rw_wdata[35];
  assign T46[34] = io_rw_rdata[34] | io_rw_wdata[34];
  assign T46[33] = io_rw_rdata[33] | io_rw_wdata[33];
  assign T46[32] = io_rw_rdata[32] | io_rw_wdata[32];
  assign T46[31] = io_rw_rdata[31] | io_rw_wdata[31];
  assign T46[30] = io_rw_rdata[30] | io_rw_wdata[30];
  assign T46[29] = io_rw_rdata[29] | io_rw_wdata[29];
  assign T46[28] = io_rw_rdata[28] | io_rw_wdata[28];
  assign T46[27] = io_rw_rdata[27] | io_rw_wdata[27];
  assign T46[26] = io_rw_rdata[26] | io_rw_wdata[26];
  assign T46[25] = io_rw_rdata[25] | io_rw_wdata[25];
  assign T46[24] = io_rw_rdata[24] | io_rw_wdata[24];
  assign T46[23] = io_rw_rdata[23] | io_rw_wdata[23];
  assign T46[22] = io_rw_rdata[22] | io_rw_wdata[22];
  assign T46[21] = io_rw_rdata[21] | io_rw_wdata[21];
  assign T46[20] = io_rw_rdata[20] | io_rw_wdata[20];
  assign T46[19] = io_rw_rdata[19] | io_rw_wdata[19];
  assign T46[18] = io_rw_rdata[18] | io_rw_wdata[18];
  assign T46[17] = io_rw_rdata[17] | io_rw_wdata[17];
  assign T46[16] = io_rw_rdata[16] | io_rw_wdata[16];
  assign T46[15] = io_rw_rdata[15] | io_rw_wdata[15];
  assign T46[14] = io_rw_rdata[14] | io_rw_wdata[14];
  assign T46[13] = io_rw_rdata[13] | io_rw_wdata[13];
  assign T46[12] = io_rw_rdata[12] | io_rw_wdata[12];
  assign T46[11] = io_rw_rdata[11] | io_rw_wdata[11];
  assign T46[10] = io_rw_rdata[10] | io_rw_wdata[10];
  assign T46[9] = io_rw_rdata[9] | io_rw_wdata[9];
  assign T46[8] = io_rw_rdata[8] | io_rw_wdata[8];
  assign T46[7] = io_rw_rdata[7] | io_rw_wdata[7];
  assign T46[6] = io_rw_rdata[6] | io_rw_wdata[6];
  assign T46[5] = io_rw_rdata[5] | io_rw_wdata[5];
  assign T46[4] = io_rw_rdata[4] | io_rw_wdata[4];
  assign T46[3] = io_rw_rdata[3] | io_rw_wdata[3];
  assign T46[2] = io_rw_rdata[2] | io_rw_wdata[2];
  assign T46[1] = io_rw_rdata[1] | io_rw_wdata[1];
  assign T46[0] = io_rw_rdata[0] | io_rw_wdata[0];
  assign T48[63] = io_rw_rdata[63] & T49[63];
  assign T48[62] = io_rw_rdata[62] & T49[62];
  assign T48[61] = io_rw_rdata[61] & T49[61];
  assign T48[60] = io_rw_rdata[60] & T49[60];
  assign T48[59] = io_rw_rdata[59] & T49[59];
  assign T48[58] = io_rw_rdata[58] & T49[58];
  assign T48[57] = io_rw_rdata[57] & T49[57];
  assign T48[56] = io_rw_rdata[56] & T49[56];
  assign T48[55] = io_rw_rdata[55] & T49[55];
  assign T48[54] = io_rw_rdata[54] & T49[54];
  assign T48[53] = io_rw_rdata[53] & T49[53];
  assign T48[52] = io_rw_rdata[52] & T49[52];
  assign T48[51] = io_rw_rdata[51] & T49[51];
  assign T48[50] = io_rw_rdata[50] & T49[50];
  assign T48[49] = io_rw_rdata[49] & T49[49];
  assign T48[48] = io_rw_rdata[48] & T49[48];
  assign T48[47] = io_rw_rdata[47] & T49[47];
  assign T48[46] = io_rw_rdata[46] & T49[46];
  assign T48[45] = io_rw_rdata[45] & T49[45];
  assign T48[44] = io_rw_rdata[44] & T49[44];
  assign T48[43] = io_rw_rdata[43] & T49[43];
  assign T48[42] = io_rw_rdata[42] & T49[42];
  assign T48[41] = io_rw_rdata[41] & T49[41];
  assign T48[40] = io_rw_rdata[40] & T49[40];
  assign T48[39] = io_rw_rdata[39] & T49[39];
  assign T48[38] = io_rw_rdata[38] & T49[38];
  assign T48[37] = io_rw_rdata[37] & T49[37];
  assign T48[36] = io_rw_rdata[36] & T49[36];
  assign T48[35] = io_rw_rdata[35] & T49[35];
  assign T48[34] = io_rw_rdata[34] & T49[34];
  assign T48[33] = io_rw_rdata[33] & T49[33];
  assign T48[32] = io_rw_rdata[32] & T49[32];
  assign T48[31] = io_rw_rdata[31] & T49[31];
  assign T48[30] = io_rw_rdata[30] & T49[30];
  assign T48[29] = io_rw_rdata[29] & T49[29];
  assign T48[28] = io_rw_rdata[28] & T49[28];
  assign T48[27] = io_rw_rdata[27] & T49[27];
  assign T48[26] = io_rw_rdata[26] & T49[26];
  assign T48[25] = io_rw_rdata[25] & T49[25];
  assign T48[24] = io_rw_rdata[24] & T49[24];
  assign T48[23] = io_rw_rdata[23] & T49[23];
  assign T48[22] = io_rw_rdata[22] & T49[22];
  assign T48[21] = io_rw_rdata[21] & T49[21];
  assign T48[20] = io_rw_rdata[20] & T49[20];
  assign T48[19] = io_rw_rdata[19] & T49[19];
  assign T48[18] = io_rw_rdata[18] & T49[18];
  assign T48[17] = io_rw_rdata[17] & T49[17];
  assign T48[16] = io_rw_rdata[16] & T49[16];
  assign T48[15] = io_rw_rdata[15] & T49[15];
  assign T48[14] = io_rw_rdata[14] & T49[14];
  assign T48[13] = io_rw_rdata[13] & T49[13];
  assign T48[12] = io_rw_rdata[12] & T49[12];
  assign T48[11] = io_rw_rdata[11] & T49[11];
  assign T48[10] = io_rw_rdata[10] & T49[10];
  assign T48[9] = io_rw_rdata[9] & T49[9];
  assign T48[8] = io_rw_rdata[8] & T49[8];
  assign T48[7] = io_rw_rdata[7] & T49[7];
  assign T48[6] = io_rw_rdata[6] & T49[6];
  assign T48[5] = io_rw_rdata[5] & T49[5];
  assign T48[4] = io_rw_rdata[4] & T49[4];
  assign T48[3] = io_rw_rdata[3] & T49[3];
  assign T48[2] = io_rw_rdata[2] & T49[2];
  assign T48[1] = io_rw_rdata[1] & T49[1];
  assign T48[0] = io_rw_rdata[0] & T49[0];
  assign T49[63] = ~io_rw_wdata[63];
  assign T49[62] = ~io_rw_wdata[62];
  assign T49[61] = ~io_rw_wdata[61];
  assign T49[60] = ~io_rw_wdata[60];
  assign T49[59] = ~io_rw_wdata[59];
  assign T49[58] = ~io_rw_wdata[58];
  assign T49[57] = ~io_rw_wdata[57];
  assign T49[56] = ~io_rw_wdata[56];
  assign T49[55] = ~io_rw_wdata[55];
  assign T49[54] = ~io_rw_wdata[54];
  assign T49[53] = ~io_rw_wdata[53];
  assign T49[52] = ~io_rw_wdata[52];
  assign T49[51] = ~io_rw_wdata[51];
  assign T49[50] = ~io_rw_wdata[50];
  assign T49[49] = ~io_rw_wdata[49];
  assign T49[48] = ~io_rw_wdata[48];
  assign T49[47] = ~io_rw_wdata[47];
  assign T49[46] = ~io_rw_wdata[46];
  assign T49[45] = ~io_rw_wdata[45];
  assign T49[44] = ~io_rw_wdata[44];
  assign T49[43] = ~io_rw_wdata[43];
  assign T49[42] = ~io_rw_wdata[42];
  assign T49[41] = ~io_rw_wdata[41];
  assign T49[40] = ~io_rw_wdata[40];
  assign T49[39] = ~io_rw_wdata[39];
  assign T49[38] = ~io_rw_wdata[38];
  assign T49[37] = ~io_rw_wdata[37];
  assign T49[36] = ~io_rw_wdata[36];
  assign T49[35] = ~io_rw_wdata[35];
  assign T49[34] = ~io_rw_wdata[34];
  assign T49[33] = ~io_rw_wdata[33];
  assign T49[32] = ~io_rw_wdata[32];
  assign T49[31] = ~io_rw_wdata[31];
  assign T49[30] = ~io_rw_wdata[30];
  assign T49[29] = ~io_rw_wdata[29];
  assign T49[28] = ~io_rw_wdata[28];
  assign T49[27] = ~io_rw_wdata[27];
  assign T49[26] = ~io_rw_wdata[26];
  assign T49[25] = ~io_rw_wdata[25];
  assign T49[24] = ~io_rw_wdata[24];
  assign T49[23] = ~io_rw_wdata[23];
  assign T49[22] = ~io_rw_wdata[22];
  assign T49[21] = ~io_rw_wdata[21];
  assign T49[20] = ~io_rw_wdata[20];
  assign T49[19] = ~io_rw_wdata[19];
  assign T49[18] = ~io_rw_wdata[18];
  assign T49[17] = ~io_rw_wdata[17];
  assign T49[16] = ~io_rw_wdata[16];
  assign T49[15] = ~io_rw_wdata[15];
  assign T49[14] = ~io_rw_wdata[14];
  assign T49[13] = ~io_rw_wdata[13];
  assign T49[12] = ~io_rw_wdata[12];
  assign T49[11] = ~io_rw_wdata[11];
  assign T49[10] = ~io_rw_wdata[10];
  assign T49[9] = ~io_rw_wdata[9];
  assign T49[8] = ~io_rw_wdata[8];
  assign T49[7] = ~io_rw_wdata[7];
  assign T49[6] = ~io_rw_wdata[6];
  assign T49[5] = ~io_rw_wdata[5];
  assign T49[4] = ~io_rw_wdata[4];
  assign T49[3] = ~io_rw_wdata[3];
  assign T49[2] = ~io_rw_wdata[2];
  assign T49[1] = ~io_rw_wdata[1];
  assign T49[0] = ~io_rw_wdata[0];
  assign T52 = T58 & T53;
  assign T53 = T55 | N2299;
  assign T55 = N2310 | N2312;
  assign T58 = io_rocc_csr_wen & N2953;
  assign N163 = ~cpu_ren;
  assign io_rocc_csr_wen = T63 | T61;
  assign T61 = host_csr_req_fire & host_csr_bits_rw;
  assign T63 = cpu_wen & T64;
  assign T64 = ~N2394;
  assign cpu_wen = T66 & priv_sufficient;
  assign T66 = cpu_ren & N2399;
  assign T69 = T58 & T70;
  assign T70 = T72 | N2296;
  assign T72 = N2307 | N2309;
  assign T76 = io_rocc_csr_wen & N2527;
  assign T914[0] = T78 & priv_sufficient;
  assign T78 = T79 & N3100;
  assign T79 = T82 & T80;
  assign T80 = ~io_rw_addr[0];
  assign T82 = io_rw_addr[8] & T83;
  assign T83 = ~io_rw_addr[1];
  assign T216[0] = maybe_insn_redirect_trap & priv_sufficient;
  assign maybe_insn_redirect_trap = io_rw_addr[2] & N3100;
  assign T88 = T58 & T89;
  assign T89 = T91 | N2306;
  assign T91 = N2320 | N2322;
  assign T94 = T214 | T95;
  assign T95 = cpu_ren & T96;
  assign T96 = T104 | T97;
  assign T97 = fp_csr & T98;
  assign T98 = ~T99;
  assign fp_csr = T101 | N3073;
  assign T101 = N3085 | N3097;
  assign T104 = T213 | T105;
  assign T105 = ~addr_valid;
  assign addr_valid = T107 | N2413;
  assign T107 = T109 | N2426;
  assign T109 = T111 | N2439;
  assign T111 = T113 | N2451;
  assign T113 = T115 | N2466;
  assign T115 = T117 | N2478;
  assign T117 = T119 | N2490;
  assign T119 = T121 | N2503;
  assign T121 = T123 | N2515;
  assign T123 = T124 | N2527;
  assign T124 = T126 | N2540;
  assign T126 = T128 | N2552;
  assign T128 = T130 | N2564;
  assign T130 = T132 | N2576;
  assign T132 = T134 | N2588;
  assign T134 = T136 | N2600;
  assign T136 = T138 | N2612;
  assign T138 = T140 | N2624;
  assign T140 = T142 | N2636;
  assign T142 = T144 | N2648;
  assign T144 = T146 | N2660;
  assign T146 = T148 | N2672;
  assign T148 = T150 | N2684;
  assign T150 = T152 | N2696;
  assign T152 = T154 | N2708;
  assign T154 = T156 | N2720;
  assign T156 = T158 | N2732;
  assign T158 = T160 | N2744;
  assign T160 = T162 | N2757;
  assign T162 = T164 | N2769;
  assign T164 = T166 | N2781;
  assign T166 = T168 | N2794;
  assign T168 = T170 | N2809;
  assign T170 = T172 | N2821;
  assign T172 = T174 | N2833;
  assign T174 = T176 | N2845;
  assign T176 = T178 | N2857;
  assign T178 = T180 | N2869;
  assign T180 = T182 | N2881;
  assign T182 = T184 | N2893;
  assign T184 = T186 | N2905;
  assign T186 = T188 | N2917;
  assign T188 = T190 | N2929;
  assign T190 = T192 | N2941;
  assign T192 = T193 | N2953;
  assign T193 = T195 | N2965;
  assign T195 = T197 | N2977;
  assign T197 = T199 | N2989;
  assign T199 = T201 | N3001;
  assign T201 = T203 | N3013;
  assign T203 = T205 | N3025;
  assign T205 = T207 | N3037;
  assign T207 = T209 | N3049;
  assign T209 = T211 | N3061;
  assign T211 = T212 | N3073;
  assign T212 = N3085 | N3097;
  assign T213 = ~priv_sufficient;
  assign T214 = cpu_wen & N2394;
  assign N164 = ~T312;
  assign N165 = ~T300;
  assign T218[1] = T300;
  assign N166 = ~T285;
  assign N167 = ~T273;
  assign T220_0 = T273;
  assign N168 = ~T260;
  assign T222[63] = T223;
  assign T223 = T247 & T224;
  assign T224 = T246 | T225;
  assign T225 = N2319 & io_status_ie;
  assign T246 = ~N3101;
  assign N3101 = io_status_prv[1] | io_status_prv[0];
  assign T247 = T497_1 & T515_1;
  assign T251 = io_rocc_csr_wen & N2881;
  assign T253 = io_rocc_csr_wen & N2515;
  assign T257 = io_rocc_csr_wen & N2869;
  assign T259 = io_rocc_csr_wen & N2503;
  assign T260 = T265 & T261;
  assign T261 = T264 | T262;
  assign T262 = N2303 & io_status_ie;
  assign T265 = T848[3] & T858[3];
  assign T270 = io_rocc_csr_wen & N2893;
  assign T273 = T278 & T274;
  assign T274 = T277 | T275;
  assign T275 = N2293 & io_status_ie;
  assign T277 = ~N3102;
  assign N3102 = io_status_prv[1] | io_status_prv[0];
  assign T278 = T497[5] & T515[5];
  assign T285 = T290 & T286;
  assign T286 = T289 | T287;
  assign T287 = N2160 & io_status_ie;
  assign T290 = T848_7 & T858_7;
  assign T295 = io_rocc_csr_wen & N2989;
  assign T297 = io_rocc_csr_wen & N2809;
  assign T300 = N2385 & T301;
  assign T301 = T304 | T302;
  assign T302 = N2088 & io_status_ie;
  assign T307 = T311 & T308;
  assign T308 = N2152 | T309;
  assign T309 = ~host_csr_req_fire;
  assign T311 = io_rocc_csr_wen & N2757;
  assign T312 = io_rocc_interrupt & T313;
  assign T313 = T316 | T314;
  assign T314 = N2082 & io_status_ie;
  assign N169 = ~T322;
  assign N170 = ~T320;
  assign T320 = io_rocc_csr_wen & N3097;
  assign T322 = io_rocc_csr_wen & N3073;
  assign io_fatc = T331 & priv_sufficient;
  assign T331 = T332 & N3100;
  assign T332 = T334 & io_rw_addr[0];
  assign T334 = io_rw_addr[8] & T335;
  assign T335 = ~io_rw_addr[1];
  assign N171 = ~T369;
  assign N172 = ~maybe_insn_redirect_trap;
  assign N173 = ~io_status_prv[1];
  assign N174 = ~T346;
  assign N175 = ~T216[0];
  assign T343[39] = ~T344[39];
  assign T343[38] = ~T344[38];
  assign T343[37] = ~T344[37];
  assign T343[36] = ~T344[36];
  assign T343[35] = ~T344[35];
  assign T343[34] = ~T344[34];
  assign T343[33] = ~T344[33];
  assign T343[32] = ~T344[32];
  assign T343[31] = ~T344[31];
  assign T343[30] = ~T344[30];
  assign T343[29] = ~T344[29];
  assign T343[28] = ~T344[28];
  assign T343[27] = ~T344[27];
  assign T343[26] = ~T344[26];
  assign T343[25] = ~T344[25];
  assign T343[24] = ~T344[24];
  assign T343[23] = ~T344[23];
  assign T343[22] = ~T344[22];
  assign T343[21] = ~T344[21];
  assign T343[20] = ~T344[20];
  assign T343[19] = ~T344[19];
  assign T343[18] = ~T344[18];
  assign T343[17] = ~T344[17];
  assign T343[16] = ~T344[16];
  assign T343[15] = ~T344[15];
  assign T343[14] = ~T344[14];
  assign T343[13] = ~T344[13];
  assign T343[12] = ~T344[12];
  assign T343[11] = ~T344[11];
  assign T343[10] = ~T344[10];
  assign T343[9] = ~T344[9];
  assign T343[8] = ~T344[8];
  assign T343[7] = ~T344[7];
  assign T343[6] = ~T344[6];
  assign T343[5] = ~T344[5];
  assign T343[4] = ~T344[4];
  assign T343[3] = ~T344[3];
  assign T343[2] = ~T344[2];
  assign T343[1] = ~1'b1;
  assign T343[0] = ~1'b1;
  assign T344[39] = ~io_rocc_csr_wdata[39];
  assign T344[38] = ~io_rocc_csr_wdata[38];
  assign T344[37] = ~io_rocc_csr_wdata[37];
  assign T344[36] = ~io_rocc_csr_wdata[36];
  assign T344[35] = ~io_rocc_csr_wdata[35];
  assign T344[34] = ~io_rocc_csr_wdata[34];
  assign T344[33] = ~io_rocc_csr_wdata[33];
  assign T344[32] = ~io_rocc_csr_wdata[32];
  assign T344[31] = ~io_rocc_csr_wdata[31];
  assign T344[30] = ~io_rocc_csr_wdata[30];
  assign T344[29] = ~io_rocc_csr_wdata[29];
  assign T344[28] = ~io_rocc_csr_wdata[28];
  assign T344[27] = ~io_rocc_csr_wdata[27];
  assign T344[26] = ~io_rocc_csr_wdata[26];
  assign T344[25] = ~io_rocc_csr_wdata[25];
  assign T344[24] = ~io_rocc_csr_wdata[24];
  assign T344[23] = ~io_rocc_csr_wdata[23];
  assign T344[22] = ~io_rocc_csr_wdata[22];
  assign T344[21] = ~io_rocc_csr_wdata[21];
  assign T344[20] = ~io_rocc_csr_wdata[20];
  assign T344[19] = ~io_rocc_csr_wdata[19];
  assign T344[18] = ~io_rocc_csr_wdata[18];
  assign T344[17] = ~io_rocc_csr_wdata[17];
  assign T344[16] = ~io_rocc_csr_wdata[16];
  assign T344[15] = ~io_rocc_csr_wdata[15];
  assign T344[14] = ~io_rocc_csr_wdata[14];
  assign T344[13] = ~io_rocc_csr_wdata[13];
  assign T344[12] = ~io_rocc_csr_wdata[12];
  assign T344[11] = ~io_rocc_csr_wdata[11];
  assign T344[10] = ~io_rocc_csr_wdata[10];
  assign T344[9] = ~io_rocc_csr_wdata[9];
  assign T344[8] = ~io_rocc_csr_wdata[8];
  assign T344[7] = ~io_rocc_csr_wdata[7];
  assign T344[6] = ~io_rocc_csr_wdata[6];
  assign T344[5] = ~io_rocc_csr_wdata[5];
  assign T344[4] = ~io_rocc_csr_wdata[4];
  assign T344[3] = ~io_rocc_csr_wdata[3];
  assign T344[2] = ~io_rocc_csr_wdata[2];
  assign T346 = io_rocc_csr_wen & N2426;
  assign N176 = ~T355;
  assign N177 = ~T25;
  assign T349[39] = ~T350[39];
  assign T349[38] = ~T350[38];
  assign T349[37] = ~T350[37];
  assign T349[36] = ~T350[36];
  assign T349[35] = ~T350[35];
  assign T349[34] = ~T350[34];
  assign T349[33] = ~T350[33];
  assign T349[32] = ~T350[32];
  assign T349[31] = ~T350[31];
  assign T349[30] = ~T350[30];
  assign T349[29] = ~T350[29];
  assign T349[28] = ~T350[28];
  assign T349[27] = ~T350[27];
  assign T349[26] = ~T350[26];
  assign T349[25] = ~T350[25];
  assign T349[24] = ~T350[24];
  assign T349[23] = ~T350[23];
  assign T349[22] = ~T350[22];
  assign T349[21] = ~T350[21];
  assign T349[20] = ~T350[20];
  assign T349[19] = ~T350[19];
  assign T349[18] = ~T350[18];
  assign T349[17] = ~T350[17];
  assign T349[16] = ~T350[16];
  assign T349[15] = ~T350[15];
  assign T349[14] = ~T350[14];
  assign T349[13] = ~T350[13];
  assign T349[12] = ~T350[12];
  assign T349[11] = ~T350[11];
  assign T349[10] = ~T350[10];
  assign T349[9] = ~T350[9];
  assign T349[8] = ~T350[8];
  assign T349[7] = ~T350[7];
  assign T349[6] = ~T350[6];
  assign T349[5] = ~T350[5];
  assign T349[4] = ~T350[4];
  assign T349[3] = ~T350[3];
  assign T349[2] = ~T350[2];
  assign T349[1] = ~1'b1;
  assign T349[0] = ~1'b1;
  assign T350[39] = ~io_pc[39];
  assign T350[38] = ~io_pc[38];
  assign T350[37] = ~io_pc[37];
  assign T350[36] = ~io_pc[36];
  assign T350[35] = ~io_pc[35];
  assign T350[34] = ~io_pc[34];
  assign T350[33] = ~io_pc[33];
  assign T350[32] = ~io_pc[32];
  assign T350[31] = ~io_pc[31];
  assign T350[30] = ~io_pc[30];
  assign T350[29] = ~io_pc[29];
  assign T350[28] = ~io_pc[28];
  assign T350[27] = ~io_pc[27];
  assign T350[26] = ~io_pc[26];
  assign T350[25] = ~io_pc[25];
  assign T350[24] = ~io_pc[24];
  assign T350[23] = ~io_pc[23];
  assign T350[22] = ~io_pc[22];
  assign T350[21] = ~io_pc[21];
  assign T350[20] = ~io_pc[20];
  assign T350[19] = ~io_pc[19];
  assign T350[18] = ~io_pc[18];
  assign T350[17] = ~io_pc[17];
  assign T350[16] = ~io_pc[16];
  assign T350[15] = ~io_pc[15];
  assign T350[14] = ~io_pc[14];
  assign T350[13] = ~io_pc[13];
  assign T350[12] = ~io_pc[12];
  assign T350[11] = ~io_pc[11];
  assign T350[10] = ~io_pc[10];
  assign T350[9] = ~io_pc[9];
  assign T350[8] = ~io_pc[8];
  assign T350[7] = ~io_pc[7];
  assign T350[6] = ~io_pc[6];
  assign T350[5] = ~io_pc[5];
  assign T350[4] = ~io_pc[4];
  assign T350[3] = ~io_pc[3];
  assign T350[2] = ~io_pc[2];
  assign T352[39] = ~T353[39];
  assign T352[38] = ~T353[38];
  assign T352[37] = ~T353[37];
  assign T352[36] = ~T353[36];
  assign T352[35] = ~T353[35];
  assign T352[34] = ~T353[34];
  assign T352[33] = ~T353[33];
  assign T352[32] = ~T353[32];
  assign T352[31] = ~T353[31];
  assign T352[30] = ~T353[30];
  assign T352[29] = ~T353[29];
  assign T352[28] = ~T353[28];
  assign T352[27] = ~T353[27];
  assign T352[26] = ~T353[26];
  assign T352[25] = ~T353[25];
  assign T352[24] = ~T353[24];
  assign T352[23] = ~T353[23];
  assign T352[22] = ~T353[22];
  assign T352[21] = ~T353[21];
  assign T352[20] = ~T353[20];
  assign T352[19] = ~T353[19];
  assign T352[18] = ~T353[18];
  assign T352[17] = ~T353[17];
  assign T352[16] = ~T353[16];
  assign T352[15] = ~T353[15];
  assign T352[14] = ~T353[14];
  assign T352[13] = ~T353[13];
  assign T352[12] = ~T353[12];
  assign T352[11] = ~T353[11];
  assign T352[10] = ~T353[10];
  assign T352[9] = ~T353[9];
  assign T352[8] = ~T353[8];
  assign T352[7] = ~T353[7];
  assign T352[6] = ~T353[6];
  assign T352[5] = ~T353[5];
  assign T352[4] = ~T353[4];
  assign T352[3] = ~T353[3];
  assign T352[2] = ~T353[2];
  assign T352[1] = ~1'b1;
  assign T352[0] = ~1'b1;
  assign T353[39] = ~io_rocc_csr_wdata[39];
  assign T353[38] = ~io_rocc_csr_wdata[38];
  assign T353[37] = ~io_rocc_csr_wdata[37];
  assign T353[36] = ~io_rocc_csr_wdata[36];
  assign T353[35] = ~io_rocc_csr_wdata[35];
  assign T353[34] = ~io_rocc_csr_wdata[34];
  assign T353[33] = ~io_rocc_csr_wdata[33];
  assign T353[32] = ~io_rocc_csr_wdata[32];
  assign T353[31] = ~io_rocc_csr_wdata[31];
  assign T353[30] = ~io_rocc_csr_wdata[30];
  assign T353[29] = ~io_rocc_csr_wdata[29];
  assign T353[28] = ~io_rocc_csr_wdata[28];
  assign T353[27] = ~io_rocc_csr_wdata[27];
  assign T353[26] = ~io_rocc_csr_wdata[26];
  assign T353[25] = ~io_rocc_csr_wdata[25];
  assign T353[24] = ~io_rocc_csr_wdata[24];
  assign T353[23] = ~io_rocc_csr_wdata[23];
  assign T353[22] = ~io_rocc_csr_wdata[22];
  assign T353[21] = ~io_rocc_csr_wdata[21];
  assign T353[20] = ~io_rocc_csr_wdata[20];
  assign T353[19] = ~io_rocc_csr_wdata[19];
  assign T353[18] = ~io_rocc_csr_wdata[18];
  assign T353[17] = ~io_rocc_csr_wdata[17];
  assign T353[16] = ~io_rocc_csr_wdata[16];
  assign T353[15] = ~io_rocc_csr_wdata[15];
  assign T353[14] = ~io_rocc_csr_wdata[14];
  assign T353[13] = ~io_rocc_csr_wdata[13];
  assign T353[12] = ~io_rocc_csr_wdata[12];
  assign T353[11] = ~io_rocc_csr_wdata[11];
  assign T353[10] = ~io_rocc_csr_wdata[10];
  assign T353[9] = ~io_rocc_csr_wdata[9];
  assign T353[8] = ~io_rocc_csr_wdata[8];
  assign T353[7] = ~io_rocc_csr_wdata[7];
  assign T353[6] = ~io_rocc_csr_wdata[6];
  assign T353[5] = ~io_rocc_csr_wdata[5];
  assign T353[4] = ~io_rocc_csr_wdata[4];
  assign T353[3] = ~io_rocc_csr_wdata[3];
  assign T353[2] = ~io_rocc_csr_wdata[2];
  assign T355 = io_rocc_csr_wen & N2845;
  assign N178 = ~T362;
  assign T359[38] = ~T360[38];
  assign T359[37] = ~T360[37];
  assign T359[36] = ~T360[36];
  assign T359[35] = ~T360[35];
  assign T359[34] = ~T360[34];
  assign T359[33] = ~T360[33];
  assign T359[32] = ~T360[32];
  assign T359[31] = ~T360[31];
  assign T359[30] = ~T360[30];
  assign T359[29] = ~T360[29];
  assign T359[28] = ~T360[28];
  assign T359[27] = ~T360[27];
  assign T359[26] = ~T360[26];
  assign T359[25] = ~T360[25];
  assign T359[24] = ~T360[24];
  assign T359[23] = ~T360[23];
  assign T359[22] = ~T360[22];
  assign T359[21] = ~T360[21];
  assign T359[20] = ~T360[20];
  assign T359[19] = ~T360[19];
  assign T359[18] = ~T360[18];
  assign T359[17] = ~T360[17];
  assign T359[16] = ~T360[16];
  assign T359[15] = ~T360[15];
  assign T359[14] = ~T360[14];
  assign T359[13] = ~T360[13];
  assign T359[12] = ~T360[12];
  assign T359[11] = ~T360[11];
  assign T359[10] = ~T360[10];
  assign T359[9] = ~T360[9];
  assign T359[8] = ~T360[8];
  assign T359[7] = ~T360[7];
  assign T359[6] = ~T360[6];
  assign T359[5] = ~T360[5];
  assign T359[4] = ~T360[4];
  assign T359[3] = ~T360[3];
  assign T359[2] = ~T360[2];
  assign T359[1] = ~1'b1;
  assign T359[0] = ~1'b1;
  assign T360[38] = ~io_rocc_csr_wdata[38];
  assign T360[37] = ~io_rocc_csr_wdata[37];
  assign T360[36] = ~io_rocc_csr_wdata[36];
  assign T360[35] = ~io_rocc_csr_wdata[35];
  assign T360[34] = ~io_rocc_csr_wdata[34];
  assign T360[33] = ~io_rocc_csr_wdata[33];
  assign T360[32] = ~io_rocc_csr_wdata[32];
  assign T360[31] = ~io_rocc_csr_wdata[31];
  assign T360[30] = ~io_rocc_csr_wdata[30];
  assign T360[29] = ~io_rocc_csr_wdata[29];
  assign T360[28] = ~io_rocc_csr_wdata[28];
  assign T360[27] = ~io_rocc_csr_wdata[27];
  assign T360[26] = ~io_rocc_csr_wdata[26];
  assign T360[25] = ~io_rocc_csr_wdata[25];
  assign T360[24] = ~io_rocc_csr_wdata[24];
  assign T360[23] = ~io_rocc_csr_wdata[23];
  assign T360[22] = ~io_rocc_csr_wdata[22];
  assign T360[21] = ~io_rocc_csr_wdata[21];
  assign T360[20] = ~io_rocc_csr_wdata[20];
  assign T360[19] = ~io_rocc_csr_wdata[19];
  assign T360[18] = ~io_rocc_csr_wdata[18];
  assign T360[17] = ~io_rocc_csr_wdata[17];
  assign T360[16] = ~io_rocc_csr_wdata[16];
  assign T360[15] = ~io_rocc_csr_wdata[15];
  assign T360[14] = ~io_rocc_csr_wdata[14];
  assign T360[13] = ~io_rocc_csr_wdata[13];
  assign T360[12] = ~io_rocc_csr_wdata[12];
  assign T360[11] = ~io_rocc_csr_wdata[11];
  assign T360[10] = ~io_rocc_csr_wdata[10];
  assign T360[9] = ~io_rocc_csr_wdata[9];
  assign T360[8] = ~io_rocc_csr_wdata[8];
  assign T360[7] = ~io_rocc_csr_wdata[7];
  assign T360[6] = ~io_rocc_csr_wdata[6];
  assign T360[5] = ~io_rocc_csr_wdata[5];
  assign T360[4] = ~io_rocc_csr_wdata[4];
  assign T360[3] = ~io_rocc_csr_wdata[3];
  assign T360[2] = ~io_rocc_csr_wdata[2];
  assign T362 = io_rocc_csr_wen & N2413;
  assign T367 = io_rocc_csr_wen & N2917;
  assign T369 = io_exception | io_csr_xcpt;
  assign T373 = io_rocc_csr_wen & N2451;
  assign T399 = T58 & N2087;
  assign T402 = T58 & N2159;
  assign io_status_sd = T409 | T408;
  assign io_eret = T914[0] | T216[0];
  assign insn_wfi = T413 & priv_sufficient;
  assign T413 = T414 & N3100;
  assign T414 = T417 & T415;
  assign T415 = ~io_rw_addr[0];
  assign T417 = io_rw_addr[8] & io_rw_addr[1];
  assign N179 = ~T435;
  assign N180 = ~T433;
  assign N181 = ~T431;
  assign N182 = ~T429;
  assign N183 = ~T427;
  assign T425 = T247 & T426;
  assign T427 = T265 & T428;
  assign T429 = T278 & T430;
  assign T431 = T290 & T432;
  assign T433 = N2385 & T434;
  assign T435 = io_rocc_interrupt & T436;
  assign io_rw_rdata[63] = T442[63] | T438[63];
  assign io_rw_rdata[62] = T442[62] | T438[62];
  assign io_rw_rdata[61] = T442[61] | T438[61];
  assign io_rw_rdata[60] = T442[60] | T438[60];
  assign io_rw_rdata[59] = T442[59] | T438[59];
  assign io_rw_rdata[58] = T442[58] | T438[58];
  assign io_rw_rdata[57] = T442[57] | T438[57];
  assign io_rw_rdata[56] = T442[56] | T438[56];
  assign io_rw_rdata[55] = T442[55] | T438[55];
  assign io_rw_rdata[54] = T442[54] | T438[54];
  assign io_rw_rdata[53] = T442[53] | T438[53];
  assign io_rw_rdata[52] = T442[52] | T438[52];
  assign io_rw_rdata[51] = T442[51] | T438[51];
  assign io_rw_rdata[50] = T442[50] | T438[50];
  assign io_rw_rdata[49] = T442[49] | T438[49];
  assign io_rw_rdata[48] = T442[48] | T438[48];
  assign io_rw_rdata[47] = T442[47] | T438[47];
  assign io_rw_rdata[46] = T442[46] | T438[46];
  assign io_rw_rdata[45] = T442[45] | T438[45];
  assign io_rw_rdata[44] = T442[44] | T438[44];
  assign io_rw_rdata[43] = T442[43] | T438[43];
  assign io_rw_rdata[42] = T442[42] | T438[42];
  assign io_rw_rdata[41] = T442[41] | T438[41];
  assign io_rw_rdata[40] = T442[40] | T438[40];
  assign io_rw_rdata[39] = T442[39] | T438[39];
  assign io_rw_rdata[38] = T442[38] | T438[38];
  assign io_rw_rdata[37] = T442[37] | T438[37];
  assign io_rw_rdata[36] = T442[36] | T438[36];
  assign io_rw_rdata[35] = T442[35] | T438[35];
  assign io_rw_rdata[34] = T442[34] | T438[34];
  assign io_rw_rdata[33] = T442[33] | T438[33];
  assign io_rw_rdata[32] = T442[32] | T438[32];
  assign io_rw_rdata[31] = T442[31] | T438[31];
  assign io_rw_rdata[30] = T442[30] | T438[30];
  assign io_rw_rdata[29] = T442[29] | T438[29];
  assign io_rw_rdata[28] = T442[28] | T438[28];
  assign io_rw_rdata[27] = T442[27] | T438[27];
  assign io_rw_rdata[26] = T442[26] | T438[26];
  assign io_rw_rdata[25] = T442[25] | T438[25];
  assign io_rw_rdata[24] = T442[24] | T438[24];
  assign io_rw_rdata[23] = T442[23] | T438[23];
  assign io_rw_rdata[22] = T442[22] | T438[22];
  assign io_rw_rdata[21] = T442[21] | T438[21];
  assign io_rw_rdata[20] = T442[20] | T438[20];
  assign io_rw_rdata[19] = T442[19] | T438[19];
  assign io_rw_rdata[18] = T442[18] | T438[18];
  assign io_rw_rdata[17] = T442[17] | T438[17];
  assign io_rw_rdata[16] = T442[16] | T438[16];
  assign io_rw_rdata[15] = T442[15] | T438[15];
  assign io_rw_rdata[14] = T442[14] | T438[14];
  assign io_rw_rdata[13] = T442[13] | T438[13];
  assign io_rw_rdata[12] = T442[12] | T438[12];
  assign io_rw_rdata[11] = T442[11] | T438[11];
  assign io_rw_rdata[10] = T442[10] | T438[10];
  assign io_rw_rdata[9] = T442[9] | T438[9];
  assign io_rw_rdata[8] = T442[8] | T438[8];
  assign io_rw_rdata[7] = T442[7] | T438[7];
  assign io_rw_rdata[6] = T442[6] | T438[6];
  assign io_rw_rdata[5] = T442[5] | T438[5];
  assign io_rw_rdata[4] = T442[4] | T438[4];
  assign io_rw_rdata[3] = T442[3] | T438[3];
  assign io_rw_rdata[2] = T442[2] | T438[2];
  assign io_rw_rdata[1] = T442[1] | T438[1];
  assign io_rw_rdata[0] = T442[0] | T438[0];
  assign T442[63] = T447[63] | T443[63];
  assign T442[62] = T447[62] | T443[62];
  assign T442[61] = T447[61] | T443[61];
  assign T442[60] = T447[60] | T443[60];
  assign T442[59] = T447[59] | T443[59];
  assign T442[58] = T447[58] | T443[58];
  assign T442[57] = T447[57] | T443[57];
  assign T442[56] = T447[56] | T443[56];
  assign T442[55] = T447[55] | T443[55];
  assign T442[54] = T447[54] | T443[54];
  assign T442[53] = T447[53] | T443[53];
  assign T442[52] = T447[52] | T443[52];
  assign T442[51] = T447[51] | T443[51];
  assign T442[50] = T447[50] | T443[50];
  assign T442[49] = T447[49] | T443[49];
  assign T442[48] = T447[48] | T443[48];
  assign T442[47] = T447[47] | T443[47];
  assign T442[46] = T447[46] | T443[46];
  assign T442[45] = T447[45] | T443[45];
  assign T442[44] = T447[44] | T443[44];
  assign T442[43] = T447[43] | T443[43];
  assign T442[42] = T447[42] | T443[42];
  assign T442[41] = T447[41] | T443[41];
  assign T442[40] = T447[40] | T443[40];
  assign T442[39] = T447[39] | T443[39];
  assign T442[38] = T447[38] | T443[38];
  assign T442[37] = T447[37] | T443[37];
  assign T442[36] = T447[36] | T443[36];
  assign T442[35] = T447[35] | T443[35];
  assign T442[34] = T447[34] | T443[34];
  assign T442[33] = T447[33] | T443[33];
  assign T442[32] = T447[32] | T443[32];
  assign T442[31] = T447[31] | T443[31];
  assign T442[30] = T447[30] | T443[30];
  assign T442[29] = T447[29] | T443[29];
  assign T442[28] = T447[28] | T443[28];
  assign T442[27] = T447[27] | T443[27];
  assign T442[26] = T447[26] | T443[26];
  assign T442[25] = T447[25] | T443[25];
  assign T442[24] = T447[24] | T443[24];
  assign T442[23] = T447[23] | T443[23];
  assign T442[22] = T447[22] | T443[22];
  assign T442[21] = T447[21] | T443[21];
  assign T442[20] = T447[20] | T443[20];
  assign T442[19] = T447[19] | T443[19];
  assign T442[18] = T447[18] | T443[18];
  assign T442[17] = T447[17] | T443[17];
  assign T442[16] = T447[16] | T443[16];
  assign T442[15] = T447[15] | T443[15];
  assign T442[14] = T447[14] | T443[14];
  assign T442[13] = T447[13] | T443[13];
  assign T442[12] = T447[12] | T443[12];
  assign T442[11] = T447[11] | T443[11];
  assign T442[10] = T447[10] | T443[10];
  assign T442[9] = T447[9] | T443[9];
  assign T442[8] = T447[8] | T443[8];
  assign T442[7] = T447[7] | T443[7];
  assign T442[6] = T447[6] | T443[6];
  assign T442[5] = T447[5] | T443[5];
  assign T442[4] = T447[4] | T443[4];
  assign T442[3] = T447[3] | T443[3];
  assign T442[2] = T447[2] | T443[2];
  assign T442[1] = T447[1] | T443[1];
  assign T442[0] = T447[0] | T443[0];
  assign T447[63] = T450[63] | 1'b0;
  assign T447[62] = T450[62] | 1'b0;
  assign T447[61] = T450[61] | 1'b0;
  assign T447[60] = T450[60] | 1'b0;
  assign T447[59] = T450[59] | 1'b0;
  assign T447[58] = T450[58] | 1'b0;
  assign T447[57] = T450[57] | 1'b0;
  assign T447[56] = T450[56] | 1'b0;
  assign T447[55] = T450[55] | 1'b0;
  assign T447[54] = T450[54] | 1'b0;
  assign T447[53] = T450[53] | 1'b0;
  assign T447[52] = T450[52] | 1'b0;
  assign T447[51] = T450[51] | 1'b0;
  assign T447[50] = T450[50] | 1'b0;
  assign T447[49] = T450[49] | 1'b0;
  assign T447[48] = T450[48] | 1'b0;
  assign T447[47] = T450[47] | 1'b0;
  assign T447[46] = T450[46] | 1'b0;
  assign T447[45] = T450[45] | 1'b0;
  assign T447[44] = T450[44] | 1'b0;
  assign T447[43] = T450[43] | 1'b0;
  assign T447[42] = T450[42] | 1'b0;
  assign T447[41] = T450[41] | 1'b0;
  assign T447[40] = T450[40] | 1'b0;
  assign T447[39] = T450[39] | 1'b0;
  assign T447[38] = T450[38] | 1'b0;
  assign T447[37] = T450[37] | 1'b0;
  assign T447[36] = T450[36] | 1'b0;
  assign T447[35] = T450[35] | 1'b0;
  assign T447[34] = T450[34] | 1'b0;
  assign T447[33] = T450[33] | 1'b0;
  assign T447[32] = T450[32] | 1'b0;
  assign T447[31] = T450[31] | T945[31];
  assign T447[30] = T450[30] | T945[30];
  assign T447[29] = T450[29] | T945[29];
  assign T447[28] = T450[28] | T945[28];
  assign T447[27] = T450[27] | T945[27];
  assign T447[26] = T450[26] | T945[26];
  assign T447[25] = T450[25] | T945[25];
  assign T447[24] = T450[24] | T945[24];
  assign T447[23] = T450[23] | T945[23];
  assign T447[22] = T450[22] | T945[22];
  assign T447[21] = T450[21] | T945[21];
  assign T447[20] = T450[20] | T945[20];
  assign T447[19] = T450[19] | T945[19];
  assign T447[18] = T450[18] | T945[18];
  assign T447[17] = T450[17] | T945[17];
  assign T447[16] = T450[16] | T945[16];
  assign T447[15] = T450[15] | T945[15];
  assign T447[14] = T450[14] | T945[14];
  assign T447[13] = T450[13] | T945[13];
  assign T447[12] = T450[12] | T945[12];
  assign T447[11] = T450[11] | T945[11];
  assign T447[10] = T450[10] | T945[10];
  assign T447[9] = T450[9] | T945[9];
  assign T447[8] = T450[8] | T945[8];
  assign T447[7] = T450[7] | T945[7];
  assign T447[6] = T450[6] | T945[6];
  assign T447[5] = T450[5] | T945[5];
  assign T447[4] = T450[4] | T945[4];
  assign T447[3] = T450[3] | T945[3];
  assign T447[2] = T450[2] | T945[2];
  assign T447[1] = T450[1] | T945[1];
  assign T447[0] = T450[0] | T945[0];
  assign T450[63] = T477[63] | T451[63];
  assign T450[62] = T477[62] | T451[62];
  assign T450[61] = T477[61] | T451[61];
  assign T450[60] = T477[60] | T451[60];
  assign T450[59] = T477[59] | T451[59];
  assign T450[58] = T477[58] | T451[58];
  assign T450[57] = T477[57] | T451[57];
  assign T450[56] = T477[56] | T451[56];
  assign T450[55] = T477[55] | T451[55];
  assign T450[54] = T477[54] | T451[54];
  assign T450[53] = T477[53] | T451[53];
  assign T450[52] = T477[52] | T451[52];
  assign T450[51] = T477[51] | T451[51];
  assign T450[50] = T477[50] | T451[50];
  assign T450[49] = T477[49] | T451[49];
  assign T450[48] = T477[48] | T451[48];
  assign T450[47] = T477[47] | T451[47];
  assign T450[46] = T477[46] | T451[46];
  assign T450[45] = T477[45] | T451[45];
  assign T450[44] = T477[44] | T451[44];
  assign T450[43] = T477[43] | T451[43];
  assign T450[42] = T477[42] | T451[42];
  assign T450[41] = T477[41] | T451[41];
  assign T450[40] = T477[40] | T451[40];
  assign T450[39] = T477[39] | T451[39];
  assign T450[38] = T477[38] | T451[38];
  assign T450[37] = T477[37] | T451[37];
  assign T450[36] = T477[36] | T451[36];
  assign T450[35] = T477[35] | T451[35];
  assign T450[34] = T477[34] | T451[34];
  assign T450[33] = T477[33] | T451[33];
  assign T450[32] = T477[32] | T451[32];
  assign T450[31] = T477[31] | T451[31];
  assign T450[30] = T477[30] | T451[30];
  assign T450[29] = T477[29] | T451[29];
  assign T450[28] = T477[28] | T451[28];
  assign T450[27] = T477[27] | T451[27];
  assign T450[26] = T477[26] | T451[26];
  assign T450[25] = T477[25] | T451[25];
  assign T450[24] = T477[24] | T451[24];
  assign T450[23] = T477[23] | T451[23];
  assign T450[22] = T477[22] | T451[22];
  assign T450[21] = T477[21] | T451[21];
  assign T450[20] = T477[20] | T451[20];
  assign T450[19] = T477[19] | T451[19];
  assign T450[18] = T477[18] | T451[18];
  assign T450[17] = T477[17] | T451[17];
  assign T450[16] = T477[16] | T451[16];
  assign T450[15] = T477[15] | T451[15];
  assign T450[14] = T477[14] | T451[14];
  assign T450[13] = T477[13] | T451[13];
  assign T450[12] = T477[12] | T451[12];
  assign T450[11] = T477[11] | T451[11];
  assign T450[10] = T477[10] | T451[10];
  assign T450[9] = T477[9] | T451[9];
  assign T450[8] = T477[8] | T451[8];
  assign T450[7] = T477[7] | T451[7];
  assign T450[6] = T477[6] | T451[6];
  assign T450[5] = T477[5] | T451[5];
  assign T450[4] = T477[4] | T451[4];
  assign T450[3] = T477[3] | T451[3];
  assign T450[2] = T477[2] | T451[2];
  assign T450[1] = T477[1] | T451[1];
  assign T450[0] = T477[0] | T451[0];
  assign N184 = ~T463;
  assign T465 = T25 & T466;
  assign T466 = T468 | N2226;
  assign T468 = T470 | N2302;
  assign T470 = N2315 | N2317;
  assign T474 = io_rocc_csr_wen & N2833;
  assign T477[63] = T491[63] | T478[63];
  assign T477[62] = T491[62] | T478[62];
  assign T477[61] = T491[61] | T478[61];
  assign T477[60] = T491[60] | T478[60];
  assign T477[59] = T491[59] | T478[59];
  assign T477[58] = T491[58] | T478[58];
  assign T477[57] = T491[57] | T478[57];
  assign T477[56] = T491[56] | T478[56];
  assign T477[55] = T491[55] | T478[55];
  assign T477[54] = T491[54] | T478[54];
  assign T477[53] = T491[53] | T478[53];
  assign T477[52] = T491[52] | T478[52];
  assign T477[51] = T491[51] | T478[51];
  assign T477[50] = T491[50] | T478[50];
  assign T477[49] = T491[49] | T478[49];
  assign T477[48] = T491[48] | T478[48];
  assign T477[47] = T491[47] | T478[47];
  assign T477[46] = T491[46] | T478[46];
  assign T477[45] = T491[45] | T478[45];
  assign T477[44] = T491[44] | T478[44];
  assign T477[43] = T491[43] | T478[43];
  assign T477[42] = T491[42] | T478[42];
  assign T477[41] = T491[41] | T478[41];
  assign T477[40] = T491[40] | T478[40];
  assign T477[39] = T491[39] | T478[39];
  assign T477[38] = T491[38] | T478[38];
  assign T477[37] = T491[37] | T478[37];
  assign T477[36] = T491[36] | T478[36];
  assign T477[35] = T491[35] | T478[35];
  assign T477[34] = T491[34] | T478[34];
  assign T477[33] = T491[33] | T478[33];
  assign T477[32] = T491[32] | T478[32];
  assign T477[31] = T491[31] | T478[31];
  assign T477[30] = T491[30] | T478[30];
  assign T477[29] = T491[29] | T478[29];
  assign T477[28] = T491[28] | T478[28];
  assign T477[27] = T491[27] | T478[27];
  assign T477[26] = T491[26] | T478[26];
  assign T477[25] = T491[25] | T478[25];
  assign T477[24] = T491[24] | T478[24];
  assign T477[23] = T491[23] | T478[23];
  assign T477[22] = T491[22] | T478[22];
  assign T477[21] = T491[21] | T478[21];
  assign T477[20] = T491[20] | T478[20];
  assign T477[19] = T491[19] | T478[19];
  assign T477[18] = T491[18] | T478[18];
  assign T477[17] = T491[17] | T478[17];
  assign T477[16] = T491[16] | T478[16];
  assign T477[15] = T491[15] | T478[15];
  assign T477[14] = T491[14] | T478[14];
  assign T477[13] = T491[13] | T478[13];
  assign T477[12] = T491[12] | T478[12];
  assign T477[11] = T491[11] | T478[11];
  assign T477[10] = T491[10] | T478[10];
  assign T477[9] = T491[9] | T478[9];
  assign T477[8] = T491[8] | T478[8];
  assign T477[7] = T491[7] | T478[7];
  assign T477[6] = T491[6] | T478[6];
  assign T477[5] = T491[5] | T478[5];
  assign T477[4] = T491[4] | T478[4];
  assign T477[3] = T491[3] | T478[3];
  assign T477[2] = T491[2] | T478[2];
  assign T477[1] = T491[1] | T478[1];
  assign T477[0] = T491[0] | T478[0];
  assign T485 = T25 & io_csr_xcpt;
  assign T486 = T485 & insn_break;
  assign T488 = T485 & insn_call;
  assign T490 = io_rocc_csr_wen & N2821;
  assign T491[63] = T495[63] | T492[63];
  assign T491[62] = T495[62] | T492[62];
  assign T491[61] = T495[61] | T492[61];
  assign T491[60] = T495[60] | T492[60];
  assign T491[59] = T495[59] | T492[59];
  assign T491[58] = T495[58] | T492[58];
  assign T491[57] = T495[57] | T492[57];
  assign T491[56] = T495[56] | T492[56];
  assign T491[55] = T495[55] | T492[55];
  assign T491[54] = T495[54] | T492[54];
  assign T491[53] = T495[53] | T492[53];
  assign T491[52] = T495[52] | T492[52];
  assign T491[51] = T495[51] | T492[51];
  assign T491[50] = T495[50] | T492[50];
  assign T491[49] = T495[49] | T492[49];
  assign T491[48] = T495[48] | T492[48];
  assign T491[47] = T495[47] | T492[47];
  assign T491[46] = T495[46] | T492[46];
  assign T491[45] = T495[45] | T492[45];
  assign T491[44] = T495[44] | T492[44];
  assign T491[43] = T495[43] | T492[43];
  assign T491[42] = T495[42] | T492[42];
  assign T491[41] = T495[41] | T492[41];
  assign T491[40] = T495[40] | T492[40];
  assign T491[39] = T495[39] | T492[39];
  assign T491[38] = T495[38] | T492[38];
  assign T491[37] = T495[37] | T492[37];
  assign T491[36] = T495[36] | T492[36];
  assign T491[35] = T495[35] | T492[35];
  assign T491[34] = T495[34] | T492[34];
  assign T491[33] = T495[33] | T492[33];
  assign T491[32] = T495[32] | T492[32];
  assign T491[31] = T495[31] | T492[31];
  assign T491[30] = T495[30] | T492[30];
  assign T491[29] = T495[29] | T492[29];
  assign T491[28] = T495[28] | T492[28];
  assign T491[27] = T495[27] | T492[27];
  assign T491[26] = T495[26] | T492[26];
  assign T491[25] = T495[25] | T492[25];
  assign T491[24] = T495[24] | T492[24];
  assign T491[23] = T495[23] | T492[23];
  assign T491[22] = T495[22] | T492[22];
  assign T491[21] = T495[21] | T492[21];
  assign T491[20] = T495[20] | T492[20];
  assign T491[19] = T495[19] | T492[19];
  assign T491[18] = T495[18] | T492[18];
  assign T491[17] = T495[17] | T492[17];
  assign T491[16] = T495[16] | T492[16];
  assign T491[15] = T495[15] | T492[15];
  assign T491[14] = T495[14] | T492[14];
  assign T491[13] = T495[13] | T492[13];
  assign T491[12] = T495[12] | T492[12];
  assign T491[11] = T495[11] | T492[11];
  assign T491[10] = T495[10] | T492[10];
  assign T491[9] = T495[9] | T492[9];
  assign T491[8] = T495[8] | T492[8];
  assign T491[7] = T495[7] | T492[7];
  assign T491[6] = T495[6] | T492[6];
  assign T491[5] = T495[5] | T492[5];
  assign T491[4] = T495[4] | T492[4];
  assign T491[3] = T495[3] | T492[3];
  assign T491[2] = T495[2] | T492[2];
  assign T491[1] = T495[1] | T492[1];
  assign T491[0] = T495[0] | T492[0];
  assign T494 = io_rocc_csr_wen & N2490;
  assign T495[63] = T513[63] | 1'b0;
  assign T495[62] = T513[62] | 1'b0;
  assign T495[61] = T513[61] | 1'b0;
  assign T495[60] = T513[60] | 1'b0;
  assign T495[59] = T513[59] | 1'b0;
  assign T495[58] = T513[58] | 1'b0;
  assign T495[57] = T513[57] | 1'b0;
  assign T495[56] = T513[56] | 1'b0;
  assign T495[55] = T513[55] | 1'b0;
  assign T495[54] = T513[54] | 1'b0;
  assign T495[53] = T513[53] | 1'b0;
  assign T495[52] = T513[52] | 1'b0;
  assign T495[51] = T513[51] | 1'b0;
  assign T495[50] = T513[50] | 1'b0;
  assign T495[49] = T513[49] | 1'b0;
  assign T495[48] = T513[48] | 1'b0;
  assign T495[47] = T513[47] | 1'b0;
  assign T495[46] = T513[46] | 1'b0;
  assign T495[45] = T513[45] | 1'b0;
  assign T495[44] = T513[44] | 1'b0;
  assign T495[43] = T513[43] | 1'b0;
  assign T495[42] = T513[42] | 1'b0;
  assign T495[41] = T513[41] | 1'b0;
  assign T495[40] = T513[40] | 1'b0;
  assign T495[39] = T513[39] | 1'b0;
  assign T495[38] = T513[38] | 1'b0;
  assign T495[37] = T513[37] | 1'b0;
  assign T495[36] = T513[36] | 1'b0;
  assign T495[35] = T513[35] | 1'b0;
  assign T495[34] = T513[34] | 1'b0;
  assign T495[33] = T513[33] | 1'b0;
  assign T495[32] = T513[32] | 1'b0;
  assign T495[31] = T513[31] | 1'b0;
  assign T495[30] = T513[30] | 1'b0;
  assign T495[29] = T513[29] | 1'b0;
  assign T495[28] = T513[28] | 1'b0;
  assign T495[27] = T513[27] | 1'b0;
  assign T495[26] = T513[26] | 1'b0;
  assign T495[25] = T513[25] | 1'b0;
  assign T495[24] = T513[24] | 1'b0;
  assign T495[23] = T513[23] | 1'b0;
  assign T495[22] = T513[22] | 1'b0;
  assign T495[21] = T513[21] | 1'b0;
  assign T495[20] = T513[20] | 1'b0;
  assign T495[19] = T513[19] | 1'b0;
  assign T495[18] = T513[18] | 1'b0;
  assign T495[17] = T513[17] | 1'b0;
  assign T495[16] = T513[16] | 1'b0;
  assign T495[15] = T513[15] | 1'b0;
  assign T495[14] = T513[14] | 1'b0;
  assign T495[13] = T513[13] | 1'b0;
  assign T495[12] = T513[12] | 1'b0;
  assign T495[11] = T513[11] | 1'b0;
  assign T495[10] = T513[10] | 1'b0;
  assign T495[9] = T513[9] | 1'b0;
  assign T495[8] = T513[8] | 1'b0;
  assign T495[7] = T513[7] | 1'b0;
  assign T495[6] = T513[6] | 1'b0;
  assign T495[5] = T513[5] | T949[5];
  assign T495[4] = T513[4] | 1'b0;
  assign T495[3] = T513[3] | 1'b0;
  assign T495[2] = T513[2] | 1'b0;
  assign T495[1] = T513[1] | T949_1;
  assign T495[0] = T513[0] | 1'b0;
  assign T513[63] = T531[63] | 1'b0;
  assign T513[62] = T531[62] | 1'b0;
  assign T513[61] = T531[61] | 1'b0;
  assign T513[60] = T531[60] | 1'b0;
  assign T513[59] = T531[59] | 1'b0;
  assign T513[58] = T531[58] | 1'b0;
  assign T513[57] = T531[57] | 1'b0;
  assign T513[56] = T531[56] | 1'b0;
  assign T513[55] = T531[55] | 1'b0;
  assign T513[54] = T531[54] | 1'b0;
  assign T513[53] = T531[53] | 1'b0;
  assign T513[52] = T531[52] | 1'b0;
  assign T513[51] = T531[51] | 1'b0;
  assign T513[50] = T531[50] | 1'b0;
  assign T513[49] = T531[49] | 1'b0;
  assign T513[48] = T531[48] | 1'b0;
  assign T513[47] = T531[47] | 1'b0;
  assign T513[46] = T531[46] | 1'b0;
  assign T513[45] = T531[45] | 1'b0;
  assign T513[44] = T531[44] | 1'b0;
  assign T513[43] = T531[43] | 1'b0;
  assign T513[42] = T531[42] | 1'b0;
  assign T513[41] = T531[41] | 1'b0;
  assign T513[40] = T531[40] | 1'b0;
  assign T513[39] = T531[39] | 1'b0;
  assign T513[38] = T531[38] | 1'b0;
  assign T513[37] = T531[37] | 1'b0;
  assign T513[36] = T531[36] | 1'b0;
  assign T513[35] = T531[35] | 1'b0;
  assign T513[34] = T531[34] | 1'b0;
  assign T513[33] = T531[33] | 1'b0;
  assign T513[32] = T531[32] | 1'b0;
  assign T513[31] = T531[31] | 1'b0;
  assign T513[30] = T531[30] | 1'b0;
  assign T513[29] = T531[29] | 1'b0;
  assign T513[28] = T531[28] | 1'b0;
  assign T513[27] = T531[27] | 1'b0;
  assign T513[26] = T531[26] | 1'b0;
  assign T513[25] = T531[25] | 1'b0;
  assign T513[24] = T531[24] | 1'b0;
  assign T513[23] = T531[23] | 1'b0;
  assign T513[22] = T531[22] | 1'b0;
  assign T513[21] = T531[21] | 1'b0;
  assign T513[20] = T531[20] | 1'b0;
  assign T513[19] = T531[19] | 1'b0;
  assign T513[18] = T531[18] | 1'b0;
  assign T513[17] = T531[17] | 1'b0;
  assign T513[16] = T531[16] | 1'b0;
  assign T513[15] = T531[15] | 1'b0;
  assign T513[14] = T531[14] | 1'b0;
  assign T513[13] = T531[13] | 1'b0;
  assign T513[12] = T531[12] | 1'b0;
  assign T513[11] = T531[11] | 1'b0;
  assign T513[10] = T531[10] | 1'b0;
  assign T513[9] = T531[9] | 1'b0;
  assign T513[8] = T531[8] | 1'b0;
  assign T513[7] = T531[7] | 1'b0;
  assign T513[6] = T531[6] | 1'b0;
  assign T513[5] = T531[5] | T950[5];
  assign T513[4] = T531[4] | 1'b0;
  assign T513[3] = T531[3] | 1'b0;
  assign T513[2] = T531[2] | 1'b0;
  assign T513[1] = T531[1] | T950_1;
  assign T513[0] = T531[0] | 1'b0;
  assign T531[63] = T580[63] | T532_63;
  assign T531[62] = T580[62] | 1'b0;
  assign T531[61] = T580[61] | 1'b0;
  assign T531[60] = T580[60] | 1'b0;
  assign T531[59] = T580[59] | 1'b0;
  assign T531[58] = T580[58] | 1'b0;
  assign T531[57] = T580[57] | 1'b0;
  assign T531[56] = T580[56] | 1'b0;
  assign T531[55] = T580[55] | 1'b0;
  assign T531[54] = T580[54] | 1'b0;
  assign T531[53] = T580[53] | 1'b0;
  assign T531[52] = T580[52] | 1'b0;
  assign T531[51] = T580[51] | 1'b0;
  assign T531[50] = T580[50] | 1'b0;
  assign T531[49] = T580[49] | 1'b0;
  assign T531[48] = T580[48] | 1'b0;
  assign T531[47] = T580[47] | 1'b0;
  assign T531[46] = T580[46] | 1'b0;
  assign T531[45] = T580[45] | 1'b0;
  assign T531[44] = T580[44] | 1'b0;
  assign T531[43] = T580[43] | 1'b0;
  assign T531[42] = T580[42] | 1'b0;
  assign T531[41] = T580[41] | 1'b0;
  assign T531[40] = T580[40] | 1'b0;
  assign T531[39] = T580[39] | 1'b0;
  assign T531[38] = T580[38] | 1'b0;
  assign T531[37] = T580[37] | 1'b0;
  assign T531[36] = T580[36] | 1'b0;
  assign T531[35] = T580[35] | 1'b0;
  assign T531[34] = T580[34] | 1'b0;
  assign T531[33] = T580[33] | 1'b0;
  assign T531[32] = T580[32] | 1'b0;
  assign T531[31] = T580[31] | T532_31;
  assign T531[30] = T580[30] | 1'b0;
  assign T531[29] = T580[29] | 1'b0;
  assign T531[28] = T580[28] | 1'b0;
  assign T531[27] = T580[27] | 1'b0;
  assign T531[26] = T580[26] | 1'b0;
  assign T531[25] = T580[25] | 1'b0;
  assign T531[24] = T580[24] | 1'b0;
  assign T531[23] = T580[23] | 1'b0;
  assign T531[22] = T580[22] | 1'b0;
  assign T531[21] = T580[21] | 1'b0;
  assign T531[20] = T580[20] | 1'b0;
  assign T531[19] = T580[19] | 1'b0;
  assign T531[18] = T580[18] | 1'b0;
  assign T531[17] = T580[17] | 1'b0;
  assign T531[16] = T580[16] | T532[16];
  assign T531[15] = T580[15] | T532[15];
  assign T531[14] = T580[14] | T532[14];
  assign T531[13] = T580[13] | T532[13];
  assign T531[12] = T580[12] | T532[12];
  assign T531[11] = T580[11] | 1'b0;
  assign T531[10] = T580[10] | 1'b0;
  assign T531[9] = T580[9] | 1'b0;
  assign T531[8] = T580[8] | 1'b0;
  assign T531[7] = T580[7] | 1'b0;
  assign T531[6] = T580[6] | 1'b0;
  assign T531[5] = T580[5] | 1'b0;
  assign T531[4] = T580[4] | T532_4;
  assign T531[3] = T580[3] | T532_3;
  assign T531[2] = T580[2] | 1'b0;
  assign T531[1] = T580[1] | 1'b0;
  assign T531[0] = T580[0] | T532_0;
  assign T580[63] = T593[63] | T581[63];
  assign T580[62] = T593[62] | T581[62];
  assign T580[61] = T593[61] | T581[61];
  assign T580[60] = T593[60] | T581[60];
  assign T580[59] = T593[59] | T581[59];
  assign T580[58] = T593[58] | T581[58];
  assign T580[57] = T593[57] | T581[57];
  assign T580[56] = T593[56] | T581[56];
  assign T580[55] = T593[55] | T581[55];
  assign T580[54] = T593[54] | T581[54];
  assign T580[53] = T593[53] | T581[53];
  assign T580[52] = T593[52] | T581[52];
  assign T580[51] = T593[51] | T581[51];
  assign T580[50] = T593[50] | T581[50];
  assign T580[49] = T593[49] | T581[49];
  assign T580[48] = T593[48] | T581[48];
  assign T580[47] = T593[47] | T581[47];
  assign T580[46] = T593[46] | T581[46];
  assign T580[45] = T593[45] | T581[45];
  assign T580[44] = T593[44] | T581[44];
  assign T580[43] = T593[43] | T581[43];
  assign T580[42] = T593[42] | T581[42];
  assign T580[41] = T593[41] | T581[41];
  assign T580[40] = T593[40] | T581[40];
  assign T580[39] = T593[39] | T581[39];
  assign T580[38] = T593[38] | T581[38];
  assign T580[37] = T593[37] | T581[37];
  assign T580[36] = T593[36] | T581[36];
  assign T580[35] = T593[35] | T581[35];
  assign T580[34] = T593[34] | T581[34];
  assign T580[33] = T593[33] | T581[33];
  assign T580[32] = T593[32] | T581[32];
  assign T580[31] = T593[31] | T581[31];
  assign T580[30] = T593[30] | T581[30];
  assign T580[29] = T593[29] | T581[29];
  assign T580[28] = T593[28] | T581[28];
  assign T580[27] = T593[27] | T581[27];
  assign T580[26] = T593[26] | T581[26];
  assign T580[25] = T593[25] | T581[25];
  assign T580[24] = T593[24] | T581[24];
  assign T580[23] = T593[23] | T581[23];
  assign T580[22] = T593[22] | T581[22];
  assign T580[21] = T593[21] | T581[21];
  assign T580[20] = T593[20] | T581[20];
  assign T580[19] = T593[19] | T581[19];
  assign T580[18] = T593[18] | T581[18];
  assign T580[17] = T593[17] | T581[17];
  assign T580[16] = T593[16] | T581[16];
  assign T580[15] = T593[15] | T581[15];
  assign T580[14] = T593[14] | T581[14];
  assign T580[13] = T593[13] | T581[13];
  assign T580[12] = T593[12] | T581[12];
  assign T580[11] = T593[11] | T581[11];
  assign T580[10] = T593[10] | T581[10];
  assign T580[9] = T593[9] | T581[9];
  assign T580[8] = T593[8] | T581[8];
  assign T580[7] = T593[7] | T581[7];
  assign T580[6] = T593[6] | T581[6];
  assign T580[5] = T593[5] | T581[5];
  assign T580[4] = T593[4] | T581[4];
  assign T580[3] = T593[3] | T581[3];
  assign T580[2] = T593[2] | T581[2];
  assign T580[1] = T593[1] | T581[1];
  assign T580[0] = T593[0] | T581[0];
  assign T591 = io_uarch_counters_15 & T586[6];
  assign T593[63] = T606[63] | T594[63];
  assign T593[62] = T606[62] | T594[62];
  assign T593[61] = T606[61] | T594[61];
  assign T593[60] = T606[60] | T594[60];
  assign T593[59] = T606[59] | T594[59];
  assign T593[58] = T606[58] | T594[58];
  assign T593[57] = T606[57] | T594[57];
  assign T593[56] = T606[56] | T594[56];
  assign T593[55] = T606[55] | T594[55];
  assign T593[54] = T606[54] | T594[54];
  assign T593[53] = T606[53] | T594[53];
  assign T593[52] = T606[52] | T594[52];
  assign T593[51] = T606[51] | T594[51];
  assign T593[50] = T606[50] | T594[50];
  assign T593[49] = T606[49] | T594[49];
  assign T593[48] = T606[48] | T594[48];
  assign T593[47] = T606[47] | T594[47];
  assign T593[46] = T606[46] | T594[46];
  assign T593[45] = T606[45] | T594[45];
  assign T593[44] = T606[44] | T594[44];
  assign T593[43] = T606[43] | T594[43];
  assign T593[42] = T606[42] | T594[42];
  assign T593[41] = T606[41] | T594[41];
  assign T593[40] = T606[40] | T594[40];
  assign T593[39] = T606[39] | T594[39];
  assign T593[38] = T606[38] | T594[38];
  assign T593[37] = T606[37] | T594[37];
  assign T593[36] = T606[36] | T594[36];
  assign T593[35] = T606[35] | T594[35];
  assign T593[34] = T606[34] | T594[34];
  assign T593[33] = T606[33] | T594[33];
  assign T593[32] = T606[32] | T594[32];
  assign T593[31] = T606[31] | T594[31];
  assign T593[30] = T606[30] | T594[30];
  assign T593[29] = T606[29] | T594[29];
  assign T593[28] = T606[28] | T594[28];
  assign T593[27] = T606[27] | T594[27];
  assign T593[26] = T606[26] | T594[26];
  assign T593[25] = T606[25] | T594[25];
  assign T593[24] = T606[24] | T594[24];
  assign T593[23] = T606[23] | T594[23];
  assign T593[22] = T606[22] | T594[22];
  assign T593[21] = T606[21] | T594[21];
  assign T593[20] = T606[20] | T594[20];
  assign T593[19] = T606[19] | T594[19];
  assign T593[18] = T606[18] | T594[18];
  assign T593[17] = T606[17] | T594[17];
  assign T593[16] = T606[16] | T594[16];
  assign T593[15] = T606[15] | T594[15];
  assign T593[14] = T606[14] | T594[14];
  assign T593[13] = T606[13] | T594[13];
  assign T593[12] = T606[12] | T594[12];
  assign T593[11] = T606[11] | T594[11];
  assign T593[10] = T606[10] | T594[10];
  assign T593[9] = T606[9] | T594[9];
  assign T593[8] = T606[8] | T594[8];
  assign T593[7] = T606[7] | T594[7];
  assign T593[6] = T606[6] | T594[6];
  assign T593[5] = T606[5] | T594[5];
  assign T593[4] = T606[4] | T594[4];
  assign T593[3] = T606[3] | T594[3];
  assign T593[2] = T606[2] | T594[2];
  assign T593[1] = T606[1] | T594[1];
  assign T593[0] = T606[0] | T594[0];
  assign T604 = io_uarch_counters_14 & T599[6];
  assign T606[63] = T619[63] | T607[63];
  assign T606[62] = T619[62] | T607[62];
  assign T606[61] = T619[61] | T607[61];
  assign T606[60] = T619[60] | T607[60];
  assign T606[59] = T619[59] | T607[59];
  assign T606[58] = T619[58] | T607[58];
  assign T606[57] = T619[57] | T607[57];
  assign T606[56] = T619[56] | T607[56];
  assign T606[55] = T619[55] | T607[55];
  assign T606[54] = T619[54] | T607[54];
  assign T606[53] = T619[53] | T607[53];
  assign T606[52] = T619[52] | T607[52];
  assign T606[51] = T619[51] | T607[51];
  assign T606[50] = T619[50] | T607[50];
  assign T606[49] = T619[49] | T607[49];
  assign T606[48] = T619[48] | T607[48];
  assign T606[47] = T619[47] | T607[47];
  assign T606[46] = T619[46] | T607[46];
  assign T606[45] = T619[45] | T607[45];
  assign T606[44] = T619[44] | T607[44];
  assign T606[43] = T619[43] | T607[43];
  assign T606[42] = T619[42] | T607[42];
  assign T606[41] = T619[41] | T607[41];
  assign T606[40] = T619[40] | T607[40];
  assign T606[39] = T619[39] | T607[39];
  assign T606[38] = T619[38] | T607[38];
  assign T606[37] = T619[37] | T607[37];
  assign T606[36] = T619[36] | T607[36];
  assign T606[35] = T619[35] | T607[35];
  assign T606[34] = T619[34] | T607[34];
  assign T606[33] = T619[33] | T607[33];
  assign T606[32] = T619[32] | T607[32];
  assign T606[31] = T619[31] | T607[31];
  assign T606[30] = T619[30] | T607[30];
  assign T606[29] = T619[29] | T607[29];
  assign T606[28] = T619[28] | T607[28];
  assign T606[27] = T619[27] | T607[27];
  assign T606[26] = T619[26] | T607[26];
  assign T606[25] = T619[25] | T607[25];
  assign T606[24] = T619[24] | T607[24];
  assign T606[23] = T619[23] | T607[23];
  assign T606[22] = T619[22] | T607[22];
  assign T606[21] = T619[21] | T607[21];
  assign T606[20] = T619[20] | T607[20];
  assign T606[19] = T619[19] | T607[19];
  assign T606[18] = T619[18] | T607[18];
  assign T606[17] = T619[17] | T607[17];
  assign T606[16] = T619[16] | T607[16];
  assign T606[15] = T619[15] | T607[15];
  assign T606[14] = T619[14] | T607[14];
  assign T606[13] = T619[13] | T607[13];
  assign T606[12] = T619[12] | T607[12];
  assign T606[11] = T619[11] | T607[11];
  assign T606[10] = T619[10] | T607[10];
  assign T606[9] = T619[9] | T607[9];
  assign T606[8] = T619[8] | T607[8];
  assign T606[7] = T619[7] | T607[7];
  assign T606[6] = T619[6] | T607[6];
  assign T606[5] = T619[5] | T607[5];
  assign T606[4] = T619[4] | T607[4];
  assign T606[3] = T619[3] | T607[3];
  assign T606[2] = T619[2] | T607[2];
  assign T606[1] = T619[1] | T607[1];
  assign T606[0] = T619[0] | T607[0];
  assign T617 = io_uarch_counters_13 & T612[6];
  assign T619[63] = T632[63] | T620[63];
  assign T619[62] = T632[62] | T620[62];
  assign T619[61] = T632[61] | T620[61];
  assign T619[60] = T632[60] | T620[60];
  assign T619[59] = T632[59] | T620[59];
  assign T619[58] = T632[58] | T620[58];
  assign T619[57] = T632[57] | T620[57];
  assign T619[56] = T632[56] | T620[56];
  assign T619[55] = T632[55] | T620[55];
  assign T619[54] = T632[54] | T620[54];
  assign T619[53] = T632[53] | T620[53];
  assign T619[52] = T632[52] | T620[52];
  assign T619[51] = T632[51] | T620[51];
  assign T619[50] = T632[50] | T620[50];
  assign T619[49] = T632[49] | T620[49];
  assign T619[48] = T632[48] | T620[48];
  assign T619[47] = T632[47] | T620[47];
  assign T619[46] = T632[46] | T620[46];
  assign T619[45] = T632[45] | T620[45];
  assign T619[44] = T632[44] | T620[44];
  assign T619[43] = T632[43] | T620[43];
  assign T619[42] = T632[42] | T620[42];
  assign T619[41] = T632[41] | T620[41];
  assign T619[40] = T632[40] | T620[40];
  assign T619[39] = T632[39] | T620[39];
  assign T619[38] = T632[38] | T620[38];
  assign T619[37] = T632[37] | T620[37];
  assign T619[36] = T632[36] | T620[36];
  assign T619[35] = T632[35] | T620[35];
  assign T619[34] = T632[34] | T620[34];
  assign T619[33] = T632[33] | T620[33];
  assign T619[32] = T632[32] | T620[32];
  assign T619[31] = T632[31] | T620[31];
  assign T619[30] = T632[30] | T620[30];
  assign T619[29] = T632[29] | T620[29];
  assign T619[28] = T632[28] | T620[28];
  assign T619[27] = T632[27] | T620[27];
  assign T619[26] = T632[26] | T620[26];
  assign T619[25] = T632[25] | T620[25];
  assign T619[24] = T632[24] | T620[24];
  assign T619[23] = T632[23] | T620[23];
  assign T619[22] = T632[22] | T620[22];
  assign T619[21] = T632[21] | T620[21];
  assign T619[20] = T632[20] | T620[20];
  assign T619[19] = T632[19] | T620[19];
  assign T619[18] = T632[18] | T620[18];
  assign T619[17] = T632[17] | T620[17];
  assign T619[16] = T632[16] | T620[16];
  assign T619[15] = T632[15] | T620[15];
  assign T619[14] = T632[14] | T620[14];
  assign T619[13] = T632[13] | T620[13];
  assign T619[12] = T632[12] | T620[12];
  assign T619[11] = T632[11] | T620[11];
  assign T619[10] = T632[10] | T620[10];
  assign T619[9] = T632[9] | T620[9];
  assign T619[8] = T632[8] | T620[8];
  assign T619[7] = T632[7] | T620[7];
  assign T619[6] = T632[6] | T620[6];
  assign T619[5] = T632[5] | T620[5];
  assign T619[4] = T632[4] | T620[4];
  assign T619[3] = T632[3] | T620[3];
  assign T619[2] = T632[2] | T620[2];
  assign T619[1] = T632[1] | T620[1];
  assign T619[0] = T632[0] | T620[0];
  assign T630 = io_uarch_counters_12 & T625[6];
  assign T632[63] = T645[63] | T633[63];
  assign T632[62] = T645[62] | T633[62];
  assign T632[61] = T645[61] | T633[61];
  assign T632[60] = T645[60] | T633[60];
  assign T632[59] = T645[59] | T633[59];
  assign T632[58] = T645[58] | T633[58];
  assign T632[57] = T645[57] | T633[57];
  assign T632[56] = T645[56] | T633[56];
  assign T632[55] = T645[55] | T633[55];
  assign T632[54] = T645[54] | T633[54];
  assign T632[53] = T645[53] | T633[53];
  assign T632[52] = T645[52] | T633[52];
  assign T632[51] = T645[51] | T633[51];
  assign T632[50] = T645[50] | T633[50];
  assign T632[49] = T645[49] | T633[49];
  assign T632[48] = T645[48] | T633[48];
  assign T632[47] = T645[47] | T633[47];
  assign T632[46] = T645[46] | T633[46];
  assign T632[45] = T645[45] | T633[45];
  assign T632[44] = T645[44] | T633[44];
  assign T632[43] = T645[43] | T633[43];
  assign T632[42] = T645[42] | T633[42];
  assign T632[41] = T645[41] | T633[41];
  assign T632[40] = T645[40] | T633[40];
  assign T632[39] = T645[39] | T633[39];
  assign T632[38] = T645[38] | T633[38];
  assign T632[37] = T645[37] | T633[37];
  assign T632[36] = T645[36] | T633[36];
  assign T632[35] = T645[35] | T633[35];
  assign T632[34] = T645[34] | T633[34];
  assign T632[33] = T645[33] | T633[33];
  assign T632[32] = T645[32] | T633[32];
  assign T632[31] = T645[31] | T633[31];
  assign T632[30] = T645[30] | T633[30];
  assign T632[29] = T645[29] | T633[29];
  assign T632[28] = T645[28] | T633[28];
  assign T632[27] = T645[27] | T633[27];
  assign T632[26] = T645[26] | T633[26];
  assign T632[25] = T645[25] | T633[25];
  assign T632[24] = T645[24] | T633[24];
  assign T632[23] = T645[23] | T633[23];
  assign T632[22] = T645[22] | T633[22];
  assign T632[21] = T645[21] | T633[21];
  assign T632[20] = T645[20] | T633[20];
  assign T632[19] = T645[19] | T633[19];
  assign T632[18] = T645[18] | T633[18];
  assign T632[17] = T645[17] | T633[17];
  assign T632[16] = T645[16] | T633[16];
  assign T632[15] = T645[15] | T633[15];
  assign T632[14] = T645[14] | T633[14];
  assign T632[13] = T645[13] | T633[13];
  assign T632[12] = T645[12] | T633[12];
  assign T632[11] = T645[11] | T633[11];
  assign T632[10] = T645[10] | T633[10];
  assign T632[9] = T645[9] | T633[9];
  assign T632[8] = T645[8] | T633[8];
  assign T632[7] = T645[7] | T633[7];
  assign T632[6] = T645[6] | T633[6];
  assign T632[5] = T645[5] | T633[5];
  assign T632[4] = T645[4] | T633[4];
  assign T632[3] = T645[3] | T633[3];
  assign T632[2] = T645[2] | T633[2];
  assign T632[1] = T645[1] | T633[1];
  assign T632[0] = T645[0] | T633[0];
  assign T643 = io_uarch_counters_11 & T638[6];
  assign T645[63] = T658[63] | T646[63];
  assign T645[62] = T658[62] | T646[62];
  assign T645[61] = T658[61] | T646[61];
  assign T645[60] = T658[60] | T646[60];
  assign T645[59] = T658[59] | T646[59];
  assign T645[58] = T658[58] | T646[58];
  assign T645[57] = T658[57] | T646[57];
  assign T645[56] = T658[56] | T646[56];
  assign T645[55] = T658[55] | T646[55];
  assign T645[54] = T658[54] | T646[54];
  assign T645[53] = T658[53] | T646[53];
  assign T645[52] = T658[52] | T646[52];
  assign T645[51] = T658[51] | T646[51];
  assign T645[50] = T658[50] | T646[50];
  assign T645[49] = T658[49] | T646[49];
  assign T645[48] = T658[48] | T646[48];
  assign T645[47] = T658[47] | T646[47];
  assign T645[46] = T658[46] | T646[46];
  assign T645[45] = T658[45] | T646[45];
  assign T645[44] = T658[44] | T646[44];
  assign T645[43] = T658[43] | T646[43];
  assign T645[42] = T658[42] | T646[42];
  assign T645[41] = T658[41] | T646[41];
  assign T645[40] = T658[40] | T646[40];
  assign T645[39] = T658[39] | T646[39];
  assign T645[38] = T658[38] | T646[38];
  assign T645[37] = T658[37] | T646[37];
  assign T645[36] = T658[36] | T646[36];
  assign T645[35] = T658[35] | T646[35];
  assign T645[34] = T658[34] | T646[34];
  assign T645[33] = T658[33] | T646[33];
  assign T645[32] = T658[32] | T646[32];
  assign T645[31] = T658[31] | T646[31];
  assign T645[30] = T658[30] | T646[30];
  assign T645[29] = T658[29] | T646[29];
  assign T645[28] = T658[28] | T646[28];
  assign T645[27] = T658[27] | T646[27];
  assign T645[26] = T658[26] | T646[26];
  assign T645[25] = T658[25] | T646[25];
  assign T645[24] = T658[24] | T646[24];
  assign T645[23] = T658[23] | T646[23];
  assign T645[22] = T658[22] | T646[22];
  assign T645[21] = T658[21] | T646[21];
  assign T645[20] = T658[20] | T646[20];
  assign T645[19] = T658[19] | T646[19];
  assign T645[18] = T658[18] | T646[18];
  assign T645[17] = T658[17] | T646[17];
  assign T645[16] = T658[16] | T646[16];
  assign T645[15] = T658[15] | T646[15];
  assign T645[14] = T658[14] | T646[14];
  assign T645[13] = T658[13] | T646[13];
  assign T645[12] = T658[12] | T646[12];
  assign T645[11] = T658[11] | T646[11];
  assign T645[10] = T658[10] | T646[10];
  assign T645[9] = T658[9] | T646[9];
  assign T645[8] = T658[8] | T646[8];
  assign T645[7] = T658[7] | T646[7];
  assign T645[6] = T658[6] | T646[6];
  assign T645[5] = T658[5] | T646[5];
  assign T645[4] = T658[4] | T646[4];
  assign T645[3] = T658[3] | T646[3];
  assign T645[2] = T658[2] | T646[2];
  assign T645[1] = T658[1] | T646[1];
  assign T645[0] = T658[0] | T646[0];
  assign T656 = io_uarch_counters_10 & T651[6];
  assign T658[63] = T671[63] | T659[63];
  assign T658[62] = T671[62] | T659[62];
  assign T658[61] = T671[61] | T659[61];
  assign T658[60] = T671[60] | T659[60];
  assign T658[59] = T671[59] | T659[59];
  assign T658[58] = T671[58] | T659[58];
  assign T658[57] = T671[57] | T659[57];
  assign T658[56] = T671[56] | T659[56];
  assign T658[55] = T671[55] | T659[55];
  assign T658[54] = T671[54] | T659[54];
  assign T658[53] = T671[53] | T659[53];
  assign T658[52] = T671[52] | T659[52];
  assign T658[51] = T671[51] | T659[51];
  assign T658[50] = T671[50] | T659[50];
  assign T658[49] = T671[49] | T659[49];
  assign T658[48] = T671[48] | T659[48];
  assign T658[47] = T671[47] | T659[47];
  assign T658[46] = T671[46] | T659[46];
  assign T658[45] = T671[45] | T659[45];
  assign T658[44] = T671[44] | T659[44];
  assign T658[43] = T671[43] | T659[43];
  assign T658[42] = T671[42] | T659[42];
  assign T658[41] = T671[41] | T659[41];
  assign T658[40] = T671[40] | T659[40];
  assign T658[39] = T671[39] | T659[39];
  assign T658[38] = T671[38] | T659[38];
  assign T658[37] = T671[37] | T659[37];
  assign T658[36] = T671[36] | T659[36];
  assign T658[35] = T671[35] | T659[35];
  assign T658[34] = T671[34] | T659[34];
  assign T658[33] = T671[33] | T659[33];
  assign T658[32] = T671[32] | T659[32];
  assign T658[31] = T671[31] | T659[31];
  assign T658[30] = T671[30] | T659[30];
  assign T658[29] = T671[29] | T659[29];
  assign T658[28] = T671[28] | T659[28];
  assign T658[27] = T671[27] | T659[27];
  assign T658[26] = T671[26] | T659[26];
  assign T658[25] = T671[25] | T659[25];
  assign T658[24] = T671[24] | T659[24];
  assign T658[23] = T671[23] | T659[23];
  assign T658[22] = T671[22] | T659[22];
  assign T658[21] = T671[21] | T659[21];
  assign T658[20] = T671[20] | T659[20];
  assign T658[19] = T671[19] | T659[19];
  assign T658[18] = T671[18] | T659[18];
  assign T658[17] = T671[17] | T659[17];
  assign T658[16] = T671[16] | T659[16];
  assign T658[15] = T671[15] | T659[15];
  assign T658[14] = T671[14] | T659[14];
  assign T658[13] = T671[13] | T659[13];
  assign T658[12] = T671[12] | T659[12];
  assign T658[11] = T671[11] | T659[11];
  assign T658[10] = T671[10] | T659[10];
  assign T658[9] = T671[9] | T659[9];
  assign T658[8] = T671[8] | T659[8];
  assign T658[7] = T671[7] | T659[7];
  assign T658[6] = T671[6] | T659[6];
  assign T658[5] = T671[5] | T659[5];
  assign T658[4] = T671[4] | T659[4];
  assign T658[3] = T671[3] | T659[3];
  assign T658[2] = T671[2] | T659[2];
  assign T658[1] = T671[1] | T659[1];
  assign T658[0] = T671[0] | T659[0];
  assign T669 = io_uarch_counters_9 & T664[6];
  assign T671[63] = T684[63] | T672[63];
  assign T671[62] = T684[62] | T672[62];
  assign T671[61] = T684[61] | T672[61];
  assign T671[60] = T684[60] | T672[60];
  assign T671[59] = T684[59] | T672[59];
  assign T671[58] = T684[58] | T672[58];
  assign T671[57] = T684[57] | T672[57];
  assign T671[56] = T684[56] | T672[56];
  assign T671[55] = T684[55] | T672[55];
  assign T671[54] = T684[54] | T672[54];
  assign T671[53] = T684[53] | T672[53];
  assign T671[52] = T684[52] | T672[52];
  assign T671[51] = T684[51] | T672[51];
  assign T671[50] = T684[50] | T672[50];
  assign T671[49] = T684[49] | T672[49];
  assign T671[48] = T684[48] | T672[48];
  assign T671[47] = T684[47] | T672[47];
  assign T671[46] = T684[46] | T672[46];
  assign T671[45] = T684[45] | T672[45];
  assign T671[44] = T684[44] | T672[44];
  assign T671[43] = T684[43] | T672[43];
  assign T671[42] = T684[42] | T672[42];
  assign T671[41] = T684[41] | T672[41];
  assign T671[40] = T684[40] | T672[40];
  assign T671[39] = T684[39] | T672[39];
  assign T671[38] = T684[38] | T672[38];
  assign T671[37] = T684[37] | T672[37];
  assign T671[36] = T684[36] | T672[36];
  assign T671[35] = T684[35] | T672[35];
  assign T671[34] = T684[34] | T672[34];
  assign T671[33] = T684[33] | T672[33];
  assign T671[32] = T684[32] | T672[32];
  assign T671[31] = T684[31] | T672[31];
  assign T671[30] = T684[30] | T672[30];
  assign T671[29] = T684[29] | T672[29];
  assign T671[28] = T684[28] | T672[28];
  assign T671[27] = T684[27] | T672[27];
  assign T671[26] = T684[26] | T672[26];
  assign T671[25] = T684[25] | T672[25];
  assign T671[24] = T684[24] | T672[24];
  assign T671[23] = T684[23] | T672[23];
  assign T671[22] = T684[22] | T672[22];
  assign T671[21] = T684[21] | T672[21];
  assign T671[20] = T684[20] | T672[20];
  assign T671[19] = T684[19] | T672[19];
  assign T671[18] = T684[18] | T672[18];
  assign T671[17] = T684[17] | T672[17];
  assign T671[16] = T684[16] | T672[16];
  assign T671[15] = T684[15] | T672[15];
  assign T671[14] = T684[14] | T672[14];
  assign T671[13] = T684[13] | T672[13];
  assign T671[12] = T684[12] | T672[12];
  assign T671[11] = T684[11] | T672[11];
  assign T671[10] = T684[10] | T672[10];
  assign T671[9] = T684[9] | T672[9];
  assign T671[8] = T684[8] | T672[8];
  assign T671[7] = T684[7] | T672[7];
  assign T671[6] = T684[6] | T672[6];
  assign T671[5] = T684[5] | T672[5];
  assign T671[4] = T684[4] | T672[4];
  assign T671[3] = T684[3] | T672[3];
  assign T671[2] = T684[2] | T672[2];
  assign T671[1] = T684[1] | T672[1];
  assign T671[0] = T684[0] | T672[0];
  assign T682 = io_uarch_counters_8 & T677[6];
  assign T684[63] = T697[63] | T685[63];
  assign T684[62] = T697[62] | T685[62];
  assign T684[61] = T697[61] | T685[61];
  assign T684[60] = T697[60] | T685[60];
  assign T684[59] = T697[59] | T685[59];
  assign T684[58] = T697[58] | T685[58];
  assign T684[57] = T697[57] | T685[57];
  assign T684[56] = T697[56] | T685[56];
  assign T684[55] = T697[55] | T685[55];
  assign T684[54] = T697[54] | T685[54];
  assign T684[53] = T697[53] | T685[53];
  assign T684[52] = T697[52] | T685[52];
  assign T684[51] = T697[51] | T685[51];
  assign T684[50] = T697[50] | T685[50];
  assign T684[49] = T697[49] | T685[49];
  assign T684[48] = T697[48] | T685[48];
  assign T684[47] = T697[47] | T685[47];
  assign T684[46] = T697[46] | T685[46];
  assign T684[45] = T697[45] | T685[45];
  assign T684[44] = T697[44] | T685[44];
  assign T684[43] = T697[43] | T685[43];
  assign T684[42] = T697[42] | T685[42];
  assign T684[41] = T697[41] | T685[41];
  assign T684[40] = T697[40] | T685[40];
  assign T684[39] = T697[39] | T685[39];
  assign T684[38] = T697[38] | T685[38];
  assign T684[37] = T697[37] | T685[37];
  assign T684[36] = T697[36] | T685[36];
  assign T684[35] = T697[35] | T685[35];
  assign T684[34] = T697[34] | T685[34];
  assign T684[33] = T697[33] | T685[33];
  assign T684[32] = T697[32] | T685[32];
  assign T684[31] = T697[31] | T685[31];
  assign T684[30] = T697[30] | T685[30];
  assign T684[29] = T697[29] | T685[29];
  assign T684[28] = T697[28] | T685[28];
  assign T684[27] = T697[27] | T685[27];
  assign T684[26] = T697[26] | T685[26];
  assign T684[25] = T697[25] | T685[25];
  assign T684[24] = T697[24] | T685[24];
  assign T684[23] = T697[23] | T685[23];
  assign T684[22] = T697[22] | T685[22];
  assign T684[21] = T697[21] | T685[21];
  assign T684[20] = T697[20] | T685[20];
  assign T684[19] = T697[19] | T685[19];
  assign T684[18] = T697[18] | T685[18];
  assign T684[17] = T697[17] | T685[17];
  assign T684[16] = T697[16] | T685[16];
  assign T684[15] = T697[15] | T685[15];
  assign T684[14] = T697[14] | T685[14];
  assign T684[13] = T697[13] | T685[13];
  assign T684[12] = T697[12] | T685[12];
  assign T684[11] = T697[11] | T685[11];
  assign T684[10] = T697[10] | T685[10];
  assign T684[9] = T697[9] | T685[9];
  assign T684[8] = T697[8] | T685[8];
  assign T684[7] = T697[7] | T685[7];
  assign T684[6] = T697[6] | T685[6];
  assign T684[5] = T697[5] | T685[5];
  assign T684[4] = T697[4] | T685[4];
  assign T684[3] = T697[3] | T685[3];
  assign T684[2] = T697[2] | T685[2];
  assign T684[1] = T697[1] | T685[1];
  assign T684[0] = T697[0] | T685[0];
  assign T695 = io_uarch_counters_7 & T690[6];
  assign T697[63] = T710[63] | T698[63];
  assign T697[62] = T710[62] | T698[62];
  assign T697[61] = T710[61] | T698[61];
  assign T697[60] = T710[60] | T698[60];
  assign T697[59] = T710[59] | T698[59];
  assign T697[58] = T710[58] | T698[58];
  assign T697[57] = T710[57] | T698[57];
  assign T697[56] = T710[56] | T698[56];
  assign T697[55] = T710[55] | T698[55];
  assign T697[54] = T710[54] | T698[54];
  assign T697[53] = T710[53] | T698[53];
  assign T697[52] = T710[52] | T698[52];
  assign T697[51] = T710[51] | T698[51];
  assign T697[50] = T710[50] | T698[50];
  assign T697[49] = T710[49] | T698[49];
  assign T697[48] = T710[48] | T698[48];
  assign T697[47] = T710[47] | T698[47];
  assign T697[46] = T710[46] | T698[46];
  assign T697[45] = T710[45] | T698[45];
  assign T697[44] = T710[44] | T698[44];
  assign T697[43] = T710[43] | T698[43];
  assign T697[42] = T710[42] | T698[42];
  assign T697[41] = T710[41] | T698[41];
  assign T697[40] = T710[40] | T698[40];
  assign T697[39] = T710[39] | T698[39];
  assign T697[38] = T710[38] | T698[38];
  assign T697[37] = T710[37] | T698[37];
  assign T697[36] = T710[36] | T698[36];
  assign T697[35] = T710[35] | T698[35];
  assign T697[34] = T710[34] | T698[34];
  assign T697[33] = T710[33] | T698[33];
  assign T697[32] = T710[32] | T698[32];
  assign T697[31] = T710[31] | T698[31];
  assign T697[30] = T710[30] | T698[30];
  assign T697[29] = T710[29] | T698[29];
  assign T697[28] = T710[28] | T698[28];
  assign T697[27] = T710[27] | T698[27];
  assign T697[26] = T710[26] | T698[26];
  assign T697[25] = T710[25] | T698[25];
  assign T697[24] = T710[24] | T698[24];
  assign T697[23] = T710[23] | T698[23];
  assign T697[22] = T710[22] | T698[22];
  assign T697[21] = T710[21] | T698[21];
  assign T697[20] = T710[20] | T698[20];
  assign T697[19] = T710[19] | T698[19];
  assign T697[18] = T710[18] | T698[18];
  assign T697[17] = T710[17] | T698[17];
  assign T697[16] = T710[16] | T698[16];
  assign T697[15] = T710[15] | T698[15];
  assign T697[14] = T710[14] | T698[14];
  assign T697[13] = T710[13] | T698[13];
  assign T697[12] = T710[12] | T698[12];
  assign T697[11] = T710[11] | T698[11];
  assign T697[10] = T710[10] | T698[10];
  assign T697[9] = T710[9] | T698[9];
  assign T697[8] = T710[8] | T698[8];
  assign T697[7] = T710[7] | T698[7];
  assign T697[6] = T710[6] | T698[6];
  assign T697[5] = T710[5] | T698[5];
  assign T697[4] = T710[4] | T698[4];
  assign T697[3] = T710[3] | T698[3];
  assign T697[2] = T710[2] | T698[2];
  assign T697[1] = T710[1] | T698[1];
  assign T697[0] = T710[0] | T698[0];
  assign T708 = io_uarch_counters_6 & T703[6];
  assign T710[63] = T723[63] | T711[63];
  assign T710[62] = T723[62] | T711[62];
  assign T710[61] = T723[61] | T711[61];
  assign T710[60] = T723[60] | T711[60];
  assign T710[59] = T723[59] | T711[59];
  assign T710[58] = T723[58] | T711[58];
  assign T710[57] = T723[57] | T711[57];
  assign T710[56] = T723[56] | T711[56];
  assign T710[55] = T723[55] | T711[55];
  assign T710[54] = T723[54] | T711[54];
  assign T710[53] = T723[53] | T711[53];
  assign T710[52] = T723[52] | T711[52];
  assign T710[51] = T723[51] | T711[51];
  assign T710[50] = T723[50] | T711[50];
  assign T710[49] = T723[49] | T711[49];
  assign T710[48] = T723[48] | T711[48];
  assign T710[47] = T723[47] | T711[47];
  assign T710[46] = T723[46] | T711[46];
  assign T710[45] = T723[45] | T711[45];
  assign T710[44] = T723[44] | T711[44];
  assign T710[43] = T723[43] | T711[43];
  assign T710[42] = T723[42] | T711[42];
  assign T710[41] = T723[41] | T711[41];
  assign T710[40] = T723[40] | T711[40];
  assign T710[39] = T723[39] | T711[39];
  assign T710[38] = T723[38] | T711[38];
  assign T710[37] = T723[37] | T711[37];
  assign T710[36] = T723[36] | T711[36];
  assign T710[35] = T723[35] | T711[35];
  assign T710[34] = T723[34] | T711[34];
  assign T710[33] = T723[33] | T711[33];
  assign T710[32] = T723[32] | T711[32];
  assign T710[31] = T723[31] | T711[31];
  assign T710[30] = T723[30] | T711[30];
  assign T710[29] = T723[29] | T711[29];
  assign T710[28] = T723[28] | T711[28];
  assign T710[27] = T723[27] | T711[27];
  assign T710[26] = T723[26] | T711[26];
  assign T710[25] = T723[25] | T711[25];
  assign T710[24] = T723[24] | T711[24];
  assign T710[23] = T723[23] | T711[23];
  assign T710[22] = T723[22] | T711[22];
  assign T710[21] = T723[21] | T711[21];
  assign T710[20] = T723[20] | T711[20];
  assign T710[19] = T723[19] | T711[19];
  assign T710[18] = T723[18] | T711[18];
  assign T710[17] = T723[17] | T711[17];
  assign T710[16] = T723[16] | T711[16];
  assign T710[15] = T723[15] | T711[15];
  assign T710[14] = T723[14] | T711[14];
  assign T710[13] = T723[13] | T711[13];
  assign T710[12] = T723[12] | T711[12];
  assign T710[11] = T723[11] | T711[11];
  assign T710[10] = T723[10] | T711[10];
  assign T710[9] = T723[9] | T711[9];
  assign T710[8] = T723[8] | T711[8];
  assign T710[7] = T723[7] | T711[7];
  assign T710[6] = T723[6] | T711[6];
  assign T710[5] = T723[5] | T711[5];
  assign T710[4] = T723[4] | T711[4];
  assign T710[3] = T723[3] | T711[3];
  assign T710[2] = T723[2] | T711[2];
  assign T710[1] = T723[1] | T711[1];
  assign T710[0] = T723[0] | T711[0];
  assign T721 = io_uarch_counters_5 & T716[6];
  assign T723[63] = T736[63] | T724[63];
  assign T723[62] = T736[62] | T724[62];
  assign T723[61] = T736[61] | T724[61];
  assign T723[60] = T736[60] | T724[60];
  assign T723[59] = T736[59] | T724[59];
  assign T723[58] = T736[58] | T724[58];
  assign T723[57] = T736[57] | T724[57];
  assign T723[56] = T736[56] | T724[56];
  assign T723[55] = T736[55] | T724[55];
  assign T723[54] = T736[54] | T724[54];
  assign T723[53] = T736[53] | T724[53];
  assign T723[52] = T736[52] | T724[52];
  assign T723[51] = T736[51] | T724[51];
  assign T723[50] = T736[50] | T724[50];
  assign T723[49] = T736[49] | T724[49];
  assign T723[48] = T736[48] | T724[48];
  assign T723[47] = T736[47] | T724[47];
  assign T723[46] = T736[46] | T724[46];
  assign T723[45] = T736[45] | T724[45];
  assign T723[44] = T736[44] | T724[44];
  assign T723[43] = T736[43] | T724[43];
  assign T723[42] = T736[42] | T724[42];
  assign T723[41] = T736[41] | T724[41];
  assign T723[40] = T736[40] | T724[40];
  assign T723[39] = T736[39] | T724[39];
  assign T723[38] = T736[38] | T724[38];
  assign T723[37] = T736[37] | T724[37];
  assign T723[36] = T736[36] | T724[36];
  assign T723[35] = T736[35] | T724[35];
  assign T723[34] = T736[34] | T724[34];
  assign T723[33] = T736[33] | T724[33];
  assign T723[32] = T736[32] | T724[32];
  assign T723[31] = T736[31] | T724[31];
  assign T723[30] = T736[30] | T724[30];
  assign T723[29] = T736[29] | T724[29];
  assign T723[28] = T736[28] | T724[28];
  assign T723[27] = T736[27] | T724[27];
  assign T723[26] = T736[26] | T724[26];
  assign T723[25] = T736[25] | T724[25];
  assign T723[24] = T736[24] | T724[24];
  assign T723[23] = T736[23] | T724[23];
  assign T723[22] = T736[22] | T724[22];
  assign T723[21] = T736[21] | T724[21];
  assign T723[20] = T736[20] | T724[20];
  assign T723[19] = T736[19] | T724[19];
  assign T723[18] = T736[18] | T724[18];
  assign T723[17] = T736[17] | T724[17];
  assign T723[16] = T736[16] | T724[16];
  assign T723[15] = T736[15] | T724[15];
  assign T723[14] = T736[14] | T724[14];
  assign T723[13] = T736[13] | T724[13];
  assign T723[12] = T736[12] | T724[12];
  assign T723[11] = T736[11] | T724[11];
  assign T723[10] = T736[10] | T724[10];
  assign T723[9] = T736[9] | T724[9];
  assign T723[8] = T736[8] | T724[8];
  assign T723[7] = T736[7] | T724[7];
  assign T723[6] = T736[6] | T724[6];
  assign T723[5] = T736[5] | T724[5];
  assign T723[4] = T736[4] | T724[4];
  assign T723[3] = T736[3] | T724[3];
  assign T723[2] = T736[2] | T724[2];
  assign T723[1] = T736[1] | T724[1];
  assign T723[0] = T736[0] | T724[0];
  assign T734 = io_uarch_counters_4 & T729[6];
  assign T736[63] = T749[63] | T737[63];
  assign T736[62] = T749[62] | T737[62];
  assign T736[61] = T749[61] | T737[61];
  assign T736[60] = T749[60] | T737[60];
  assign T736[59] = T749[59] | T737[59];
  assign T736[58] = T749[58] | T737[58];
  assign T736[57] = T749[57] | T737[57];
  assign T736[56] = T749[56] | T737[56];
  assign T736[55] = T749[55] | T737[55];
  assign T736[54] = T749[54] | T737[54];
  assign T736[53] = T749[53] | T737[53];
  assign T736[52] = T749[52] | T737[52];
  assign T736[51] = T749[51] | T737[51];
  assign T736[50] = T749[50] | T737[50];
  assign T736[49] = T749[49] | T737[49];
  assign T736[48] = T749[48] | T737[48];
  assign T736[47] = T749[47] | T737[47];
  assign T736[46] = T749[46] | T737[46];
  assign T736[45] = T749[45] | T737[45];
  assign T736[44] = T749[44] | T737[44];
  assign T736[43] = T749[43] | T737[43];
  assign T736[42] = T749[42] | T737[42];
  assign T736[41] = T749[41] | T737[41];
  assign T736[40] = T749[40] | T737[40];
  assign T736[39] = T749[39] | T737[39];
  assign T736[38] = T749[38] | T737[38];
  assign T736[37] = T749[37] | T737[37];
  assign T736[36] = T749[36] | T737[36];
  assign T736[35] = T749[35] | T737[35];
  assign T736[34] = T749[34] | T737[34];
  assign T736[33] = T749[33] | T737[33];
  assign T736[32] = T749[32] | T737[32];
  assign T736[31] = T749[31] | T737[31];
  assign T736[30] = T749[30] | T737[30];
  assign T736[29] = T749[29] | T737[29];
  assign T736[28] = T749[28] | T737[28];
  assign T736[27] = T749[27] | T737[27];
  assign T736[26] = T749[26] | T737[26];
  assign T736[25] = T749[25] | T737[25];
  assign T736[24] = T749[24] | T737[24];
  assign T736[23] = T749[23] | T737[23];
  assign T736[22] = T749[22] | T737[22];
  assign T736[21] = T749[21] | T737[21];
  assign T736[20] = T749[20] | T737[20];
  assign T736[19] = T749[19] | T737[19];
  assign T736[18] = T749[18] | T737[18];
  assign T736[17] = T749[17] | T737[17];
  assign T736[16] = T749[16] | T737[16];
  assign T736[15] = T749[15] | T737[15];
  assign T736[14] = T749[14] | T737[14];
  assign T736[13] = T749[13] | T737[13];
  assign T736[12] = T749[12] | T737[12];
  assign T736[11] = T749[11] | T737[11];
  assign T736[10] = T749[10] | T737[10];
  assign T736[9] = T749[9] | T737[9];
  assign T736[8] = T749[8] | T737[8];
  assign T736[7] = T749[7] | T737[7];
  assign T736[6] = T749[6] | T737[6];
  assign T736[5] = T749[5] | T737[5];
  assign T736[4] = T749[4] | T737[4];
  assign T736[3] = T749[3] | T737[3];
  assign T736[2] = T749[2] | T737[2];
  assign T736[1] = T749[1] | T737[1];
  assign T736[0] = T749[0] | T737[0];
  assign T747 = io_uarch_counters_3 & T742[6];
  assign T749[63] = T762[63] | T750[63];
  assign T749[62] = T762[62] | T750[62];
  assign T749[61] = T762[61] | T750[61];
  assign T749[60] = T762[60] | T750[60];
  assign T749[59] = T762[59] | T750[59];
  assign T749[58] = T762[58] | T750[58];
  assign T749[57] = T762[57] | T750[57];
  assign T749[56] = T762[56] | T750[56];
  assign T749[55] = T762[55] | T750[55];
  assign T749[54] = T762[54] | T750[54];
  assign T749[53] = T762[53] | T750[53];
  assign T749[52] = T762[52] | T750[52];
  assign T749[51] = T762[51] | T750[51];
  assign T749[50] = T762[50] | T750[50];
  assign T749[49] = T762[49] | T750[49];
  assign T749[48] = T762[48] | T750[48];
  assign T749[47] = T762[47] | T750[47];
  assign T749[46] = T762[46] | T750[46];
  assign T749[45] = T762[45] | T750[45];
  assign T749[44] = T762[44] | T750[44];
  assign T749[43] = T762[43] | T750[43];
  assign T749[42] = T762[42] | T750[42];
  assign T749[41] = T762[41] | T750[41];
  assign T749[40] = T762[40] | T750[40];
  assign T749[39] = T762[39] | T750[39];
  assign T749[38] = T762[38] | T750[38];
  assign T749[37] = T762[37] | T750[37];
  assign T749[36] = T762[36] | T750[36];
  assign T749[35] = T762[35] | T750[35];
  assign T749[34] = T762[34] | T750[34];
  assign T749[33] = T762[33] | T750[33];
  assign T749[32] = T762[32] | T750[32];
  assign T749[31] = T762[31] | T750[31];
  assign T749[30] = T762[30] | T750[30];
  assign T749[29] = T762[29] | T750[29];
  assign T749[28] = T762[28] | T750[28];
  assign T749[27] = T762[27] | T750[27];
  assign T749[26] = T762[26] | T750[26];
  assign T749[25] = T762[25] | T750[25];
  assign T749[24] = T762[24] | T750[24];
  assign T749[23] = T762[23] | T750[23];
  assign T749[22] = T762[22] | T750[22];
  assign T749[21] = T762[21] | T750[21];
  assign T749[20] = T762[20] | T750[20];
  assign T749[19] = T762[19] | T750[19];
  assign T749[18] = T762[18] | T750[18];
  assign T749[17] = T762[17] | T750[17];
  assign T749[16] = T762[16] | T750[16];
  assign T749[15] = T762[15] | T750[15];
  assign T749[14] = T762[14] | T750[14];
  assign T749[13] = T762[13] | T750[13];
  assign T749[12] = T762[12] | T750[12];
  assign T749[11] = T762[11] | T750[11];
  assign T749[10] = T762[10] | T750[10];
  assign T749[9] = T762[9] | T750[9];
  assign T749[8] = T762[8] | T750[8];
  assign T749[7] = T762[7] | T750[7];
  assign T749[6] = T762[6] | T750[6];
  assign T749[5] = T762[5] | T750[5];
  assign T749[4] = T762[4] | T750[4];
  assign T749[3] = T762[3] | T750[3];
  assign T749[2] = T762[2] | T750[2];
  assign T749[1] = T762[1] | T750[1];
  assign T749[0] = T762[0] | T750[0];
  assign T760 = io_uarch_counters_2 & T755[6];
  assign T762[63] = T775[63] | T763[63];
  assign T762[62] = T775[62] | T763[62];
  assign T762[61] = T775[61] | T763[61];
  assign T762[60] = T775[60] | T763[60];
  assign T762[59] = T775[59] | T763[59];
  assign T762[58] = T775[58] | T763[58];
  assign T762[57] = T775[57] | T763[57];
  assign T762[56] = T775[56] | T763[56];
  assign T762[55] = T775[55] | T763[55];
  assign T762[54] = T775[54] | T763[54];
  assign T762[53] = T775[53] | T763[53];
  assign T762[52] = T775[52] | T763[52];
  assign T762[51] = T775[51] | T763[51];
  assign T762[50] = T775[50] | T763[50];
  assign T762[49] = T775[49] | T763[49];
  assign T762[48] = T775[48] | T763[48];
  assign T762[47] = T775[47] | T763[47];
  assign T762[46] = T775[46] | T763[46];
  assign T762[45] = T775[45] | T763[45];
  assign T762[44] = T775[44] | T763[44];
  assign T762[43] = T775[43] | T763[43];
  assign T762[42] = T775[42] | T763[42];
  assign T762[41] = T775[41] | T763[41];
  assign T762[40] = T775[40] | T763[40];
  assign T762[39] = T775[39] | T763[39];
  assign T762[38] = T775[38] | T763[38];
  assign T762[37] = T775[37] | T763[37];
  assign T762[36] = T775[36] | T763[36];
  assign T762[35] = T775[35] | T763[35];
  assign T762[34] = T775[34] | T763[34];
  assign T762[33] = T775[33] | T763[33];
  assign T762[32] = T775[32] | T763[32];
  assign T762[31] = T775[31] | T763[31];
  assign T762[30] = T775[30] | T763[30];
  assign T762[29] = T775[29] | T763[29];
  assign T762[28] = T775[28] | T763[28];
  assign T762[27] = T775[27] | T763[27];
  assign T762[26] = T775[26] | T763[26];
  assign T762[25] = T775[25] | T763[25];
  assign T762[24] = T775[24] | T763[24];
  assign T762[23] = T775[23] | T763[23];
  assign T762[22] = T775[22] | T763[22];
  assign T762[21] = T775[21] | T763[21];
  assign T762[20] = T775[20] | T763[20];
  assign T762[19] = T775[19] | T763[19];
  assign T762[18] = T775[18] | T763[18];
  assign T762[17] = T775[17] | T763[17];
  assign T762[16] = T775[16] | T763[16];
  assign T762[15] = T775[15] | T763[15];
  assign T762[14] = T775[14] | T763[14];
  assign T762[13] = T775[13] | T763[13];
  assign T762[12] = T775[12] | T763[12];
  assign T762[11] = T775[11] | T763[11];
  assign T762[10] = T775[10] | T763[10];
  assign T762[9] = T775[9] | T763[9];
  assign T762[8] = T775[8] | T763[8];
  assign T762[7] = T775[7] | T763[7];
  assign T762[6] = T775[6] | T763[6];
  assign T762[5] = T775[5] | T763[5];
  assign T762[4] = T775[4] | T763[4];
  assign T762[3] = T775[3] | T763[3];
  assign T762[2] = T775[2] | T763[2];
  assign T762[1] = T775[1] | T763[1];
  assign T762[0] = T775[0] | T763[0];
  assign T773 = io_uarch_counters_1 & T768[6];
  assign T775[63] = T788[63] | T776[63];
  assign T775[62] = T788[62] | T776[62];
  assign T775[61] = T788[61] | T776[61];
  assign T775[60] = T788[60] | T776[60];
  assign T775[59] = T788[59] | T776[59];
  assign T775[58] = T788[58] | T776[58];
  assign T775[57] = T788[57] | T776[57];
  assign T775[56] = T788[56] | T776[56];
  assign T775[55] = T788[55] | T776[55];
  assign T775[54] = T788[54] | T776[54];
  assign T775[53] = T788[53] | T776[53];
  assign T775[52] = T788[52] | T776[52];
  assign T775[51] = T788[51] | T776[51];
  assign T775[50] = T788[50] | T776[50];
  assign T775[49] = T788[49] | T776[49];
  assign T775[48] = T788[48] | T776[48];
  assign T775[47] = T788[47] | T776[47];
  assign T775[46] = T788[46] | T776[46];
  assign T775[45] = T788[45] | T776[45];
  assign T775[44] = T788[44] | T776[44];
  assign T775[43] = T788[43] | T776[43];
  assign T775[42] = T788[42] | T776[42];
  assign T775[41] = T788[41] | T776[41];
  assign T775[40] = T788[40] | T776[40];
  assign T775[39] = T788[39] | T776[39];
  assign T775[38] = T788[38] | T776[38];
  assign T775[37] = T788[37] | T776[37];
  assign T775[36] = T788[36] | T776[36];
  assign T775[35] = T788[35] | T776[35];
  assign T775[34] = T788[34] | T776[34];
  assign T775[33] = T788[33] | T776[33];
  assign T775[32] = T788[32] | T776[32];
  assign T775[31] = T788[31] | T776[31];
  assign T775[30] = T788[30] | T776[30];
  assign T775[29] = T788[29] | T776[29];
  assign T775[28] = T788[28] | T776[28];
  assign T775[27] = T788[27] | T776[27];
  assign T775[26] = T788[26] | T776[26];
  assign T775[25] = T788[25] | T776[25];
  assign T775[24] = T788[24] | T776[24];
  assign T775[23] = T788[23] | T776[23];
  assign T775[22] = T788[22] | T776[22];
  assign T775[21] = T788[21] | T776[21];
  assign T775[20] = T788[20] | T776[20];
  assign T775[19] = T788[19] | T776[19];
  assign T775[18] = T788[18] | T776[18];
  assign T775[17] = T788[17] | T776[17];
  assign T775[16] = T788[16] | T776[16];
  assign T775[15] = T788[15] | T776[15];
  assign T775[14] = T788[14] | T776[14];
  assign T775[13] = T788[13] | T776[13];
  assign T775[12] = T788[12] | T776[12];
  assign T775[11] = T788[11] | T776[11];
  assign T775[10] = T788[10] | T776[10];
  assign T775[9] = T788[9] | T776[9];
  assign T775[8] = T788[8] | T776[8];
  assign T775[7] = T788[7] | T776[7];
  assign T775[6] = T788[6] | T776[6];
  assign T775[5] = T788[5] | T776[5];
  assign T775[4] = T788[4] | T776[4];
  assign T775[3] = T788[3] | T776[3];
  assign T775[2] = T788[2] | T776[2];
  assign T775[1] = T788[1] | T776[1];
  assign T775[0] = T788[0] | T776[0];
  assign T786 = io_uarch_counters_0 & T781[6];
  assign T788[63] = T806[63] | T789[63];
  assign T788[62] = T806[62] | T789[62];
  assign T788[61] = T806[61] | T789[61];
  assign T788[60] = T806[60] | T789[60];
  assign T788[59] = T806[59] | T789[59];
  assign T788[58] = T806[58] | T789[58];
  assign T788[57] = T806[57] | T789[57];
  assign T788[56] = T806[56] | T789[56];
  assign T788[55] = T806[55] | T789[55];
  assign T788[54] = T806[54] | T789[54];
  assign T788[53] = T806[53] | T789[53];
  assign T788[52] = T806[52] | T789[52];
  assign T788[51] = T806[51] | T789[51];
  assign T788[50] = T806[50] | T789[50];
  assign T788[49] = T806[49] | T789[49];
  assign T788[48] = T806[48] | T789[48];
  assign T788[47] = T806[47] | T789[47];
  assign T788[46] = T806[46] | T789[46];
  assign T788[45] = T806[45] | T789[45];
  assign T788[44] = T806[44] | T789[44];
  assign T788[43] = T806[43] | T789[43];
  assign T788[42] = T806[42] | T789[42];
  assign T788[41] = T806[41] | T789[41];
  assign T788[40] = T806[40] | T789[40];
  assign T788[39] = T806[39] | T789[39];
  assign T788[38] = T806[38] | T789[38];
  assign T788[37] = T806[37] | T789[37];
  assign T788[36] = T806[36] | T789[36];
  assign T788[35] = T806[35] | T789[35];
  assign T788[34] = T806[34] | T789[34];
  assign T788[33] = T806[33] | T789[33];
  assign T788[32] = T806[32] | T789[32];
  assign T788[31] = T806[31] | T789[31];
  assign T788[30] = T806[30] | T789[30];
  assign T788[29] = T806[29] | T789[29];
  assign T788[28] = T806[28] | T789[28];
  assign T788[27] = T806[27] | T789[27];
  assign T788[26] = T806[26] | T789[26];
  assign T788[25] = T806[25] | T789[25];
  assign T788[24] = T806[24] | T789[24];
  assign T788[23] = T806[23] | T789[23];
  assign T788[22] = T806[22] | T789[22];
  assign T788[21] = T806[21] | T789[21];
  assign T788[20] = T806[20] | T789[20];
  assign T788[19] = T806[19] | T789[19];
  assign T788[18] = T806[18] | T789[18];
  assign T788[17] = T806[17] | T789[17];
  assign T788[16] = T806[16] | T789[16];
  assign T788[15] = T806[15] | T789[15];
  assign T788[14] = T806[14] | T789[14];
  assign T788[13] = T806[13] | T789[13];
  assign T788[12] = T806[12] | T789[12];
  assign T788[11] = T806[11] | T789[11];
  assign T788[10] = T806[10] | T789[10];
  assign T788[9] = T806[9] | T789[9];
  assign T788[8] = T806[8] | T789[8];
  assign T788[7] = T806[7] | T789[7];
  assign T788[6] = T806[6] | T789[6];
  assign T788[5] = T806[5] | T789[5];
  assign T788[4] = T806[4] | T789[4];
  assign T788[3] = T806[3] | T789[3];
  assign T788[2] = T806[2] | T789[2];
  assign T788[1] = T806[1] | T789[1];
  assign T788[0] = T806[0] | T789[0];
  assign T798 = io_rocc_csr_wen & N2732;
  assign T803 = io_retire & T795[6];
  assign T806[63] = T808[63] | T807[63];
  assign T806[62] = T808[62] | T807[62];
  assign T806[61] = T808[61] | T807[61];
  assign T806[60] = T808[60] | T807[60];
  assign T806[59] = T808[59] | T807[59];
  assign T806[58] = T808[58] | T807[58];
  assign T806[57] = T808[57] | T807[57];
  assign T806[56] = T808[56] | T807[56];
  assign T806[55] = T808[55] | T807[55];
  assign T806[54] = T808[54] | T807[54];
  assign T806[53] = T808[53] | T807[53];
  assign T806[52] = T808[52] | T807[52];
  assign T806[51] = T808[51] | T807[51];
  assign T806[50] = T808[50] | T807[50];
  assign T806[49] = T808[49] | T807[49];
  assign T806[48] = T808[48] | T807[48];
  assign T806[47] = T808[47] | T807[47];
  assign T806[46] = T808[46] | T807[46];
  assign T806[45] = T808[45] | T807[45];
  assign T806[44] = T808[44] | T807[44];
  assign T806[43] = T808[43] | T807[43];
  assign T806[42] = T808[42] | T807[42];
  assign T806[41] = T808[41] | T807[41];
  assign T806[40] = T808[40] | T807[40];
  assign T806[39] = T808[39] | T807[39];
  assign T806[38] = T808[38] | T807[38];
  assign T806[37] = T808[37] | T807[37];
  assign T806[36] = T808[36] | T807[36];
  assign T806[35] = T808[35] | T807[35];
  assign T806[34] = T808[34] | T807[34];
  assign T806[33] = T808[33] | T807[33];
  assign T806[32] = T808[32] | T807[32];
  assign T806[31] = T808[31] | T807[31];
  assign T806[30] = T808[30] | T807[30];
  assign T806[29] = T808[29] | T807[29];
  assign T806[28] = T808[28] | T807[28];
  assign T806[27] = T808[27] | T807[27];
  assign T806[26] = T808[26] | T807[26];
  assign T806[25] = T808[25] | T807[25];
  assign T806[24] = T808[24] | T807[24];
  assign T806[23] = T808[23] | T807[23];
  assign T806[22] = T808[22] | T807[22];
  assign T806[21] = T808[21] | T807[21];
  assign T806[20] = T808[20] | T807[20];
  assign T806[19] = T808[19] | T807[19];
  assign T806[18] = T808[18] | T807[18];
  assign T806[17] = T808[17] | T807[17];
  assign T806[16] = T808[16] | T807[16];
  assign T806[15] = T808[15] | T807[15];
  assign T806[14] = T808[14] | T807[14];
  assign T806[13] = T808[13] | T807[13];
  assign T806[12] = T808[12] | T807[12];
  assign T806[11] = T808[11] | T807[11];
  assign T806[10] = T808[10] | T807[10];
  assign T806[9] = T808[9] | T807[9];
  assign T806[8] = T808[8] | T807[8];
  assign T806[7] = T808[7] | T807[7];
  assign T806[6] = T808[6] | T807[6];
  assign T806[5] = T808[5] | T807[5];
  assign T806[4] = T808[4] | T807[4];
  assign T806[3] = T808[3] | T807[3];
  assign T806[2] = T808[2] | T807[2];
  assign T806[1] = T808[1] | T807[1];
  assign T806[0] = T808[0] | T807[0];
  assign T808[63] = T810[63] | T809[63];
  assign T808[62] = T810[62] | T809[62];
  assign T808[61] = T810[61] | T809[61];
  assign T808[60] = T810[60] | T809[60];
  assign T808[59] = T810[59] | T809[59];
  assign T808[58] = T810[58] | T809[58];
  assign T808[57] = T810[57] | T809[57];
  assign T808[56] = T810[56] | T809[56];
  assign T808[55] = T810[55] | T809[55];
  assign T808[54] = T810[54] | T809[54];
  assign T808[53] = T810[53] | T809[53];
  assign T808[52] = T810[52] | T809[52];
  assign T808[51] = T810[51] | T809[51];
  assign T808[50] = T810[50] | T809[50];
  assign T808[49] = T810[49] | T809[49];
  assign T808[48] = T810[48] | T809[48];
  assign T808[47] = T810[47] | T809[47];
  assign T808[46] = T810[46] | T809[46];
  assign T808[45] = T810[45] | T809[45];
  assign T808[44] = T810[44] | T809[44];
  assign T808[43] = T810[43] | T809[43];
  assign T808[42] = T810[42] | T809[42];
  assign T808[41] = T810[41] | T809[41];
  assign T808[40] = T810[40] | T809[40];
  assign T808[39] = T810[39] | T809[39];
  assign T808[38] = T810[38] | T809[38];
  assign T808[37] = T810[37] | T809[37];
  assign T808[36] = T810[36] | T809[36];
  assign T808[35] = T810[35] | T809[35];
  assign T808[34] = T810[34] | T809[34];
  assign T808[33] = T810[33] | T809[33];
  assign T808[32] = T810[32] | T809[32];
  assign T808[31] = T810[31] | T809[31];
  assign T808[30] = T810[30] | T809[30];
  assign T808[29] = T810[29] | T809[29];
  assign T808[28] = T810[28] | T809[28];
  assign T808[27] = T810[27] | T809[27];
  assign T808[26] = T810[26] | T809[26];
  assign T808[25] = T810[25] | T809[25];
  assign T808[24] = T810[24] | T809[24];
  assign T808[23] = T810[23] | T809[23];
  assign T808[22] = T810[22] | T809[22];
  assign T808[21] = T810[21] | T809[21];
  assign T808[20] = T810[20] | T809[20];
  assign T808[19] = T810[19] | T809[19];
  assign T808[18] = T810[18] | T809[18];
  assign T808[17] = T810[17] | T809[17];
  assign T808[16] = T810[16] | T809[16];
  assign T808[15] = T810[15] | T809[15];
  assign T808[14] = T810[14] | T809[14];
  assign T808[13] = T810[13] | T809[13];
  assign T808[12] = T810[12] | T809[12];
  assign T808[11] = T810[11] | T809[11];
  assign T808[10] = T810[10] | T809[10];
  assign T808[9] = T810[9] | T809[9];
  assign T808[8] = T810[8] | T809[8];
  assign T808[7] = T810[7] | T809[7];
  assign T808[6] = T810[6] | T809[6];
  assign T808[5] = T810[5] | T809[5];
  assign T808[4] = T810[4] | T809[4];
  assign T808[3] = T810[3] | T809[3];
  assign T808[2] = T810[2] | T809[2];
  assign T808[1] = T810[1] | T809[1];
  assign T808[0] = T810[0] | T809[0];
  assign T810[63] = T821[63] | T811[63];
  assign T810[62] = T821[62] | T811[62];
  assign T810[61] = T821[61] | T811[61];
  assign T810[60] = T821[60] | T811[60];
  assign T810[59] = T821[59] | T811[59];
  assign T810[58] = T821[58] | T811[58];
  assign T810[57] = T821[57] | T811[57];
  assign T810[56] = T821[56] | T811[56];
  assign T810[55] = T821[55] | T811[55];
  assign T810[54] = T821[54] | T811[54];
  assign T810[53] = T821[53] | T811[53];
  assign T810[52] = T821[52] | T811[52];
  assign T810[51] = T821[51] | T811[51];
  assign T810[50] = T821[50] | T811[50];
  assign T810[49] = T821[49] | T811[49];
  assign T810[48] = T821[48] | T811[48];
  assign T810[47] = T821[47] | T811[47];
  assign T810[46] = T821[46] | T811[46];
  assign T810[45] = T821[45] | T811[45];
  assign T810[44] = T821[44] | T811[44];
  assign T810[43] = T821[43] | T811[43];
  assign T810[42] = T821[42] | T811[42];
  assign T810[41] = T821[41] | T811[41];
  assign T810[40] = T821[40] | T811[40];
  assign T810[39] = T821[39] | T811[39];
  assign T810[38] = T821[38] | T811[38];
  assign T810[37] = T821[37] | T811[37];
  assign T810[36] = T821[36] | T811[36];
  assign T810[35] = T821[35] | T811[35];
  assign T810[34] = T821[34] | T811[34];
  assign T810[33] = T821[33] | T811[33];
  assign T810[32] = T821[32] | T811[32];
  assign T810[31] = T821[31] | T811[31];
  assign T810[30] = T821[30] | T811[30];
  assign T810[29] = T821[29] | T811[29];
  assign T810[28] = T821[28] | T811[28];
  assign T810[27] = T821[27] | T811[27];
  assign T810[26] = T821[26] | T811[26];
  assign T810[25] = T821[25] | T811[25];
  assign T810[24] = T821[24] | T811[24];
  assign T810[23] = T821[23] | T811[23];
  assign T810[22] = T821[22] | T811[22];
  assign T810[21] = T821[21] | T811[21];
  assign T810[20] = T821[20] | T811[20];
  assign T810[19] = T821[19] | T811[19];
  assign T810[18] = T821[18] | T811[18];
  assign T810[17] = T821[17] | T811[17];
  assign T810[16] = T821[16] | T811[16];
  assign T810[15] = T821[15] | T811[15];
  assign T810[14] = T821[14] | T811[14];
  assign T810[13] = T821[13] | T811[13];
  assign T810[12] = T821[12] | T811[12];
  assign T810[11] = T821[11] | T811[11];
  assign T810[10] = T821[10] | T811[10];
  assign T810[9] = T821[9] | T811[9];
  assign T810[8] = T821[8] | T811[8];
  assign T810[7] = T821[7] | T811[7];
  assign T810[6] = T821[6] | T811[6];
  assign T810[5] = T821[5] | T811[5];
  assign T810[4] = T821[4] | T811[4];
  assign T810[3] = T821[3] | T811[3];
  assign T810[2] = T821[2] | T811[2];
  assign T810[1] = T821[1] | T811[1];
  assign T810[0] = T821[0] | T811[0];
  assign T814 = T815 & N2769;
  assign T815 = host_csr_req_fire & T816;
  assign T816 = ~host_csr_bits_rw;
  assign T817 = T820 & T818;
  assign T818 = N2290 | host_csr_req_fire;
  assign T820 = io_rocc_csr_wen & N2769;
  assign T821[63] = T826[63] | 1'b0;
  assign T821[62] = T826[62] | 1'b0;
  assign T821[61] = T826[61] | 1'b0;
  assign T821[60] = T826[60] | 1'b0;
  assign T821[59] = T826[59] | 1'b0;
  assign T821[58] = T826[58] | 1'b0;
  assign T821[57] = T826[57] | 1'b0;
  assign T821[56] = T826[56] | 1'b0;
  assign T821[55] = T826[55] | 1'b0;
  assign T821[54] = T826[54] | 1'b0;
  assign T821[53] = T826[53] | 1'b0;
  assign T821[52] = T826[52] | 1'b0;
  assign T821[51] = T826[51] | 1'b0;
  assign T821[50] = T826[50] | 1'b0;
  assign T821[49] = T826[49] | 1'b0;
  assign T821[48] = T826[48] | 1'b0;
  assign T821[47] = T826[47] | 1'b0;
  assign T821[46] = T826[46] | 1'b0;
  assign T821[45] = T826[45] | 1'b0;
  assign T821[44] = T826[44] | 1'b0;
  assign T821[43] = T826[43] | 1'b0;
  assign T821[42] = T826[42] | 1'b0;
  assign T821[41] = T826[41] | 1'b0;
  assign T821[40] = T826[40] | 1'b0;
  assign T821[39] = T826[39] | 1'b0;
  assign T821[38] = T826[38] | 1'b0;
  assign T821[37] = T826[37] | 1'b0;
  assign T821[36] = T826[36] | 1'b0;
  assign T821[35] = T826[35] | 1'b0;
  assign T821[34] = T826[34] | 1'b0;
  assign T821[33] = T826[33] | 1'b0;
  assign T821[32] = T826[32] | 1'b0;
  assign T821[31] = T826[31] | 1'b0;
  assign T821[30] = T826[30] | 1'b0;
  assign T821[29] = T826[29] | 1'b0;
  assign T821[28] = T826[28] | 1'b0;
  assign T821[27] = T826[27] | 1'b0;
  assign T821[26] = T826[26] | 1'b0;
  assign T821[25] = T826[25] | 1'b0;
  assign T821[24] = T826[24] | 1'b0;
  assign T821[23] = T826[23] | 1'b0;
  assign T821[22] = T826[22] | 1'b0;
  assign T821[21] = T826[21] | 1'b0;
  assign T821[20] = T826[20] | 1'b0;
  assign T821[19] = T826[19] | 1'b0;
  assign T821[18] = T826[18] | 1'b0;
  assign T821[17] = T826[17] | 1'b0;
  assign T821[16] = T826[16] | 1'b0;
  assign T821[15] = T826[15] | 1'b0;
  assign T821[14] = T826[14] | 1'b0;
  assign T821[13] = T826[13] | 1'b0;
  assign T821[12] = T826[12] | 1'b0;
  assign T821[11] = T826[11] | 1'b0;
  assign T821[10] = T826[10] | 1'b0;
  assign T821[9] = T826[9] | 1'b0;
  assign T821[8] = T826[8] | 1'b0;
  assign T821[7] = T826[7] | 1'b0;
  assign T821[6] = T826[6] | 1'b0;
  assign T821[5] = T826[5] | 1'b0;
  assign T821[4] = T826[4] | 1'b0;
  assign T821[3] = T826[3] | 1'b0;
  assign T821[2] = T826[2] | 1'b0;
  assign T821[1] = T826[1] | 1'b0;
  assign T821[0] = T826[0] | T1003[0];
  assign T825 = io_rocc_csr_wen & N2781;
  assign T826[63] = T828[63] | 1'b0;
  assign T826[62] = T828[62] | 1'b0;
  assign T826[61] = T828[61] | 1'b0;
  assign T826[60] = T828[60] | 1'b0;
  assign T826[59] = T828[59] | 1'b0;
  assign T826[58] = T828[58] | 1'b0;
  assign T826[57] = T828[57] | 1'b0;
  assign T826[56] = T828[56] | 1'b0;
  assign T826[55] = T828[55] | 1'b0;
  assign T826[54] = T828[54] | 1'b0;
  assign T826[53] = T828[53] | 1'b0;
  assign T826[52] = T828[52] | 1'b0;
  assign T826[51] = T828[51] | 1'b0;
  assign T826[50] = T828[50] | 1'b0;
  assign T826[49] = T828[49] | 1'b0;
  assign T826[48] = T828[48] | 1'b0;
  assign T826[47] = T828[47] | 1'b0;
  assign T826[46] = T828[46] | 1'b0;
  assign T826[45] = T828[45] | 1'b0;
  assign T826[44] = T828[44] | 1'b0;
  assign T826[43] = T828[43] | 1'b0;
  assign T826[42] = T828[42] | 1'b0;
  assign T826[41] = T828[41] | 1'b0;
  assign T826[40] = T828[40] | 1'b0;
  assign T826[39] = T828[39] | 1'b0;
  assign T826[38] = T828[38] | 1'b0;
  assign T826[37] = T828[37] | 1'b0;
  assign T826[36] = T828[36] | 1'b0;
  assign T826[35] = T828[35] | 1'b0;
  assign T826[34] = T828[34] | 1'b0;
  assign T826[33] = T828[33] | 1'b0;
  assign T826[32] = T828[32] | 1'b0;
  assign T826[31] = T828[31] | 1'b0;
  assign T826[30] = T828[30] | 1'b0;
  assign T826[29] = T828[29] | 1'b0;
  assign T826[28] = T828[28] | 1'b0;
  assign T826[27] = T828[27] | 1'b0;
  assign T826[26] = T828[26] | 1'b0;
  assign T826[25] = T828[25] | 1'b0;
  assign T826[24] = T828[24] | 1'b0;
  assign T826[23] = T828[23] | 1'b0;
  assign T826[22] = T828[22] | 1'b0;
  assign T826[21] = T828[21] | 1'b0;
  assign T826[20] = T828[20] | 1'b0;
  assign T826[19] = T828[19] | 1'b0;
  assign T826[18] = T828[18] | 1'b0;
  assign T826[17] = T828[17] | 1'b0;
  assign T826[16] = T828[16] | 1'b0;
  assign T826[15] = T828[15] | 1'b0;
  assign T826[14] = T828[14] | 1'b0;
  assign T826[13] = T828[13] | 1'b0;
  assign T826[12] = T828[12] | 1'b0;
  assign T826[11] = T828[11] | 1'b0;
  assign T826[10] = T828[10] | 1'b0;
  assign T826[9] = T828[9] | 1'b0;
  assign T826[8] = T828[8] | 1'b0;
  assign T826[7] = T828[7] | 1'b0;
  assign T826[6] = T828[6] | 1'b0;
  assign T826[5] = T828[5] | 1'b0;
  assign T826[4] = T828[4] | 1'b0;
  assign T826[3] = T828[3] | 1'b0;
  assign T826[2] = T828[2] | 1'b0;
  assign T826[1] = T828[1] | 1'b0;
  assign T826[0] = T828[0] | T1005[0];
  assign T828[63] = T830[63] | T829[63];
  assign T828[62] = T830[62] | T829[62];
  assign T828[61] = T830[61] | T829[61];
  assign T828[60] = T830[60] | T829[60];
  assign T828[59] = T830[59] | T829[59];
  assign T828[58] = T830[58] | T829[58];
  assign T828[57] = T830[57] | T829[57];
  assign T828[56] = T830[56] | T829[56];
  assign T828[55] = T830[55] | T829[55];
  assign T828[54] = T830[54] | T829[54];
  assign T828[53] = T830[53] | T829[53];
  assign T828[52] = T830[52] | T829[52];
  assign T828[51] = T830[51] | T829[51];
  assign T828[50] = T830[50] | T829[50];
  assign T828[49] = T830[49] | T829[49];
  assign T828[48] = T830[48] | T829[48];
  assign T828[47] = T830[47] | T829[47];
  assign T828[46] = T830[46] | T829[46];
  assign T828[45] = T830[45] | T829[45];
  assign T828[44] = T830[44] | T829[44];
  assign T828[43] = T830[43] | T829[43];
  assign T828[42] = T830[42] | T829[42];
  assign T828[41] = T830[41] | T829[41];
  assign T828[40] = T830[40] | T829[40];
  assign T828[39] = T830[39] | T829[39];
  assign T828[38] = T830[38] | T829[38];
  assign T828[37] = T830[37] | T829[37];
  assign T828[36] = T830[36] | T829[36];
  assign T828[35] = T830[35] | T829[35];
  assign T828[34] = T830[34] | T829[34];
  assign T828[33] = T830[33] | T829[33];
  assign T828[32] = T830[32] | T829[32];
  assign T828[31] = T830[31] | T829[31];
  assign T828[30] = T830[30] | T829[30];
  assign T828[29] = T830[29] | T829[29];
  assign T828[28] = T830[28] | T829[28];
  assign T828[27] = T830[27] | T829[27];
  assign T828[26] = T830[26] | T829[26];
  assign T828[25] = T830[25] | T829[25];
  assign T828[24] = T830[24] | T829[24];
  assign T828[23] = T830[23] | T829[23];
  assign T828[22] = T830[22] | T829[22];
  assign T828[21] = T830[21] | T829[21];
  assign T828[20] = T830[20] | T829[20];
  assign T828[19] = T830[19] | T829[19];
  assign T828[18] = T830[18] | T829[18];
  assign T828[17] = T830[17] | T829[17];
  assign T828[16] = T830[16] | T829[16];
  assign T828[15] = T830[15] | T829[15];
  assign T828[14] = T830[14] | T829[14];
  assign T828[13] = T830[13] | T829[13];
  assign T828[12] = T830[12] | T829[12];
  assign T828[11] = T830[11] | T829[11];
  assign T828[10] = T830[10] | T829[10];
  assign T828[9] = T830[9] | T829[9];
  assign T828[8] = T830[8] | T829[8];
  assign T828[7] = T830[7] | T829[7];
  assign T828[6] = T830[6] | T829[6];
  assign T828[5] = T830[5] | T829[5];
  assign T828[4] = T830[4] | T829[4];
  assign T828[3] = T830[3] | T829[3];
  assign T828[2] = T830[2] | T829[2];
  assign T828[1] = T830[1] | T829[1];
  assign T828[0] = T830[0] | T829[0];
  assign T830[63] = T832[63] | T831[63];
  assign T830[62] = T832[62] | T831[62];
  assign T830[61] = T832[61] | T831[61];
  assign T830[60] = T832[60] | T831[60];
  assign T830[59] = T832[59] | T831[59];
  assign T830[58] = T832[58] | T831[58];
  assign T830[57] = T832[57] | T831[57];
  assign T830[56] = T832[56] | T831[56];
  assign T830[55] = T832[55] | T831[55];
  assign T830[54] = T832[54] | T831[54];
  assign T830[53] = T832[53] | T831[53];
  assign T830[52] = T832[52] | T831[52];
  assign T830[51] = T832[51] | T831[51];
  assign T830[50] = T832[50] | T831[50];
  assign T830[49] = T832[49] | T831[49];
  assign T830[48] = T832[48] | T831[48];
  assign T830[47] = T832[47] | T831[47];
  assign T830[46] = T832[46] | T831[46];
  assign T830[45] = T832[45] | T831[45];
  assign T830[44] = T832[44] | T831[44];
  assign T830[43] = T832[43] | T831[43];
  assign T830[42] = T832[42] | T831[42];
  assign T830[41] = T832[41] | T831[41];
  assign T830[40] = T832[40] | T831[40];
  assign T830[39] = T832[39] | T831[39];
  assign T830[38] = T832[38] | T831[38];
  assign T830[37] = T832[37] | T831[37];
  assign T830[36] = T832[36] | T831[36];
  assign T830[35] = T832[35] | T831[35];
  assign T830[34] = T832[34] | T831[34];
  assign T830[33] = T832[33] | T831[33];
  assign T830[32] = T832[32] | T831[32];
  assign T830[31] = T832[31] | T831[31];
  assign T830[30] = T832[30] | T831[30];
  assign T830[29] = T832[29] | T831[29];
  assign T830[28] = T832[28] | T831[28];
  assign T830[27] = T832[27] | T831[27];
  assign T830[26] = T832[26] | T831[26];
  assign T830[25] = T832[25] | T831[25];
  assign T830[24] = T832[24] | T831[24];
  assign T830[23] = T832[23] | T831[23];
  assign T830[22] = T832[22] | T831[22];
  assign T830[21] = T832[21] | T831[21];
  assign T830[20] = T832[20] | T831[20];
  assign T830[19] = T832[19] | T831[19];
  assign T830[18] = T832[18] | T831[18];
  assign T830[17] = T832[17] | T831[17];
  assign T830[16] = T832[16] | T831[16];
  assign T830[15] = T832[15] | T831[15];
  assign T830[14] = T832[14] | T831[14];
  assign T830[13] = T832[13] | T831[13];
  assign T830[12] = T832[12] | T831[12];
  assign T830[11] = T832[11] | T831[11];
  assign T830[10] = T832[10] | T831[10];
  assign T830[9] = T832[9] | T831[9];
  assign T830[8] = T832[8] | T831[8];
  assign T830[7] = T832[7] | T831[7];
  assign T830[6] = T832[6] | T831[6];
  assign T830[5] = T832[5] | T831[5];
  assign T830[4] = T832[4] | T831[4];
  assign T830[3] = T832[3] | T831[3];
  assign T830[2] = T832[2] | T831[2];
  assign T830[1] = T832[1] | T831[1];
  assign T830[0] = T832[0] | T831[0];
  assign T832[63] = T837[63] | T833[63];
  assign T832[62] = T837[62] | T833[62];
  assign T832[61] = T837[61] | T833[61];
  assign T832[60] = T837[60] | T833[60];
  assign T832[59] = T837[59] | T833[59];
  assign T832[58] = T837[58] | T833[58];
  assign T832[57] = T837[57] | T833[57];
  assign T832[56] = T837[56] | T833[56];
  assign T832[55] = T837[55] | T833[55];
  assign T832[54] = T837[54] | T833[54];
  assign T832[53] = T837[53] | T833[53];
  assign T832[52] = T837[52] | T833[52];
  assign T832[51] = T837[51] | T833[51];
  assign T832[50] = T837[50] | T833[50];
  assign T832[49] = T837[49] | T833[49];
  assign T832[48] = T837[48] | T833[48];
  assign T832[47] = T837[47] | T833[47];
  assign T832[46] = T837[46] | T833[46];
  assign T832[45] = T837[45] | T833[45];
  assign T832[44] = T837[44] | T833[44];
  assign T832[43] = T837[43] | T833[43];
  assign T832[42] = T837[42] | T833[42];
  assign T832[41] = T837[41] | T833[41];
  assign T832[40] = T837[40] | T833[40];
  assign T832[39] = T837[39] | T833[39];
  assign T832[38] = T837[38] | T833[38];
  assign T832[37] = T837[37] | T833[37];
  assign T832[36] = T837[36] | T833[36];
  assign T832[35] = T837[35] | T833[35];
  assign T832[34] = T837[34] | T833[34];
  assign T832[33] = T837[33] | T833[33];
  assign T832[32] = T837[32] | T833[32];
  assign T832[31] = T837[31] | T833[31];
  assign T832[30] = T837[30] | T833[30];
  assign T832[29] = T837[29] | T833[29];
  assign T832[28] = T837[28] | T833[28];
  assign T832[27] = T837[27] | T833[27];
  assign T832[26] = T837[26] | T833[26];
  assign T832[25] = T837[25] | T833[25];
  assign T832[24] = T837[24] | T833[24];
  assign T832[23] = T837[23] | T833[23];
  assign T832[22] = T837[22] | T833[22];
  assign T832[21] = T837[21] | T833[21];
  assign T832[20] = T837[20] | T833[20];
  assign T832[19] = T837[19] | T833[19];
  assign T832[18] = T837[18] | T833[18];
  assign T832[17] = T837[17] | T833[17];
  assign T832[16] = T837[16] | T833[16];
  assign T832[15] = T837[15] | T833[15];
  assign T832[14] = T837[14] | T833[14];
  assign T832[13] = T837[13] | T833[13];
  assign T832[12] = T837[12] | T833[12];
  assign T832[11] = T837[11] | T833[11];
  assign T832[10] = T837[10] | T833[10];
  assign T832[9] = T837[9] | T833[9];
  assign T832[8] = T837[8] | T833[8];
  assign T832[7] = T837[7] | T833[7];
  assign T832[6] = T837[6] | T833[6];
  assign T832[5] = T837[5] | T833[5];
  assign T832[4] = T837[4] | T833[4];
  assign T832[3] = T837[3] | T833[3];
  assign T832[2] = T837[2] | T833[2];
  assign T832[1] = T837[1] | T833[1];
  assign T832[0] = T837[0] | T833[0];
  assign T837[63] = T842[63] | T838[63];
  assign T837[62] = T842[62] | T838[62];
  assign T837[61] = T842[61] | T838[61];
  assign T837[60] = T842[60] | T838[60];
  assign T837[59] = T842[59] | T838[59];
  assign T837[58] = T842[58] | T838[58];
  assign T837[57] = T842[57] | T838[57];
  assign T837[56] = T842[56] | T838[56];
  assign T837[55] = T842[55] | T838[55];
  assign T837[54] = T842[54] | T838[54];
  assign T837[53] = T842[53] | T838[53];
  assign T837[52] = T842[52] | T838[52];
  assign T837[51] = T842[51] | T838[51];
  assign T837[50] = T842[50] | T838[50];
  assign T837[49] = T842[49] | T838[49];
  assign T837[48] = T842[48] | T838[48];
  assign T837[47] = T842[47] | T838[47];
  assign T837[46] = T842[46] | T838[46];
  assign T837[45] = T842[45] | T838[45];
  assign T837[44] = T842[44] | T838[44];
  assign T837[43] = T842[43] | T838[43];
  assign T837[42] = T842[42] | T838[42];
  assign T837[41] = T842[41] | T838[41];
  assign T837[40] = T842[40] | T838[40];
  assign T837[39] = T842[39] | T838[39];
  assign T837[38] = T842[38] | T838[38];
  assign T837[37] = T842[37] | T838[37];
  assign T837[36] = T842[36] | T838[36];
  assign T837[35] = T842[35] | T838[35];
  assign T837[34] = T842[34] | T838[34];
  assign T837[33] = T842[33] | T838[33];
  assign T837[32] = T842[32] | T838[32];
  assign T837[31] = T842[31] | T838[31];
  assign T837[30] = T842[30] | T838[30];
  assign T837[29] = T842[29] | T838[29];
  assign T837[28] = T842[28] | T838[28];
  assign T837[27] = T842[27] | T838[27];
  assign T837[26] = T842[26] | T838[26];
  assign T837[25] = T842[25] | T838[25];
  assign T837[24] = T842[24] | T838[24];
  assign T837[23] = T842[23] | T838[23];
  assign T837[22] = T842[22] | T838[22];
  assign T837[21] = T842[21] | T838[21];
  assign T837[20] = T842[20] | T838[20];
  assign T837[19] = T842[19] | T838[19];
  assign T837[18] = T842[18] | T838[18];
  assign T837[17] = T842[17] | T838[17];
  assign T837[16] = T842[16] | T838[16];
  assign T837[15] = T842[15] | T838[15];
  assign T837[14] = T842[14] | T838[14];
  assign T837[13] = T842[13] | T838[13];
  assign T837[12] = T842[12] | T838[12];
  assign T837[11] = T842[11] | T838[11];
  assign T837[10] = T842[10] | T838[10];
  assign T837[9] = T842[9] | T838[9];
  assign T837[8] = T842[8] | T838[8];
  assign T837[7] = T842[7] | T838[7];
  assign T837[6] = T842[6] | T838[6];
  assign T837[5] = T842[5] | T838[5];
  assign T837[4] = T842[4] | T838[4];
  assign T837[3] = T842[3] | T838[3];
  assign T837[2] = T842[2] | T838[2];
  assign T837[1] = T842[1] | T838[1];
  assign T837[0] = T842[0] | T838[0];
  assign T842[63] = T846[63] | T843[63];
  assign T842[62] = T846[62] | T843[62];
  assign T842[61] = T846[61] | T843[61];
  assign T842[60] = T846[60] | T843[60];
  assign T842[59] = T846[59] | T843[59];
  assign T842[58] = T846[58] | T843[58];
  assign T842[57] = T846[57] | T843[57];
  assign T842[56] = T846[56] | T843[56];
  assign T842[55] = T846[55] | T843[55];
  assign T842[54] = T846[54] | T843[54];
  assign T842[53] = T846[53] | T843[53];
  assign T842[52] = T846[52] | T843[52];
  assign T842[51] = T846[51] | T843[51];
  assign T842[50] = T846[50] | T843[50];
  assign T842[49] = T846[49] | T843[49];
  assign T842[48] = T846[48] | T843[48];
  assign T842[47] = T846[47] | T843[47];
  assign T842[46] = T846[46] | T843[46];
  assign T842[45] = T846[45] | T843[45];
  assign T842[44] = T846[44] | T843[44];
  assign T842[43] = T846[43] | T843[43];
  assign T842[42] = T846[42] | T843[42];
  assign T842[41] = T846[41] | T843[41];
  assign T842[40] = T846[40] | T843[40];
  assign T842[39] = T846[39] | T843[39];
  assign T842[38] = T846[38] | T843[38];
  assign T842[37] = T846[37] | T843[37];
  assign T842[36] = T846[36] | T843[36];
  assign T842[35] = T846[35] | T843[35];
  assign T842[34] = T846[34] | T843[34];
  assign T842[33] = T846[33] | T843[33];
  assign T842[32] = T846[32] | T843[32];
  assign T842[31] = T846[31] | T843[31];
  assign T842[30] = T846[30] | T843[30];
  assign T842[29] = T846[29] | T843[29];
  assign T842[28] = T846[28] | T843[28];
  assign T842[27] = T846[27] | T843[27];
  assign T842[26] = T846[26] | T843[26];
  assign T842[25] = T846[25] | T843[25];
  assign T842[24] = T846[24] | T843[24];
  assign T842[23] = T846[23] | T843[23];
  assign T842[22] = T846[22] | T843[22];
  assign T842[21] = T846[21] | T843[21];
  assign T842[20] = T846[20] | T843[20];
  assign T842[19] = T846[19] | T843[19];
  assign T842[18] = T846[18] | T843[18];
  assign T842[17] = T846[17] | T843[17];
  assign T842[16] = T846[16] | T843[16];
  assign T842[15] = T846[15] | T843[15];
  assign T842[14] = T846[14] | T843[14];
  assign T842[13] = T846[13] | T843[13];
  assign T842[12] = T846[12] | T843[12];
  assign T842[11] = T846[11] | T843[11];
  assign T842[10] = T846[10] | T843[10];
  assign T842[9] = T846[9] | T843[9];
  assign T842[8] = T846[8] | T843[8];
  assign T842[7] = T846[7] | T843[7];
  assign T842[6] = T846[6] | T843[6];
  assign T842[5] = T846[5] | T843[5];
  assign T842[4] = T846[4] | T843[4];
  assign T842[3] = T846[3] | T843[3];
  assign T842[2] = T846[2] | T843[2];
  assign T842[1] = T846[1] | T843[1];
  assign T842[0] = T846[0] | T843[0];
  assign T845 = io_rocc_csr_wen & N2857;
  assign T846[63] = T856[63] | 1'b0;
  assign T846[62] = T856[62] | 1'b0;
  assign T846[61] = T856[61] | 1'b0;
  assign T846[60] = T856[60] | 1'b0;
  assign T846[59] = T856[59] | 1'b0;
  assign T846[58] = T856[58] | 1'b0;
  assign T846[57] = T856[57] | 1'b0;
  assign T846[56] = T856[56] | 1'b0;
  assign T846[55] = T856[55] | 1'b0;
  assign T846[54] = T856[54] | 1'b0;
  assign T846[53] = T856[53] | 1'b0;
  assign T846[52] = T856[52] | 1'b0;
  assign T846[51] = T856[51] | 1'b0;
  assign T846[50] = T856[50] | 1'b0;
  assign T846[49] = T856[49] | 1'b0;
  assign T846[48] = T856[48] | 1'b0;
  assign T846[47] = T856[47] | 1'b0;
  assign T846[46] = T856[46] | 1'b0;
  assign T846[45] = T856[45] | 1'b0;
  assign T846[44] = T856[44] | 1'b0;
  assign T846[43] = T856[43] | 1'b0;
  assign T846[42] = T856[42] | 1'b0;
  assign T846[41] = T856[41] | 1'b0;
  assign T846[40] = T856[40] | 1'b0;
  assign T846[39] = T856[39] | 1'b0;
  assign T846[38] = T856[38] | 1'b0;
  assign T846[37] = T856[37] | 1'b0;
  assign T846[36] = T856[36] | 1'b0;
  assign T846[35] = T856[35] | 1'b0;
  assign T846[34] = T856[34] | 1'b0;
  assign T846[33] = T856[33] | 1'b0;
  assign T846[32] = T856[32] | 1'b0;
  assign T846[31] = T856[31] | 1'b0;
  assign T846[30] = T856[30] | 1'b0;
  assign T846[29] = T856[29] | 1'b0;
  assign T846[28] = T856[28] | 1'b0;
  assign T846[27] = T856[27] | 1'b0;
  assign T846[26] = T856[26] | 1'b0;
  assign T846[25] = T856[25] | 1'b0;
  assign T846[24] = T856[24] | 1'b0;
  assign T846[23] = T856[23] | 1'b0;
  assign T846[22] = T856[22] | 1'b0;
  assign T846[21] = T856[21] | 1'b0;
  assign T846[20] = T856[20] | 1'b0;
  assign T846[19] = T856[19] | 1'b0;
  assign T846[18] = T856[18] | 1'b0;
  assign T846[17] = T856[17] | 1'b0;
  assign T846[16] = T856[16] | 1'b0;
  assign T846[15] = T856[15] | 1'b0;
  assign T846[14] = T856[14] | 1'b0;
  assign T846[13] = T856[13] | 1'b0;
  assign T846[12] = T856[12] | 1'b0;
  assign T846[11] = T856[11] | 1'b0;
  assign T846[10] = T856[10] | 1'b0;
  assign T846[9] = T856[9] | 1'b0;
  assign T846[8] = T856[8] | 1'b0;
  assign T846[7] = T856[7] | T1008[7];
  assign T846[6] = T856[6] | T1008[6];
  assign T846[5] = T856[5] | T1008[5];
  assign T846[4] = T856[4] | T1008[4];
  assign T846[3] = T856[3] | T1008[3];
  assign T846[2] = T856[2] | T1008[2];
  assign T846[1] = T856[1] | T1008[1];
  assign T846[0] = T856[0] | T1008[0];
  assign T856[63] = T866[63] | 1'b0;
  assign T856[62] = T866[62] | 1'b0;
  assign T856[61] = T866[61] | 1'b0;
  assign T856[60] = T866[60] | 1'b0;
  assign T856[59] = T866[59] | 1'b0;
  assign T856[58] = T866[58] | 1'b0;
  assign T856[57] = T866[57] | 1'b0;
  assign T856[56] = T866[56] | 1'b0;
  assign T856[55] = T866[55] | 1'b0;
  assign T856[54] = T866[54] | 1'b0;
  assign T856[53] = T866[53] | 1'b0;
  assign T856[52] = T866[52] | 1'b0;
  assign T856[51] = T866[51] | 1'b0;
  assign T856[50] = T866[50] | 1'b0;
  assign T856[49] = T866[49] | 1'b0;
  assign T856[48] = T866[48] | 1'b0;
  assign T856[47] = T866[47] | 1'b0;
  assign T856[46] = T866[46] | 1'b0;
  assign T856[45] = T866[45] | 1'b0;
  assign T856[44] = T866[44] | 1'b0;
  assign T856[43] = T866[43] | 1'b0;
  assign T856[42] = T866[42] | 1'b0;
  assign T856[41] = T866[41] | 1'b0;
  assign T856[40] = T866[40] | 1'b0;
  assign T856[39] = T866[39] | 1'b0;
  assign T856[38] = T866[38] | 1'b0;
  assign T856[37] = T866[37] | 1'b0;
  assign T856[36] = T866[36] | 1'b0;
  assign T856[35] = T866[35] | 1'b0;
  assign T856[34] = T866[34] | 1'b0;
  assign T856[33] = T866[33] | 1'b0;
  assign T856[32] = T866[32] | 1'b0;
  assign T856[31] = T866[31] | 1'b0;
  assign T856[30] = T866[30] | 1'b0;
  assign T856[29] = T866[29] | 1'b0;
  assign T856[28] = T866[28] | 1'b0;
  assign T856[27] = T866[27] | 1'b0;
  assign T856[26] = T866[26] | 1'b0;
  assign T856[25] = T866[25] | 1'b0;
  assign T856[24] = T866[24] | 1'b0;
  assign T856[23] = T866[23] | 1'b0;
  assign T856[22] = T866[22] | 1'b0;
  assign T856[21] = T866[21] | 1'b0;
  assign T856[20] = T866[20] | 1'b0;
  assign T856[19] = T866[19] | 1'b0;
  assign T856[18] = T866[18] | 1'b0;
  assign T856[17] = T866[17] | 1'b0;
  assign T856[16] = T866[16] | 1'b0;
  assign T856[15] = T866[15] | 1'b0;
  assign T856[14] = T866[14] | 1'b0;
  assign T856[13] = T866[13] | 1'b0;
  assign T856[12] = T866[12] | 1'b0;
  assign T856[11] = T866[11] | 1'b0;
  assign T856[10] = T866[10] | 1'b0;
  assign T856[9] = T866[9] | 1'b0;
  assign T856[8] = T866[8] | 1'b0;
  assign T856[7] = T866[7] | T1013[7];
  assign T856[6] = T866[6] | T1013[6];
  assign T856[5] = T866[5] | T1013[5];
  assign T856[4] = T866[4] | T1013[4];
  assign T856[3] = T866[3] | T1013[3];
  assign T856[2] = T866[2] | T1013[2];
  assign T856[1] = T866[1] | T1013[1];
  assign T856[0] = T866[0] | T1013[0];
  assign T866[63] = T869[63] | 1'b0;
  assign T866[62] = T869[62] | 1'b0;
  assign T866[61] = T869[61] | 1'b0;
  assign T866[60] = T869[60] | 1'b0;
  assign T866[59] = T869[59] | 1'b0;
  assign T866[58] = T869[58] | 1'b0;
  assign T866[57] = T869[57] | 1'b0;
  assign T866[56] = T869[56] | 1'b0;
  assign T866[55] = T869[55] | 1'b0;
  assign T866[54] = T869[54] | 1'b0;
  assign T866[53] = T869[53] | 1'b0;
  assign T866[52] = T869[52] | 1'b0;
  assign T866[51] = T869[51] | 1'b0;
  assign T866[50] = T869[50] | 1'b0;
  assign T866[49] = T869[49] | 1'b0;
  assign T866[48] = T869[48] | 1'b0;
  assign T866[47] = T869[47] | 1'b0;
  assign T866[46] = T869[46] | 1'b0;
  assign T866[45] = T869[45] | 1'b0;
  assign T866[44] = T869[44] | 1'b0;
  assign T866[43] = T869[43] | 1'b0;
  assign T866[42] = T869[42] | 1'b0;
  assign T866[41] = T869[41] | 1'b0;
  assign T866[40] = T869[40] | 1'b0;
  assign T866[39] = T869[39] | 1'b0;
  assign T866[38] = T869[38] | 1'b0;
  assign T866[37] = T869[37] | 1'b0;
  assign T866[36] = T869[36] | 1'b0;
  assign T866[35] = T869[35] | 1'b0;
  assign T866[34] = T869[34] | 1'b0;
  assign T866[33] = T869[33] | 1'b0;
  assign T866[32] = T869[32] | 1'b0;
  assign T866[31] = T869[31] | 1'b0;
  assign T866[30] = T869[30] | T1018[30];
  assign T866[29] = T869[29] | 1'b0;
  assign T866[28] = T869[28] | 1'b0;
  assign T866[27] = T869[27] | 1'b0;
  assign T866[26] = T869[26] | 1'b0;
  assign T866[25] = T869[25] | 1'b0;
  assign T866[24] = T869[24] | 1'b0;
  assign T866[23] = T869[23] | 1'b0;
  assign T866[22] = T869[22] | 1'b0;
  assign T866[21] = T869[21] | 1'b0;
  assign T866[20] = T869[20] | 1'b0;
  assign T866[19] = T869[19] | 1'b0;
  assign T866[18] = T869[18] | 1'b0;
  assign T866[17] = T869[17] | 1'b0;
  assign T866[16] = T869[16] | 1'b0;
  assign T866[15] = T869[15] | 1'b0;
  assign T866[14] = T869[14] | 1'b0;
  assign T866[13] = T869[13] | 1'b0;
  assign T866[12] = T869[12] | 1'b0;
  assign T866[11] = T869[11] | 1'b0;
  assign T866[10] = T869[10] | 1'b0;
  assign T866[9] = T869[9] | 1'b0;
  assign T866[8] = T869[8] | 1'b0;
  assign T866[7] = T869[7] | 1'b0;
  assign T866[6] = T869[6] | 1'b0;
  assign T866[5] = T869[5] | 1'b0;
  assign T866[4] = T869[4] | 1'b0;
  assign T866[3] = T869[3] | 1'b0;
  assign T866[2] = T869[2] | 1'b0;
  assign T866[1] = T869[1] | 1'b0;
  assign T866[0] = T869[0] | 1'b0;
  assign T1018[30] = N2905;
  assign T869[63] = T871[63] | T870[63];
  assign T869[62] = T871[62] | T870[62];
  assign T869[61] = T871[61] | T870[61];
  assign T869[60] = T871[60] | T870[60];
  assign T869[59] = T871[59] | T870[59];
  assign T869[58] = T871[58] | T870[58];
  assign T869[57] = T871[57] | T870[57];
  assign T869[56] = T871[56] | T870[56];
  assign T869[55] = T871[55] | T870[55];
  assign T869[54] = T871[54] | T870[54];
  assign T869[53] = T871[53] | T870[53];
  assign T869[52] = T871[52] | T870[52];
  assign T869[51] = T871[51] | T870[51];
  assign T869[50] = T871[50] | T870[50];
  assign T869[49] = T871[49] | T870[49];
  assign T869[48] = T871[48] | T870[48];
  assign T869[47] = T871[47] | T870[47];
  assign T869[46] = T871[46] | T870[46];
  assign T869[45] = T871[45] | T870[45];
  assign T869[44] = T871[44] | T870[44];
  assign T869[43] = T871[43] | T870[43];
  assign T869[42] = T871[42] | T870[42];
  assign T869[41] = T871[41] | T870[41];
  assign T869[40] = T871[40] | T870[40];
  assign T869[39] = T871[39] | T870[39];
  assign T869[38] = T871[38] | T870[38];
  assign T869[37] = T871[37] | T870[37];
  assign T869[36] = T871[36] | T870[36];
  assign T869[35] = T871[35] | T870[35];
  assign T869[34] = T871[34] | T870[34];
  assign T869[33] = T871[33] | T870[33];
  assign T869[32] = T871[32] | T870[32];
  assign T869[31] = T871[31] | T870[31];
  assign T869[30] = T871[30] | T870[30];
  assign T869[29] = T871[29] | T870[29];
  assign T869[28] = T871[28] | T870[28];
  assign T869[27] = T871[27] | T870[27];
  assign T869[26] = T871[26] | T870[26];
  assign T869[25] = T871[25] | T870[25];
  assign T869[24] = T871[24] | T870[24];
  assign T869[23] = T871[23] | T870[23];
  assign T869[22] = T871[22] | T870[22];
  assign T869[21] = T871[21] | T870[21];
  assign T869[20] = T871[20] | T870[20];
  assign T869[19] = T871[19] | T870[19];
  assign T869[18] = T871[18] | T870[18];
  assign T869[17] = T871[17] | T870[17];
  assign T869[16] = T871[16] | T870[16];
  assign T869[15] = T871[15] | T870[15];
  assign T869[14] = T871[14] | T870[14];
  assign T869[13] = T871[13] | T870[13];
  assign T869[12] = T871[12] | T870[12];
  assign T869[11] = T871[11] | T870[11];
  assign T869[10] = T871[10] | T870[10];
  assign T869[9] = T871[9] | T870[9];
  assign T869[8] = T871[8] | T870[8];
  assign T869[7] = T871[7] | T870[7];
  assign T869[6] = T871[6] | T870[6];
  assign T869[5] = T871[5] | T870[5];
  assign T869[4] = T871[4] | T870[4];
  assign T869[3] = T871[3] | T870[3];
  assign T869[2] = T871[2] | T870[2];
  assign T869[1] = T871[1] | T870[1];
  assign T869[0] = T871[0] | T870[0];
  assign T871[63] = T875[63] | T874[63];
  assign T871[62] = T875[62] | T874[62];
  assign T871[61] = T875[61] | T874[61];
  assign T871[60] = T875[60] | T874[60];
  assign T871[59] = T875[59] | T874[59];
  assign T871[58] = T875[58] | T874[58];
  assign T871[57] = T875[57] | T874[57];
  assign T871[56] = T875[56] | T874[56];
  assign T871[55] = T875[55] | T874[55];
  assign T871[54] = T875[54] | T874[54];
  assign T871[53] = T875[53] | T874[53];
  assign T871[52] = T875[52] | T874[52];
  assign T871[51] = T875[51] | T874[51];
  assign T871[50] = T875[50] | T874[50];
  assign T871[49] = T875[49] | T874[49];
  assign T871[48] = T875[48] | T874[48];
  assign T871[47] = T875[47] | T874[47];
  assign T871[46] = T875[46] | T874[46];
  assign T871[45] = T875[45] | T874[45];
  assign T871[44] = T875[44] | T874[44];
  assign T871[43] = T875[43] | T874[43];
  assign T871[42] = T875[42] | T874[42];
  assign T871[41] = T875[41] | T874[41];
  assign T871[40] = T875[40] | T874[40];
  assign T871[39] = T875[39] | T874[39];
  assign T871[38] = T875[38] | T874[38];
  assign T871[37] = T875[37] | T874[37];
  assign T871[36] = T875[36] | T874[36];
  assign T871[35] = T875[35] | T874[35];
  assign T871[34] = T875[34] | T874[34];
  assign T871[33] = T875[33] | T874[33];
  assign T871[32] = T875[32] | T874[32];
  assign T871[31] = T875[31] | T874[31];
  assign T871[30] = T875[30] | T874[30];
  assign T871[29] = T875[29] | T874[29];
  assign T871[28] = T875[28] | T874[28];
  assign T871[27] = T875[27] | T874[27];
  assign T871[26] = T875[26] | T874[26];
  assign T871[25] = T875[25] | T874[25];
  assign T871[24] = T875[24] | T874[24];
  assign T871[23] = T875[23] | T874[23];
  assign T871[22] = T875[22] | T874[22];
  assign T871[21] = T875[21] | T874[21];
  assign T871[20] = T875[20] | T874[20];
  assign T871[19] = T875[19] | T874[19];
  assign T871[18] = T875[18] | T874[18];
  assign T871[17] = T875[17] | T874[17];
  assign T871[16] = T875[16] | T874[16];
  assign T871[15] = T875[15] | T874[15];
  assign T871[14] = T875[14] | T874[14];
  assign T871[13] = T875[13] | T874[13];
  assign T871[12] = T875[12] | T874[12];
  assign T871[11] = T875[11] | T874[11];
  assign T871[10] = T875[10] | T874[10];
  assign T871[9] = T875[9] | T874[9];
  assign T871[8] = T875[8] | T874[8];
  assign T871[7] = T875[7] | T874[7];
  assign T871[6] = T875[6] | T874[6];
  assign T871[5] = T875[5] | T874[5];
  assign T871[4] = T875[4] | T874[4];
  assign T871[3] = T875[3] | T874[3];
  assign T871[2] = T875[2] | T874[2];
  assign T871[1] = T875[1] | T874[1];
  assign T871[0] = T875[0] | T874[0];
  assign T875[63] = T876[63] | 1'b0;
  assign T875[62] = T876[62] | 1'b0;
  assign T875[61] = T876[61] | 1'b0;
  assign T875[60] = T876[60] | 1'b0;
  assign T875[59] = T876[59] | 1'b0;
  assign T875[58] = T876[58] | 1'b0;
  assign T875[57] = T876[57] | 1'b0;
  assign T875[56] = T876[56] | 1'b0;
  assign T875[55] = T876[55] | 1'b0;
  assign T875[54] = T876[54] | 1'b0;
  assign T875[53] = T876[53] | 1'b0;
  assign T875[52] = T876[52] | 1'b0;
  assign T875[51] = T876[51] | 1'b0;
  assign T875[50] = T876[50] | 1'b0;
  assign T875[49] = T876[49] | 1'b0;
  assign T875[48] = T876[48] | 1'b0;
  assign T875[47] = T876[47] | 1'b0;
  assign T875[46] = T876[46] | 1'b0;
  assign T875[45] = T876[45] | 1'b0;
  assign T875[44] = T876[44] | 1'b0;
  assign T875[43] = T876[43] | 1'b0;
  assign T875[42] = T876[42] | 1'b0;
  assign T875[41] = T876[41] | 1'b0;
  assign T875[40] = T876[40] | 1'b0;
  assign T875[39] = T876[39] | 1'b0;
  assign T875[38] = T876[38] | 1'b0;
  assign T875[37] = T876[37] | 1'b0;
  assign T875[36] = T876[36] | 1'b0;
  assign T875[35] = T876[35] | 1'b0;
  assign T875[34] = T876[34] | 1'b0;
  assign T875[33] = T876[33] | 1'b0;
  assign T875[32] = T876[32] | 1'b0;
  assign T875[31] = T876[31] | 1'b0;
  assign T875[30] = T876[30] | 1'b0;
  assign T875[29] = T876[29] | 1'b0;
  assign T875[28] = T876[28] | 1'b0;
  assign T875[27] = T876[27] | 1'b0;
  assign T875[26] = T876[26] | 1'b0;
  assign T875[25] = T876[25] | 1'b0;
  assign T875[24] = T876[24] | 1'b0;
  assign T875[23] = T876[23] | 1'b0;
  assign T875[22] = T876[22] | 1'b0;
  assign T875[21] = T876[21] | 1'b0;
  assign T875[20] = T876[20] | 1'b0;
  assign T875[19] = T876[19] | 1'b0;
  assign T875[18] = T876[18] | 1'b0;
  assign T875[17] = T876[17] | 1'b0;
  assign T875[16] = T876[16] | 1'b0;
  assign T875[15] = T876[15] | 1'b0;
  assign T875[14] = T876[14] | 1'b0;
  assign T875[13] = T876[13] | 1'b0;
  assign T875[12] = T876[12] | 1'b0;
  assign T875[11] = T876[11] | 1'b0;
  assign T875[10] = T876[10] | 1'b0;
  assign T875[9] = T876[9] | 1'b0;
  assign T875[8] = T876[8] | 1'b0;
  assign T875[7] = T876[7] | 1'b0;
  assign T875[6] = T876[6] | 1'b0;
  assign T875[5] = T876[5] | 1'b0;
  assign T875[4] = T876[4] | 1'b0;
  assign T875[3] = T876[3] | 1'b0;
  assign T875[2] = T876[2] | 1'b0;
  assign T875[1] = T876[1] | 1'b0;
  assign T875[0] = T876[0] | N2965;
  assign T876[63] = T878[63] | T877[63];
  assign T876[62] = T878[62] | 1'b0;
  assign T876[61] = T878[61] | 1'b0;
  assign T876[60] = T878[60] | 1'b0;
  assign T876[59] = T878[59] | 1'b0;
  assign T876[58] = T878[58] | 1'b0;
  assign T876[57] = T878[57] | 1'b0;
  assign T876[56] = T878[56] | 1'b0;
  assign T876[55] = T878[55] | 1'b0;
  assign T876[54] = T878[54] | 1'b0;
  assign T876[53] = T878[53] | 1'b0;
  assign T876[52] = T878[52] | 1'b0;
  assign T876[51] = T878[51] | 1'b0;
  assign T876[50] = T878[50] | 1'b0;
  assign T876[49] = T878[49] | 1'b0;
  assign T876[48] = T878[48] | 1'b0;
  assign T876[47] = T878[47] | 1'b0;
  assign T876[46] = T878[46] | 1'b0;
  assign T876[45] = T878[45] | 1'b0;
  assign T876[44] = T878[44] | 1'b0;
  assign T876[43] = T878[43] | 1'b0;
  assign T876[42] = T878[42] | 1'b0;
  assign T876[41] = T878[41] | 1'b0;
  assign T876[40] = T878[40] | 1'b0;
  assign T876[39] = T878[39] | 1'b0;
  assign T876[38] = T878[38] | 1'b0;
  assign T876[37] = T878[37] | 1'b0;
  assign T876[36] = T878[36] | 1'b0;
  assign T876[35] = T878[35] | 1'b0;
  assign T876[34] = T878[34] | 1'b0;
  assign T876[33] = T878[33] | 1'b0;
  assign T876[32] = T878[32] | 1'b0;
  assign T876[31] = T878[31] | 1'b0;
  assign T876[30] = T878[30] | 1'b0;
  assign T876[29] = T878[29] | 1'b0;
  assign T876[28] = T878[28] | 1'b0;
  assign T876[27] = T878[27] | 1'b0;
  assign T876[26] = T878[26] | 1'b0;
  assign T876[25] = T878[25] | 1'b0;
  assign T876[24] = T878[24] | 1'b0;
  assign T876[23] = T878[23] | T877[63];
  assign T876[22] = T878[22] | 1'b0;
  assign T876[21] = T878[21] | 1'b0;
  assign T876[20] = T878[20] | 1'b0;
  assign T876[19] = T878[19] | 1'b0;
  assign T876[18] = T878[18] | T877[63];
  assign T876[17] = T878[17] | 1'b0;
  assign T876[16] = T878[16] | 1'b0;
  assign T876[15] = T878[15] | 1'b0;
  assign T876[14] = T878[14] | 1'b0;
  assign T876[13] = T878[13] | 1'b0;
  assign T876[12] = T878[12] | T877[63];
  assign T876[11] = T878[11] | 1'b0;
  assign T876[10] = T878[10] | 1'b0;
  assign T876[9] = T878[9] | 1'b0;
  assign T876[8] = T878[8] | T877[63];
  assign T876[7] = T878[7] | 1'b0;
  assign T876[6] = T878[6] | 1'b0;
  assign T876[5] = T878[5] | T877[63];
  assign T876[4] = T878[4] | 1'b0;
  assign T876[3] = T878[3] | T877[63];
  assign T876[2] = T878[2] | 1'b0;
  assign T876[1] = T878[1] | 1'b0;
  assign T876[0] = T878[0] | T877[63];
  assign T877[63] = N2977;
  assign T878[63] = T880[63] | T879[63];
  assign T878[62] = T880[62] | T879[62];
  assign T878[61] = T880[61] | T879[61];
  assign T878[60] = T880[60] | T879[60];
  assign T878[59] = T880[59] | T879[59];
  assign T878[58] = T880[58] | T879[58];
  assign T878[57] = T880[57] | T879[57];
  assign T878[56] = T880[56] | T879[56];
  assign T878[55] = T880[55] | T879[55];
  assign T878[54] = T880[54] | T879[54];
  assign T878[53] = T880[53] | T879[53];
  assign T878[52] = T880[52] | T879[52];
  assign T878[51] = T880[51] | T879[51];
  assign T878[50] = T880[50] | T879[50];
  assign T878[49] = T880[49] | T879[49];
  assign T878[48] = T880[48] | T879[48];
  assign T878[47] = T880[47] | T879[47];
  assign T878[46] = T880[46] | T879[46];
  assign T878[45] = T880[45] | T879[45];
  assign T878[44] = T880[44] | T879[44];
  assign T878[43] = T880[43] | T879[43];
  assign T878[42] = T880[42] | T879[42];
  assign T878[41] = T880[41] | T879[41];
  assign T878[40] = T880[40] | T879[40];
  assign T878[39] = T880[39] | T879[39];
  assign T878[38] = T880[38] | T879[38];
  assign T878[37] = T880[37] | T879[37];
  assign T878[36] = T880[36] | T879[36];
  assign T878[35] = T880[35] | T879[35];
  assign T878[34] = T880[34] | T879[34];
  assign T878[33] = T880[33] | T879[33];
  assign T878[32] = T880[32] | T879[32];
  assign T878[31] = T880[31] | T879[31];
  assign T878[30] = T880[30] | T879[30];
  assign T878[29] = T880[29] | T879[29];
  assign T878[28] = T880[28] | T879[28];
  assign T878[27] = T880[27] | T879[27];
  assign T878[26] = T880[26] | T879[26];
  assign T878[25] = T880[25] | T879[25];
  assign T878[24] = T880[24] | T879[24];
  assign T878[23] = T880[23] | T879[23];
  assign T878[22] = T880[22] | T879[22];
  assign T878[21] = T880[21] | T879[21];
  assign T878[20] = T880[20] | T879[20];
  assign T878[19] = T880[19] | T879[19];
  assign T878[18] = T880[18] | T879[18];
  assign T878[17] = T880[17] | T879[17];
  assign T878[16] = T880[16] | T879[16];
  assign T878[15] = T880[15] | T879[15];
  assign T878[14] = T880[14] | T879[14];
  assign T878[13] = T880[13] | T879[13];
  assign T878[12] = T880[12] | T879[12];
  assign T878[11] = T880[11] | T879[11];
  assign T878[10] = T880[10] | T879[10];
  assign T878[9] = T880[9] | T879[9];
  assign T878[8] = T880[8] | T879[8];
  assign T878[7] = T880[7] | T879[7];
  assign T878[6] = T880[6] | T879[6];
  assign T878[5] = T880[5] | T879[5];
  assign T878[4] = T880[4] | T879[4];
  assign T878[3] = T880[3] | T879[3];
  assign T878[2] = T880[2] | T879[2];
  assign T878[1] = T880[1] | T879[1];
  assign T878[0] = T880[0] | T879[0];
  assign T880[63] = T882[63] | T881[63];
  assign T880[62] = T882[62] | T881[62];
  assign T880[61] = T882[61] | T881[61];
  assign T880[60] = T882[60] | T881[60];
  assign T880[59] = T882[59] | T881[59];
  assign T880[58] = T882[58] | T881[58];
  assign T880[57] = T882[57] | T881[57];
  assign T880[56] = T882[56] | T881[56];
  assign T880[55] = T882[55] | T881[55];
  assign T880[54] = T882[54] | T881[54];
  assign T880[53] = T882[53] | T881[53];
  assign T880[52] = T882[52] | T881[52];
  assign T880[51] = T882[51] | T881[51];
  assign T880[50] = T882[50] | T881[50];
  assign T880[49] = T882[49] | T881[49];
  assign T880[48] = T882[48] | T881[48];
  assign T880[47] = T882[47] | T881[47];
  assign T880[46] = T882[46] | T881[46];
  assign T880[45] = T882[45] | T881[45];
  assign T880[44] = T882[44] | T881[44];
  assign T880[43] = T882[43] | T881[43];
  assign T880[42] = T882[42] | T881[42];
  assign T880[41] = T882[41] | T881[41];
  assign T880[40] = T882[40] | T881[40];
  assign T880[39] = T882[39] | T881[39];
  assign T880[38] = T882[38] | T881[38];
  assign T880[37] = T882[37] | T881[37];
  assign T880[36] = T882[36] | T881[36];
  assign T880[35] = T882[35] | T881[35];
  assign T880[34] = T882[34] | T881[34];
  assign T880[33] = T882[33] | T881[33];
  assign T880[32] = T882[32] | T881[32];
  assign T880[31] = T882[31] | T881[31];
  assign T880[30] = T882[30] | T881[30];
  assign T880[29] = T882[29] | T881[29];
  assign T880[28] = T882[28] | T881[28];
  assign T880[27] = T882[27] | T881[27];
  assign T880[26] = T882[26] | T881[26];
  assign T880[25] = T882[25] | T881[25];
  assign T880[24] = T882[24] | T881[24];
  assign T880[23] = T882[23] | T881[23];
  assign T880[22] = T882[22] | T881[22];
  assign T880[21] = T882[21] | T881[21];
  assign T880[20] = T882[20] | T881[20];
  assign T880[19] = T882[19] | T881[19];
  assign T880[18] = T882[18] | T881[18];
  assign T880[17] = T882[17] | T881[17];
  assign T880[16] = T882[16] | T881[16];
  assign T880[15] = T882[15] | T881[15];
  assign T880[14] = T882[14] | T881[14];
  assign T880[13] = T882[13] | T881[13];
  assign T880[12] = T882[12] | T881[12];
  assign T880[11] = T882[11] | T881[11];
  assign T880[10] = T882[10] | T881[10];
  assign T880[9] = T882[9] | T881[9];
  assign T880[8] = T882[8] | T881[8];
  assign T880[7] = T882[7] | T881[7];
  assign T880[6] = T882[6] | T881[6];
  assign T880[5] = T882[5] | T881[5];
  assign T880[4] = T882[4] | T881[4];
  assign T880[3] = T882[3] | T881[3];
  assign T880[2] = T882[2] | T881[2];
  assign T880[1] = T882[1] | T881[1];
  assign T880[0] = T882[0] | T881[0];
  assign T882[63] = T884[63] | T883[63];
  assign T882[62] = T884[62] | T883[62];
  assign T882[61] = T884[61] | T883[61];
  assign T882[60] = T884[60] | T883[60];
  assign T882[59] = T884[59] | T883[59];
  assign T882[58] = T884[58] | T883[58];
  assign T882[57] = T884[57] | T883[57];
  assign T882[56] = T884[56] | T883[56];
  assign T882[55] = T884[55] | T883[55];
  assign T882[54] = T884[54] | T883[54];
  assign T882[53] = T884[53] | T883[53];
  assign T882[52] = T884[52] | T883[52];
  assign T882[51] = T884[51] | T883[51];
  assign T882[50] = T884[50] | T883[50];
  assign T882[49] = T884[49] | T883[49];
  assign T882[48] = T884[48] | T883[48];
  assign T882[47] = T884[47] | T883[47];
  assign T882[46] = T884[46] | T883[46];
  assign T882[45] = T884[45] | T883[45];
  assign T882[44] = T884[44] | T883[44];
  assign T882[43] = T884[43] | T883[43];
  assign T882[42] = T884[42] | T883[42];
  assign T882[41] = T884[41] | T883[41];
  assign T882[40] = T884[40] | T883[40];
  assign T882[39] = T884[39] | T883[39];
  assign T882[38] = T884[38] | T883[38];
  assign T882[37] = T884[37] | T883[37];
  assign T882[36] = T884[36] | T883[36];
  assign T882[35] = T884[35] | T883[35];
  assign T882[34] = T884[34] | T883[34];
  assign T882[33] = T884[33] | T883[33];
  assign T882[32] = T884[32] | T883[32];
  assign T882[31] = T884[31] | T883[31];
  assign T882[30] = T884[30] | T883[30];
  assign T882[29] = T884[29] | T883[29];
  assign T882[28] = T884[28] | T883[28];
  assign T882[27] = T884[27] | T883[27];
  assign T882[26] = T884[26] | T883[26];
  assign T882[25] = T884[25] | T883[25];
  assign T882[24] = T884[24] | T883[24];
  assign T882[23] = T884[23] | T883[23];
  assign T882[22] = T884[22] | T883[22];
  assign T882[21] = T884[21] | T883[21];
  assign T882[20] = T884[20] | T883[20];
  assign T882[19] = T884[19] | T883[19];
  assign T882[18] = T884[18] | T883[18];
  assign T882[17] = T884[17] | T883[17];
  assign T882[16] = T884[16] | T883[16];
  assign T882[15] = T884[15] | T883[15];
  assign T882[14] = T884[14] | T883[14];
  assign T882[13] = T884[13] | T883[13];
  assign T882[12] = T884[12] | T883[12];
  assign T882[11] = T884[11] | T883[11];
  assign T882[10] = T884[10] | T883[10];
  assign T882[9] = T884[9] | T883[9];
  assign T882[8] = T884[8] | T883[8];
  assign T882[7] = T884[7] | T883[7];
  assign T882[6] = T884[6] | T883[6];
  assign T882[5] = T884[5] | T883[5];
  assign T882[4] = T884[4] | T883[4];
  assign T882[3] = T884[3] | T883[3];
  assign T882[2] = T884[2] | T883[2];
  assign T882[1] = T884[1] | T883[1];
  assign T882[0] = T884[0] | T883[0];
  assign T884[63] = T886[63] | T885[63];
  assign T884[62] = T886[62] | T885[62];
  assign T884[61] = T886[61] | T885[61];
  assign T884[60] = T886[60] | T885[60];
  assign T884[59] = T886[59] | T885[59];
  assign T884[58] = T886[58] | T885[58];
  assign T884[57] = T886[57] | T885[57];
  assign T884[56] = T886[56] | T885[56];
  assign T884[55] = T886[55] | T885[55];
  assign T884[54] = T886[54] | T885[54];
  assign T884[53] = T886[53] | T885[53];
  assign T884[52] = T886[52] | T885[52];
  assign T884[51] = T886[51] | T885[51];
  assign T884[50] = T886[50] | T885[50];
  assign T884[49] = T886[49] | T885[49];
  assign T884[48] = T886[48] | T885[48];
  assign T884[47] = T886[47] | T885[47];
  assign T884[46] = T886[46] | T885[46];
  assign T884[45] = T886[45] | T885[45];
  assign T884[44] = T886[44] | T885[44];
  assign T884[43] = T886[43] | T885[43];
  assign T884[42] = T886[42] | T885[42];
  assign T884[41] = T886[41] | T885[41];
  assign T884[40] = T886[40] | T885[40];
  assign T884[39] = T886[39] | T885[39];
  assign T884[38] = T886[38] | T885[38];
  assign T884[37] = T886[37] | T885[37];
  assign T884[36] = T886[36] | T885[36];
  assign T884[35] = T886[35] | T885[35];
  assign T884[34] = T886[34] | T885[34];
  assign T884[33] = T886[33] | T885[33];
  assign T884[32] = T886[32] | T885[32];
  assign T884[31] = T886[31] | T885[31];
  assign T884[30] = T886[30] | T885[30];
  assign T884[29] = T886[29] | T885[29];
  assign T884[28] = T886[28] | T885[28];
  assign T884[27] = T886[27] | T885[27];
  assign T884[26] = T886[26] | T885[26];
  assign T884[25] = T886[25] | T885[25];
  assign T884[24] = T886[24] | T885[24];
  assign T884[23] = T886[23] | T885[23];
  assign T884[22] = T886[22] | T885[22];
  assign T884[21] = T886[21] | T885[21];
  assign T884[20] = T886[20] | T885[20];
  assign T884[19] = T886[19] | T885[19];
  assign T884[18] = T886[18] | T885[18];
  assign T884[17] = T886[17] | T885[17];
  assign T884[16] = T886[16] | T885[16];
  assign T884[15] = T886[15] | T885[15];
  assign T884[14] = T886[14] | T885[14];
  assign T884[13] = T886[13] | T885[13];
  assign T884[12] = T886[12] | T885[12];
  assign T884[11] = T886[11] | T885[11];
  assign T884[10] = T886[10] | T885[10];
  assign T884[9] = T886[9] | T885[9];
  assign T884[8] = T886[8] | T885[8];
  assign T884[7] = T886[7] | T885[7];
  assign T884[6] = T886[6] | T885[6];
  assign T884[5] = T886[5] | T885[5];
  assign T884[4] = T886[4] | T885[4];
  assign T884[3] = T886[3] | T885[3];
  assign T884[2] = T886[2] | T885[2];
  assign T884[1] = T886[1] | T885[1];
  assign T884[0] = T886[0] | T885[0];
  assign T886[63] = T888[63] | T887[63];
  assign T886[62] = T888[62] | T887[62];
  assign T886[61] = T888[61] | T887[61];
  assign T886[60] = T888[60] | T887[60];
  assign T886[59] = T888[59] | T887[59];
  assign T886[58] = T888[58] | T887[58];
  assign T886[57] = T888[57] | T887[57];
  assign T886[56] = T888[56] | T887[56];
  assign T886[55] = T888[55] | T887[55];
  assign T886[54] = T888[54] | T887[54];
  assign T886[53] = T888[53] | T887[53];
  assign T886[52] = T888[52] | T887[52];
  assign T886[51] = T888[51] | T887[51];
  assign T886[50] = T888[50] | T887[50];
  assign T886[49] = T888[49] | T887[49];
  assign T886[48] = T888[48] | T887[48];
  assign T886[47] = T888[47] | T887[47];
  assign T886[46] = T888[46] | T887[46];
  assign T886[45] = T888[45] | T887[45];
  assign T886[44] = T888[44] | T887[44];
  assign T886[43] = T888[43] | T887[43];
  assign T886[42] = T888[42] | T887[42];
  assign T886[41] = T888[41] | T887[41];
  assign T886[40] = T888[40] | T887[40];
  assign T886[39] = T888[39] | T887[39];
  assign T886[38] = T888[38] | T887[38];
  assign T886[37] = T888[37] | T887[37];
  assign T886[36] = T888[36] | T887[36];
  assign T886[35] = T888[35] | T887[35];
  assign T886[34] = T888[34] | T887[34];
  assign T886[33] = T888[33] | T887[33];
  assign T886[32] = T888[32] | T887[32];
  assign T886[31] = T888[31] | T887[31];
  assign T886[30] = T888[30] | T887[30];
  assign T886[29] = T888[29] | T887[29];
  assign T886[28] = T888[28] | T887[28];
  assign T886[27] = T888[27] | T887[27];
  assign T886[26] = T888[26] | T887[26];
  assign T886[25] = T888[25] | T887[25];
  assign T886[24] = T888[24] | T887[24];
  assign T886[23] = T888[23] | T887[23];
  assign T886[22] = T888[22] | T887[22];
  assign T886[21] = T888[21] | T887[21];
  assign T886[20] = T888[20] | T887[20];
  assign T886[19] = T888[19] | T887[19];
  assign T886[18] = T888[18] | T887[18];
  assign T886[17] = T888[17] | T887[17];
  assign T886[16] = T888[16] | T887[16];
  assign T886[15] = T888[15] | T887[15];
  assign T886[14] = T888[14] | T887[14];
  assign T886[13] = T888[13] | T887[13];
  assign T886[12] = T888[12] | T887[12];
  assign T886[11] = T888[11] | T887[11];
  assign T886[10] = T888[10] | T887[10];
  assign T886[9] = T888[9] | T887[9];
  assign T886[8] = T888[8] | T887[8];
  assign T886[7] = T888[7] | T887[7];
  assign T886[6] = T888[6] | T887[6];
  assign T886[5] = T888[5] | T887[5];
  assign T886[4] = T888[4] | T887[4];
  assign T886[3] = T888[3] | T887[3];
  assign T886[2] = T888[2] | T887[2];
  assign T886[1] = T888[1] | T887[1];
  assign T886[0] = T888[0] | T887[0];
  assign T888[63] = T890[63] | T889[63];
  assign T888[62] = T890[62] | T889[62];
  assign T888[61] = T890[61] | T889[61];
  assign T888[60] = T890[60] | T889[60];
  assign T888[59] = T890[59] | T889[59];
  assign T888[58] = T890[58] | T889[58];
  assign T888[57] = T890[57] | T889[57];
  assign T888[56] = T890[56] | T889[56];
  assign T888[55] = T890[55] | T889[55];
  assign T888[54] = T890[54] | T889[54];
  assign T888[53] = T890[53] | T889[53];
  assign T888[52] = T890[52] | T889[52];
  assign T888[51] = T890[51] | T889[51];
  assign T888[50] = T890[50] | T889[50];
  assign T888[49] = T890[49] | T889[49];
  assign T888[48] = T890[48] | T889[48];
  assign T888[47] = T890[47] | T889[47];
  assign T888[46] = T890[46] | T889[46];
  assign T888[45] = T890[45] | T889[45];
  assign T888[44] = T890[44] | T889[44];
  assign T888[43] = T890[43] | T889[43];
  assign T888[42] = T890[42] | T889[42];
  assign T888[41] = T890[41] | T889[41];
  assign T888[40] = T890[40] | T889[40];
  assign T888[39] = T890[39] | T889[39];
  assign T888[38] = T890[38] | T889[38];
  assign T888[37] = T890[37] | T889[37];
  assign T888[36] = T890[36] | T889[36];
  assign T888[35] = T890[35] | T889[35];
  assign T888[34] = T890[34] | T889[34];
  assign T888[33] = T890[33] | T889[33];
  assign T888[32] = T890[32] | T889[32];
  assign T888[31] = T890[31] | T889[31];
  assign T888[30] = T890[30] | T889[30];
  assign T888[29] = T890[29] | T889[29];
  assign T888[28] = T890[28] | T889[28];
  assign T888[27] = T890[27] | T889[27];
  assign T888[26] = T890[26] | T889[26];
  assign T888[25] = T890[25] | T889[25];
  assign T888[24] = T890[24] | T889[24];
  assign T888[23] = T890[23] | T889[23];
  assign T888[22] = T890[22] | T889[22];
  assign T888[21] = T890[21] | T889[21];
  assign T888[20] = T890[20] | T889[20];
  assign T888[19] = T890[19] | T889[19];
  assign T888[18] = T890[18] | T889[18];
  assign T888[17] = T890[17] | T889[17];
  assign T888[16] = T890[16] | T889[16];
  assign T888[15] = T890[15] | T889[15];
  assign T888[14] = T890[14] | T889[14];
  assign T888[13] = T890[13] | T889[13];
  assign T888[12] = T890[12] | T889[12];
  assign T888[11] = T890[11] | T889[11];
  assign T888[10] = T890[10] | T889[10];
  assign T888[9] = T890[9] | T889[9];
  assign T888[8] = T890[8] | T889[8];
  assign T888[7] = T890[7] | T889[7];
  assign T888[6] = T890[6] | T889[6];
  assign T888[5] = T890[5] | T889[5];
  assign T888[4] = T890[4] | T889[4];
  assign T888[3] = T890[3] | T889[3];
  assign T888[2] = T890[2] | T889[2];
  assign T888[1] = T890[1] | T889[1];
  assign T888[0] = T890[0] | T889[0];
  assign T890[63] = 1'b0 | T891[63];
  assign T890[62] = 1'b0 | T891[62];
  assign T890[61] = 1'b0 | T891[61];
  assign T890[60] = 1'b0 | T891[60];
  assign T890[59] = 1'b0 | T891[59];
  assign T890[58] = 1'b0 | T891[58];
  assign T890[57] = 1'b0 | T891[57];
  assign T890[56] = 1'b0 | T891[56];
  assign T890[55] = 1'b0 | T891[55];
  assign T890[54] = 1'b0 | T891[54];
  assign T890[53] = 1'b0 | T891[53];
  assign T890[52] = 1'b0 | T891[52];
  assign T890[51] = 1'b0 | T891[51];
  assign T890[50] = 1'b0 | T891[50];
  assign T890[49] = 1'b0 | T891[49];
  assign T890[48] = 1'b0 | T891[48];
  assign T890[47] = 1'b0 | T891[47];
  assign T890[46] = 1'b0 | T891[46];
  assign T890[45] = 1'b0 | T891[45];
  assign T890[44] = 1'b0 | T891[44];
  assign T890[43] = 1'b0 | T891[43];
  assign T890[42] = 1'b0 | T891[42];
  assign T890[41] = 1'b0 | T891[41];
  assign T890[40] = 1'b0 | T891[40];
  assign T890[39] = 1'b0 | T891[39];
  assign T890[38] = 1'b0 | T891[38];
  assign T890[37] = 1'b0 | T891[37];
  assign T890[36] = 1'b0 | T891[36];
  assign T890[35] = 1'b0 | T891[35];
  assign T890[34] = 1'b0 | T891[34];
  assign T890[33] = 1'b0 | T891[33];
  assign T890[32] = 1'b0 | T891[32];
  assign T890[31] = 1'b0 | T891[31];
  assign T890[30] = 1'b0 | T891[30];
  assign T890[29] = 1'b0 | T891[29];
  assign T890[28] = 1'b0 | T891[28];
  assign T890[27] = 1'b0 | T891[27];
  assign T890[26] = 1'b0 | T891[26];
  assign T890[25] = 1'b0 | T891[25];
  assign T890[24] = 1'b0 | T891[24];
  assign T890[23] = 1'b0 | T891[23];
  assign T890[22] = 1'b0 | T891[22];
  assign T890[21] = 1'b0 | T891[21];
  assign T890[20] = 1'b0 | T891[20];
  assign T890[19] = 1'b0 | T891[19];
  assign T890[18] = 1'b0 | T891[18];
  assign T890[17] = 1'b0 | T891[17];
  assign T890[16] = 1'b0 | T891[16];
  assign T890[15] = 1'b0 | T891[15];
  assign T890[14] = 1'b0 | T891[14];
  assign T890[13] = 1'b0 | T891[13];
  assign T890[12] = 1'b0 | T891[12];
  assign T890[11] = 1'b0 | T891[11];
  assign T890[10] = 1'b0 | T891[10];
  assign T890[9] = 1'b0 | T891[9];
  assign T890[8] = 1'b0 | T891[8];
  assign T890[7] = T1020[7] | T891[7];
  assign T890[6] = T1020[6] | T891[6];
  assign T890[5] = T1020[5] | T891[5];
  assign T890[4] = T1020[4] | T891[4];
  assign T890[3] = T1020[3] | T891[3];
  assign T890[2] = T1020[2] | T891[2];
  assign T890[1] = T1020[1] | T891[1];
  assign T890[0] = T1020[0] | T891[0];
  assign T1020[7] = 1'b0 | T893[7];
  assign T1020[6] = 1'b0 | T893[6];
  assign T1020[5] = 1'b0 | T893[5];
  assign T1020[4] = T1023[4] | T893[4];
  assign T1020[3] = T1023[3] | T893[3];
  assign T1020[2] = T1023[2] | T893[2];
  assign T1020[1] = T1023[1] | T893[1];
  assign T1020[0] = T1023[0] | T893[0];
  assign N185 = ~T899;
  assign N186 = ~io_fcsr_flags_valid;
  assign T898[4] = T894[4] | io_fcsr_flags_bits[4];
  assign T898[3] = T894[3] | io_fcsr_flags_bits[3];
  assign T898[2] = T894[2] | io_fcsr_flags_bits[2];
  assign T898[1] = T894[1] | io_fcsr_flags_bits[1];
  assign T898[0] = T894[0] | io_fcsr_flags_bits[0];
  assign T899 = io_rocc_csr_wen & N3085;
  assign T1023[4] = T902[4] | 1'b0;
  assign T1023[3] = T902[3] | 1'b0;
  assign T1023[2] = T902[2] | T1024[2];
  assign T1023[1] = T902[1] | T1024[1];
  assign T1023[0] = T902[0] | T1024[0];
  assign T905 = ~io_host_csr_resp_ready;
  assign T906 = io_host_csr_resp_ready & T907;
  assign T907 = ~host_csr_req_fire;
  assign io_host_csr_req_ready = T910 & T909;
  assign T909 = ~io_host_csr_resp_valid;
  assign T910 = ~host_csr_req_valid;
  assign N187 = T88 | reset;
  assign N188 = T216[0] | N187;
  assign N189 = T914[0] | N188;
  assign N190 = T25 | N189;
  assign N191 = ~N190;
  assign N195 = T76 | reset;
  assign N196 = T69 | N195;
  assign N197 = T914[0] | N196;
  assign N198 = T25 | N197;
  assign N199 = ~N198;
  assign N203 = T52 | reset;
  assign N204 = T914[0] | N203;
  assign N205 = T25 | N204;
  assign N206 = ~N205;
  assign N210 = T40 | host_csr_req_fire;
  assign N211 = ~N210;
  assign N277 = ~host_csr_req_valid;
  assign N279 = T76 | reset;
  assign N280 = T58 | N279;
  assign N281 = T914[0] | N280;
  assign N282 = T25 | N281;
  assign N283 = ~N282;
  assign N286 = T76 | reset;
  assign N287 = T58 | N286;
  assign N288 = T914[0] | N287;
  assign N289 = T25 | N288;
  assign N290 = ~N289;
  assign N293 = T58 | reset;
  assign N294 = T914[0] | N293;
  assign N295 = T25 | N294;
  assign N296 = ~N295;
  assign N299 = T253 | reset;
  assign N300 = T251 | N299;
  assign N301 = ~N300;
  assign N304 = T259 | reset;
  assign N305 = T257 | N304;
  assign N306 = ~N305;
  assign N309 = T270 | reset;
  assign N310 = T251 | N309;
  assign N311 = ~N310;
  assign N314 = T257 | reset;
  assign N315 = ~N314;
  assign N318 = T251 | reset;
  assign N319 = ~N318;
  assign N322 = T259 | reset;
  assign N323 = T257 | N322;
  assign N324 = ~N323;
  assign N327 = T297 | reset;
  assign N328 = T293 | N327;
  assign N329 = ~N328;
  assign N332 = T257 | reset;
  assign N333 = ~N332;
  assign N336 = T307 | reset;
  assign N337 = ~N336;
  assign N403 = ~reset;
  assign N410 = T326[6] | reset;
  assign N411 = ~N410;
  assign N471 = T367 | reset;
  assign N472 = ~N471;
  assign N474 = T76 | reset;
  assign N475 = T58 | N474;
  assign N476 = ~N475;
  assign N480 = T76 | reset;
  assign N481 = T58 | N480;
  assign N482 = ~N481;
  assign N486 = T76 | reset;
  assign N487 = T58 | N486;
  assign N488 = T25 | N487;
  assign N489 = ~N488;
  assign N492 = T402 | reset;
  assign N493 = T399 | N492;
  assign N494 = ~N493;
  assign N497 = some_interrupt_pending | reset;
  assign N498 = insn_wfi | N497;
  assign N499 = ~N498;
  assign N502 = T465 | T474;
  assign N503 = T25 | N502;
  assign N504 = ~N503;
  assign N546 = T488 | T490;
  assign N547 = T486 | N546;
  assign N548 = T485 | N547;
  assign N549 = T25 | N548;
  assign N550 = ~N549;
  assign N616 = io_uarch_counters_15 | reset;
  assign N617 = ~N616;
  assign N625 = T591 | reset;
  assign N626 = ~N625;
  assign N686 = io_uarch_counters_14 | reset;
  assign N687 = ~N686;
  assign N695 = T604 | reset;
  assign N696 = ~N695;
  assign N756 = io_uarch_counters_13 | reset;
  assign N757 = ~N756;
  assign N765 = T617 | reset;
  assign N766 = ~N765;
  assign N826 = io_uarch_counters_12 | reset;
  assign N827 = ~N826;
  assign N835 = T630 | reset;
  assign N836 = ~N835;
  assign N896 = io_uarch_counters_11 | reset;
  assign N897 = ~N896;
  assign N905 = T643 | reset;
  assign N906 = ~N905;
  assign N966 = io_uarch_counters_10 | reset;
  assign N967 = ~N966;
  assign N975 = T656 | reset;
  assign N976 = ~N975;
  assign N1036 = io_uarch_counters_9 | reset;
  assign N1037 = ~N1036;
  assign N1045 = T669 | reset;
  assign N1046 = ~N1045;
  assign N1106 = io_uarch_counters_8 | reset;
  assign N1107 = ~N1106;
  assign N1115 = T682 | reset;
  assign N1116 = ~N1115;
  assign N1176 = io_uarch_counters_7 | reset;
  assign N1177 = ~N1176;
  assign N1185 = T695 | reset;
  assign N1186 = ~N1185;
  assign N1246 = io_uarch_counters_6 | reset;
  assign N1247 = ~N1246;
  assign N1255 = T708 | reset;
  assign N1256 = ~N1255;
  assign N1316 = io_uarch_counters_5 | reset;
  assign N1317 = ~N1316;
  assign N1325 = T721 | reset;
  assign N1326 = ~N1325;
  assign N1386 = io_uarch_counters_4 | reset;
  assign N1387 = ~N1386;
  assign N1395 = T734 | reset;
  assign N1396 = ~N1395;
  assign N1456 = io_uarch_counters_3 | reset;
  assign N1457 = ~N1456;
  assign N1465 = T747 | reset;
  assign N1466 = ~N1465;
  assign N1526 = io_uarch_counters_2 | reset;
  assign N1527 = ~N1526;
  assign N1535 = T760 | reset;
  assign N1536 = ~N1535;
  assign N1596 = io_uarch_counters_1 | reset;
  assign N1597 = ~N1596;
  assign N1605 = T773 | reset;
  assign N1606 = ~N1605;
  assign N1666 = io_uarch_counters_0 | reset;
  assign N1667 = ~N1666;
  assign N1675 = T786 | reset;
  assign N1676 = ~N1675;
  assign N1736 = T798 | reset;
  assign N1737 = io_retire | N1736;
  assign N1738 = ~N1737;
  assign N1746 = T798 | reset;
  assign N1747 = T803 | N1746;
  assign N1748 = ~N1747;
  assign N1808 = T817 | reset;
  assign N1809 = T814 | N1808;
  assign N1810 = ~N1809;
  assign N1876 = T825 | reset;
  assign N1877 = ~N1876;
  assign N1880 = ~io_host_csr_resp_valid;
  assign N1882 = T88 & N1901;
  assign N1883 = ~T88;
  assign N1884 = N1901 & N1883;
  assign N1885 = T216[0] & N1884;
  assign N1886 = ~T216[0];
  assign N1887 = N1884 & N1886;
  assign N1888 = T914[0] & N1887;
  assign N1889 = ~T914[0];
  assign N1890 = N1887 & N1889;
  assign N1891 = T25 & N1890;
  assign N1892 = T76 & N1901;
  assign N1893 = ~T76;
  assign N1894 = N1901 & N1893;
  assign N1895 = T69 & N1894;
  assign N1896 = ~T69;
  assign N1897 = N1894 & N1896;
  assign N1898 = T914[0] & N1897;
  assign N1899 = N1897 & N1889;
  assign N1900 = T25 & N1899;
  assign N1901 = ~reset;
  assign N1902 = T52 & N1901;
  assign N1903 = ~T52;
  assign N1904 = N1901 & N1903;
  assign N1905 = T914[0] & N1904;
  assign N1906 = N1904 & N1889;
  assign N1907 = T25 & N1906;
  assign N1908 = ~host_csr_req_fire;
  assign N1909 = T40 & N1908;
  assign N1910 = T76 & N1901;
  assign N1911 = N1901 & N1893;
  assign N1912 = T58 & N1911;
  assign N1913 = ~T58;
  assign N1914 = N1911 & N1913;
  assign N1915 = T914[0] & N1914;
  assign N1916 = N1914 & N1889;
  assign N1917 = T25 & N1916;
  assign N1918 = T76 & N1901;
  assign N1919 = N1901 & N1893;
  assign N1920 = T58 & N1919;
  assign N1921 = N1919 & N1913;
  assign N1922 = T914[0] & N1921;
  assign N1923 = N1921 & N1889;
  assign N1924 = T25 & N1923;
  assign N1925 = T58 & N1901;
  assign N1926 = N1901 & N1913;
  assign N1927 = T914[0] & N1926;
  assign N1928 = N1926 & N1889;
  assign N1929 = T25 & N1928;
  assign N1930 = T253 & N1901;
  assign N1931 = ~T253;
  assign N1932 = N1901 & N1931;
  assign N1933 = T251 & N1932;
  assign N1934 = T259 & N1901;
  assign N1935 = ~T259;
  assign N1936 = N1901 & N1935;
  assign N1937 = T257 & N1936;
  assign N1938 = T270 & N1901;
  assign N1939 = ~T270;
  assign N1940 = N1901 & N1939;
  assign N1941 = T251 & N1940;
  assign N1942 = T257 & N1901;
  assign N1943 = T251 & N1901;
  assign N1944 = T259 & N1901;
  assign N1945 = N1901 & N1935;
  assign N1946 = T257 & N1945;
  assign N1947 = T297 & N1901;
  assign N1948 = ~T297;
  assign N1949 = N1901 & N1948;
  assign N1950 = T293 & N1949;
  assign N1951 = T257 & N1901;
  assign N1952 = T307 & N1901;
  assign N1953 = T326[6] & N1901;
  assign N1954 = T367 & N1901;
  assign N1955 = T76 & N1901;
  assign N1956 = N1901 & N1893;
  assign N1957 = T58 & N1956;
  assign N1958 = T76 & N1901;
  assign N1959 = N1901 & N1893;
  assign N1960 = T58 & N1959;
  assign N1961 = T76 & N1901;
  assign N1962 = N1901 & N1893;
  assign N1963 = T58 & N1962;
  assign N1964 = N1962 & N1913;
  assign N1965 = T25 & N1964;
  assign N1966 = T402 & N1901;
  assign N1967 = ~T402;
  assign N1968 = N1901 & N1967;
  assign N1969 = T399 & N1968;
  assign N1970 = some_interrupt_pending & N1901;
  assign N1971 = ~some_interrupt_pending;
  assign N1972 = N1901 & N1971;
  assign N1973 = insn_wfi & N1972;
  assign N1974 = ~T474;
  assign N1975 = T465 & N1974;
  assign N1976 = ~T465;
  assign N1977 = N1974 & N1976;
  assign N1978 = T25 & N1977;
  assign N1979 = ~T490;
  assign N1980 = T488 & N1979;
  assign N1981 = ~T488;
  assign N1982 = N1979 & N1981;
  assign N1983 = T486 & N1982;
  assign N1984 = ~T486;
  assign N1985 = N1982 & N1984;
  assign N1986 = T485 & N1985;
  assign N1987 = ~T485;
  assign N1988 = N1985 & N1987;
  assign N1989 = T25 & N1988;
  assign N1990 = io_uarch_counters_15 & N1901;
  assign N1991 = T591 & N1901;
  assign N1992 = io_uarch_counters_14 & N1901;
  assign N1993 = T604 & N1901;
  assign N1994 = io_uarch_counters_13 & N1901;
  assign N1995 = T617 & N1901;
  assign N1996 = io_uarch_counters_12 & N1901;
  assign N1997 = T630 & N1901;
  assign N1998 = io_uarch_counters_11 & N1901;
  assign N1999 = T643 & N1901;
  assign N2000 = io_uarch_counters_10 & N1901;
  assign N2001 = T656 & N1901;
  assign N2002 = io_uarch_counters_9 & N1901;
  assign N2003 = T669 & N1901;
  assign N2004 = io_uarch_counters_8 & N1901;
  assign N2005 = T682 & N1901;
  assign N2006 = io_uarch_counters_7 & N1901;
  assign N2007 = T695 & N1901;
  assign N2008 = io_uarch_counters_6 & N1901;
  assign N2009 = T708 & N1901;
  assign N2010 = io_uarch_counters_5 & N1901;
  assign N2011 = T721 & N1901;
  assign N2012 = io_uarch_counters_4 & N1901;
  assign N2013 = T734 & N1901;
  assign N2014 = io_uarch_counters_3 & N1901;
  assign N2015 = T747 & N1901;
  assign N2016 = io_uarch_counters_2 & N1901;
  assign N2017 = T760 & N1901;
  assign N2018 = io_uarch_counters_1 & N1901;
  assign N2019 = T773 & N1901;
  assign N2020 = io_uarch_counters_0 & N1901;
  assign N2021 = T786 & N1901;
  assign N2022 = T798 & N1901;
  assign N2023 = ~T798;
  assign N2024 = N1901 & N2023;
  assign N2025 = io_retire & N2024;
  assign N2026 = T798 & N1901;
  assign N2027 = N1901 & N2023;
  assign N2028 = T803 & N2027;
  assign N2029 = T817 & N1901;
  assign N2030 = ~T817;
  assign N2031 = N1901 & N2030;
  assign N2032 = T814 & N2031;
  assign N2033 = T825 & N1901;

endmodule