module AMOALU( // @[:freechips.rocketchip.system.TinyConfig.fir@105905.2]
  input  [4:0]  io_cmd, // @[:freechips.rocketchip.system.TinyConfig.fir@105908.4]
  input  [31:0] io_lhs, // @[:freechips.rocketchip.system.TinyConfig.fir@105908.4]
  input  [31:0] io_rhs, // @[:freechips.rocketchip.system.TinyConfig.fir@105908.4]
  output [31:0] io_out_unmasked // @[:freechips.rocketchip.system.TinyConfig.fir@105908.4]
);
  wire  _T; // @[AMOALU.scala 64:20:freechips.rocketchip.system.TinyConfig.fir@105913.4]
  wire  _T_1; // @[AMOALU.scala 64:43:freechips.rocketchip.system.TinyConfig.fir@105914.4]
  wire  max; // @[AMOALU.scala 64:33:freechips.rocketchip.system.TinyConfig.fir@105915.4]
  wire  _T_2; // @[AMOALU.scala 65:20:freechips.rocketchip.system.TinyConfig.fir@105916.4]
  wire  _T_3; // @[AMOALU.scala 65:43:freechips.rocketchip.system.TinyConfig.fir@105917.4]
  wire  min; // @[AMOALU.scala 65:33:freechips.rocketchip.system.TinyConfig.fir@105918.4]
  wire  add; // @[AMOALU.scala 66:20:freechips.rocketchip.system.TinyConfig.fir@105919.4]
  wire  _T_4; // @[AMOALU.scala 67:26:freechips.rocketchip.system.TinyConfig.fir@105920.4]
  wire  _T_5; // @[AMOALU.scala 67:48:freechips.rocketchip.system.TinyConfig.fir@105921.4]
  wire  logic_and; // @[AMOALU.scala 67:38:freechips.rocketchip.system.TinyConfig.fir@105922.4]
  wire  _T_6; // @[AMOALU.scala 68:26:freechips.rocketchip.system.TinyConfig.fir@105923.4]
  wire  logic_xor; // @[AMOALU.scala 68:39:freechips.rocketchip.system.TinyConfig.fir@105925.4]
  wire [31:0] adder_out; // @[AMOALU.scala 73:21:freechips.rocketchip.system.TinyConfig.fir@105930.4]
  wire [4:0] _T_14; // @[AMOALU.scala 86:17:freechips.rocketchip.system.TinyConfig.fir@105933.4]
  wire  _T_16; // @[AMOALU.scala 86:25:freechips.rocketchip.system.TinyConfig.fir@105935.4]
  wire  _T_17; // @[AMOALU.scala 88:12:freechips.rocketchip.system.TinyConfig.fir@105936.4]
  wire  _T_18; // @[AMOALU.scala 88:23:freechips.rocketchip.system.TinyConfig.fir@105937.4]
  wire  _T_19; // @[AMOALU.scala 88:18:freechips.rocketchip.system.TinyConfig.fir@105938.4]
  wire  _T_22; // @[AMOALU.scala 79:35:freechips.rocketchip.system.TinyConfig.fir@105941.4]
  wire  _T_25; // @[AMOALU.scala 88:58:freechips.rocketchip.system.TinyConfig.fir@105944.4]
  wire  less; // @[AMOALU.scala 88:10:freechips.rocketchip.system.TinyConfig.fir@105945.4]
  wire  _T_26; // @[AMOALU.scala 94:23:freechips.rocketchip.system.TinyConfig.fir@105946.4]
  wire [31:0] minmax; // @[AMOALU.scala 94:19:freechips.rocketchip.system.TinyConfig.fir@105947.4]
  wire [31:0] _T_27; // @[AMOALU.scala 96:27:freechips.rocketchip.system.TinyConfig.fir@105948.4]
  wire [31:0] _T_28; // @[AMOALU.scala 96:8:freechips.rocketchip.system.TinyConfig.fir@105949.4]
  wire [31:0] _T_29; // @[AMOALU.scala 97:27:freechips.rocketchip.system.TinyConfig.fir@105950.4]
  wire [31:0] _T_30; // @[AMOALU.scala 97:8:freechips.rocketchip.system.TinyConfig.fir@105951.4]
  wire [31:0] logic_; // @[AMOALU.scala 96:42:freechips.rocketchip.system.TinyConfig.fir@105952.4]
  wire  _T_31; // @[AMOALU.scala 100:19:freechips.rocketchip.system.TinyConfig.fir@105953.4]
  wire [31:0] _T_32; // @[AMOALU.scala 100:8:freechips.rocketchip.system.TinyConfig.fir@105954.4]
  assign _T = io_cmd == 5'hd; // @[AMOALU.scala 64:20:freechips.rocketchip.system.TinyConfig.fir@105913.4]
  assign _T_1 = io_cmd == 5'hf; // @[AMOALU.scala 64:43:freechips.rocketchip.system.TinyConfig.fir@105914.4]
  assign max = _T | _T_1; // @[AMOALU.scala 64:33:freechips.rocketchip.system.TinyConfig.fir@105915.4]
  assign _T_2 = io_cmd == 5'hc; // @[AMOALU.scala 65:20:freechips.rocketchip.system.TinyConfig.fir@105916.4]
  assign _T_3 = io_cmd == 5'he; // @[AMOALU.scala 65:43:freechips.rocketchip.system.TinyConfig.fir@105917.4]
  assign min = _T_2 | _T_3; // @[AMOALU.scala 65:33:freechips.rocketchip.system.TinyConfig.fir@105918.4]
  assign add = io_cmd == 5'h8; // @[AMOALU.scala 66:20:freechips.rocketchip.system.TinyConfig.fir@105919.4]
  assign _T_4 = io_cmd == 5'ha; // @[AMOALU.scala 67:26:freechips.rocketchip.system.TinyConfig.fir@105920.4]
  assign _T_5 = io_cmd == 5'hb; // @[AMOALU.scala 67:48:freechips.rocketchip.system.TinyConfig.fir@105921.4]
  assign logic_and = _T_4 | _T_5; // @[AMOALU.scala 67:38:freechips.rocketchip.system.TinyConfig.fir@105922.4]
  assign _T_6 = io_cmd == 5'h9; // @[AMOALU.scala 68:26:freechips.rocketchip.system.TinyConfig.fir@105923.4]
  assign logic_xor = _T_6 | _T_4; // @[AMOALU.scala 68:39:freechips.rocketchip.system.TinyConfig.fir@105925.4]
  assign adder_out = io_lhs + io_rhs; // @[AMOALU.scala 73:21:freechips.rocketchip.system.TinyConfig.fir@105930.4]
  assign _T_14 = io_cmd & 5'h2; // @[AMOALU.scala 86:17:freechips.rocketchip.system.TinyConfig.fir@105933.4]
  assign _T_16 = _T_14 == 5'h0; // @[AMOALU.scala 86:25:freechips.rocketchip.system.TinyConfig.fir@105935.4]
  assign _T_17 = io_lhs[31]; // @[AMOALU.scala 88:12:freechips.rocketchip.system.TinyConfig.fir@105936.4]
  assign _T_18 = io_rhs[31]; // @[AMOALU.scala 88:23:freechips.rocketchip.system.TinyConfig.fir@105937.4]
  assign _T_19 = _T_17 == _T_18; // @[AMOALU.scala 88:18:freechips.rocketchip.system.TinyConfig.fir@105938.4]
  assign _T_22 = io_lhs < io_rhs; // @[AMOALU.scala 79:35:freechips.rocketchip.system.TinyConfig.fir@105941.4]
  assign _T_25 = _T_16 ? _T_17 : _T_18; // @[AMOALU.scala 88:58:freechips.rocketchip.system.TinyConfig.fir@105944.4]
  assign less = _T_19 ? _T_22 : _T_25; // @[AMOALU.scala 88:10:freechips.rocketchip.system.TinyConfig.fir@105945.4]
  assign _T_26 = less ? min : max; // @[AMOALU.scala 94:23:freechips.rocketchip.system.TinyConfig.fir@105946.4]
  assign minmax = _T_26 ? io_lhs : io_rhs; // @[AMOALU.scala 94:19:freechips.rocketchip.system.TinyConfig.fir@105947.4]
  assign _T_27 = io_lhs & io_rhs; // @[AMOALU.scala 96:27:freechips.rocketchip.system.TinyConfig.fir@105948.4]
  assign _T_28 = logic_and ? _T_27 : 32'h0; // @[AMOALU.scala 96:8:freechips.rocketchip.system.TinyConfig.fir@105949.4]
  assign _T_29 = io_lhs ^ io_rhs; // @[AMOALU.scala 97:27:freechips.rocketchip.system.TinyConfig.fir@105950.4]
  assign _T_30 = logic_xor ? _T_29 : 32'h0; // @[AMOALU.scala 97:8:freechips.rocketchip.system.TinyConfig.fir@105951.4]
  assign logic_ = _T_28 | _T_30; // @[AMOALU.scala 96:42:freechips.rocketchip.system.TinyConfig.fir@105952.4]
  assign _T_31 = logic_and | logic_xor; // @[AMOALU.scala 100:19:freechips.rocketchip.system.TinyConfig.fir@105953.4]
  assign _T_32 = _T_31 ? logic_ : minmax; // @[AMOALU.scala 100:8:freechips.rocketchip.system.TinyConfig.fir@105954.4]
  assign io_out_unmasked = add ? adder_out : _T_32; // @[AMOALU.scala 105:19:freechips.rocketchip.system.TinyConfig.fir@105976.4]
endmodule