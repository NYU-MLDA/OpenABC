module loadstore1_0_bf8b4530d8d246dd74ac53a13471bba17941dff7(clk, rst, \l_in.valid , \l_in.op , \l_in.nia , \l_in.insn , \l_in.instr_tag , \l_in.addr1 , \l_in.addr2 , \l_in.data , \l_in.write_reg , \l_in.length , \l_in.ci , \l_in.byte_reverse , \l_in.sign_extend , \l_in.update , \l_in.xerc , \l_in.reserve , \l_in.rc , \l_in.virt_mode , \l_in.priv_mode , \l_in.mode_32bit , \l_in.is_32bit , \l_in.repeat , \l_in.second , \l_in.msr , \d_in.valid , \d_in.data , \d_in.store_done , \d_in.error , \d_in.cache_paradox , \m_in.done , \m_in.err , \m_in.invalid , \m_in.badtree , \m_in.segerr , \m_in.perm_error , \m_in.rc_error , \m_in.sprval , dc_stall, \e_out.busy , \e_out.in_progress , \e_out.interrupt , \l_out.valid , \l_out.instr_tag , \l_out.write_enable , \l_out.write_reg , \l_out.write_data , \l_out.xerc , \l_out.rc , \l_out.store_done , \l_out.interrupt , \l_out.intr_vec , \l_out.srr0 , \l_out.srr1 , \d_out.valid , \d_out.hold , \d_out.load , \d_out.dcbz , \d_out.nc , \d_out.reserve , \d_out.atomic , \d_out.atomic_last , \d_out.virt_mode , \d_out.priv_mode , \d_out.addr , \d_out.data , \d_out.byte_sel , \m_out.valid , \m_out.tlbie , \m_out.slbia , \m_out.mtspr , \m_out.iside , \m_out.load , \m_out.priv , \m_out.sprn , \m_out.addr , \m_out.rs , \events.load_complete , \events.store_complete , \events.itlb_miss , log_out);
  wire [7:0] _0000_;
  wire [7:0] _0001_;
  wire [7:0] _0002_;
  wire [7:0] _0003_;
  wire [7:0] _0004_;
  wire [7:0] _0005_;
  wire [7:0] _0006_;
  wire [7:0] _0007_;
  wire [7:0] _0008_;
  wire [7:0] _0009_;
  wire [7:0] _0010_;
  wire [7:0] _0011_;
  wire [7:0] _0012_;
  wire [7:0] _0013_;
  wire [7:0] _0014_;
  wire [7:0] _0015_;
  wire [7:0] _0016_;
  wire [7:0] _0017_;
  wire [7:0] _0018_;
  wire [7:0] _0019_;
  wire [7:0] _0020_;
  wire [7:0] _0021_;
  wire [7:0] _0022_;
  wire [7:0] _0023_;
  wire [7:0] _0024_;
  wire [7:0] _0025_;
  wire [7:0] _0026_;
  wire [7:0] _0027_;
  wire [7:0] _0028_;
  wire [7:0] _0029_;
  wire [7:0] _0030_;
  wire [7:0] _0031_;
  wire [7:0] _0032_;
  wire [7:0] _0033_;
  wire [7:0] _0034_;
  wire [7:0] _0035_;
  wire [7:0] _0036_;
  wire [7:0] _0037_;
  wire [7:0] _0038_;
  wire [7:0] _0039_;
  wire [7:0] _0040_;
  wire [7:0] _0041_;
  wire [7:0] _0042_;
  wire [7:0] _0043_;
  wire [7:0] _0044_;
  wire [7:0] _0045_;
  wire [7:0] _0046_;
  wire [7:0] _0047_;
  wire [7:0] _0048_;
  wire [7:0] _0049_;
  wire [7:0] _0050_;
  wire [7:0] _0051_;
  wire [7:0] _0052_;
  wire [7:0] _0053_;
  wire [7:0] _0054_;
  wire [7:0] _0055_;
  wire [7:0] _0056_;
  wire [7:0] _0057_;
  wire [7:0] _0058_;
  wire [7:0] _0059_;
  wire [7:0] _0060_;
  wire [7:0] _0061_;
  wire [7:0] _0062_;
  wire [7:0] _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire [336:0] _0069_;
  wire _0070_;
  wire [303:0] _0071_;
  wire [2:0] _0072_;
  wire [65:0] _0073_;
  wire [1:0] _0074_;
  wire [2:0] _0075_;
  wire _0076_;
  wire [77:0] _0077_;
  wire _0078_;
  wire [63:0] _0079_;
  wire [95:0] _0080_;
  wire [38:0] _0081_;
  wire [1:0] _0082_;
  wire [94:0] _0083_;
  wire _0084_;
  reg [337:0] _0085_;
  reg [373:0] _0086_;
  reg [380:0] _0087_;
  reg _0088_;
  reg _0089_;
  wire _0090_;
  wire _0091_;
  wire [4:0] _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire [22:0] _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire [22:0] _0102_;
  wire [22:0] _0103_;
  wire [22:0] _0104_;
  wire [7:0] _0105_;
  wire _0106_;
  wire _0107_;
  wire [10:0] _0108_;
  wire _0109_;
  wire [10:0] _0110_;
  wire [4:0] _0111_;
  wire [10:0] _0112_;
  wire [4:0] _0113_;
  wire [10:0] _0114_;
  wire [4:0] _0115_;
  wire [10:0] _0116_;
  wire [4:0] _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire [22:0] _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire [22:0] _0127_;
  wire [63:0] _0128_;
  wire _0129_;
  wire [63:0] _0130_;
  wire _0131_;
  wire [60:0] _0132_;
  wire [31:0] _0133_;
  wire [31:0] _0134_;
  wire [31:0] _0135_;
  wire [31:0] _0136_;
  wire [31:0] _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire [2:0] _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire [7:0] _0147_;
  wire [15:0] _0148_;
  wire _0149_;
  wire _0150_;
  wire [2:0] _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire [63:0] _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire [2:0] _0205_;
  wire [2:0] _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire [63:0] _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire [60:0] _0243_;
  wire _0244_;
  wire [71:0] _0245_;
  wire [71:0] _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire [71:0] _0250_;
  wire [71:0] _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire [71:0] _0257_;
  wire [71:0] _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire [71:0] _0264_;
  wire [71:0] _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire [63:0] _0271_;
  wire [71:0] _0272_;
  wire [71:0] _0273_;
  wire _0274_;
  wire _0275_;
  wire [64:0] _0276_;
  wire [120:0] _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire [12:0] _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire [2:0] _0289_;
  wire [2:0] _0290_;
  wire [2:0] _0291_;
  wire [2:0] _0292_;
  wire [2:0] _0293_;
  wire [2:0] _0294_;
  wire [2:0] _0295_;
  wire [2:0] _0296_;
  wire [2:0] _0297_;
  wire [2:0] _0298_;
  wire [2:0] _0299_;
  wire [2:0] _0300_;
  wire [2:0] _0301_;
  wire [2:0] _0302_;
  wire [2:0] _0303_;
  wire [2:0] _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire [1:0] _0327_;
  wire [1:0] _0328_;
  wire [1:0] _0329_;
  wire [2:0] _0330_;
  wire [3:0] _0331_;
  wire [2:0] _0332_;
  wire [3:0] _0333_;
  wire [2:0] _0334_;
  wire [3:0] _0335_;
  wire [2:0] _0336_;
  wire [3:0] _0337_;
  wire [2:0] _0338_;
  wire [3:0] _0339_;
  wire [2:0] _0340_;
  wire [3:0] _0341_;
  wire [2:0] _0342_;
  wire [3:0] _0343_;
  wire [2:0] _0344_;
  wire [3:0] _0345_;
  wire _0346_;
  wire _0347_;
  wire [1:0] _0348_;
  wire _0349_;
  wire [303:0] _0350_;
  wire [1:0] _0351_;
  wire [66:0] _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire [1:0] _0373_;
  wire [1:0] _0374_;
  wire _0375_;
  wire _0376_;
  wire [1:0] _0377_;
  wire [1:0] _0378_;
  wire _0379_;
  wire _0380_;
  wire [1:0] _0381_;
  wire [1:0] _0382_;
  wire _0383_;
  wire _0384_;
  wire [1:0] _0385_;
  wire [1:0] _0386_;
  wire _0387_;
  wire _0388_;
  wire [1:0] _0389_;
  wire [1:0] _0390_;
  wire _0391_;
  wire _0392_;
  wire [1:0] _0393_;
  wire [1:0] _0394_;
  wire _0395_;
  wire _0396_;
  wire [1:0] _0397_;
  wire [1:0] _0398_;
  wire _0399_;
  wire _0400_;
  wire [1:0] _0401_;
  wire [1:0] _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire [7:0] _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire [7:0] _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire [7:0] _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire [7:0] _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire [7:0] _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire [7:0] _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire [7:0] _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire [7:0] _0490_;
  wire _0491_;
  wire [22:0] _0492_;
  wire [22:0] _0493_;
  wire [22:0] _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire [63:0] _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire [63:0] _0816_;
  wire [63:0] _0817_;
  wire _0818_;
  wire [63:0] _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire [63:0] _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire [1:0] _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire [1:0] _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire [1:0] _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire [1:0] _0860_;
  wire _0861_;
  wire _0862_;
  wire [63:0] _0863_;
  wire [31:0] _0864_;
  wire [95:0] _0865_;
  wire [1:0] _0866_;
  wire [95:0] _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire [95:0] _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire [1:0] _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire [1:0] _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire [1:0] _0893_;
  wire _0894_;
  wire [95:0] _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire [1:0] _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire [1:0] _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire [31:0] _0918_;
  wire [11:0] _0919_;
  wire _0920_;
  wire [11:0] _0921_;
  wire [1:0] _0922_;
  wire _0923_;
  wire _0924_;
  wire [95:0] _0925_;
  wire [11:0] _0926_;
  wire [1:0] _0927_;
  wire _0928_;
  wire _0929_;
  wire [63:0] _0930_;
  wire [31:0] _0931_;
  wire [11:0] _0932_;
  wire [1:0] _0933_;
  wire _0934_;
  wire _0935_;
  wire [95:0] _0936_;
  wire [75:0] _0937_;
  wire [1:0] _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire [63:0] _0944_;
  wire _0945_;
  wire [71:0] _0946_;
  wire [7:0] _0947_;
  wire [63:0] _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire [7:0] _0957_;
  wire [7:0] _0958_;
  wire [7:0] _0959_;
  wire [7:0] _0960_;
  wire [7:0] _0961_;
  wire [7:0] _0962_;
  wire [7:0] _0963_;
  wire [7:0] _0964_;
  wire [7:0] _0965_;
  wire [7:0] _0966_;
  wire [7:0] _0967_;
  wire [7:0] _0968_;
  wire [7:0] _0969_;
  wire [7:0] _0970_;
  wire [7:0] _0971_;
  wire [7:0] _0972_;
  wire [7:0] _0973_;
  wire [7:0] _0974_;
  wire [7:0] _0975_;
  wire [7:0] _0976_;
  wire [7:0] _0977_;
  wire [7:0] _0978_;
  wire [7:0] _0979_;
  wire [7:0] _0980_;
  wire [7:0] _0981_;
  wire [7:0] _0982_;
  wire [7:0] _0983_;
  wire [7:0] _0984_;
  wire [7:0] _0985_;
  wire [7:0] _0986_;
  wire [7:0] _0987_;
  wire [7:0] _0988_;
  wire [7:0] _0989_;
  wire [7:0] _0990_;
  wire [7:0] _0991_;
  wire [7:0] _0992_;
  wire [7:0] _0993_;
  wire [7:0] _0994_;
  wire [7:0] _0995_;
  wire [7:0] _0996_;
  wire [7:0] _0997_;
  wire [7:0] _0998_;
  wire [7:0] _0999_;
  wire [7:0] _1000_;
  wire [7:0] _1001_;
  wire [7:0] _1002_;
  wire [7:0] _1003_;
  wire [7:0] _1004_;
  wire busy;
  input clk;
  wire clk;
  wire complete;
  input \d_in.cache_paradox ;
  wire \d_in.cache_paradox ;
  input [63:0] \d_in.data ;
  wire [63:0] \d_in.data ;
  input \d_in.error ;
  wire \d_in.error ;
  input \d_in.store_done ;
  wire \d_in.store_done ;
  input \d_in.valid ;
  wire \d_in.valid ;
  output [63:0] \d_out.addr ;
  wire [63:0] \d_out.addr ;
  output \d_out.atomic ;
  wire \d_out.atomic ;
  output \d_out.atomic_last ;
  wire \d_out.atomic_last ;
  output [7:0] \d_out.byte_sel ;
  wire [7:0] \d_out.byte_sel ;
  output [63:0] \d_out.data ;
  wire [63:0] \d_out.data ;
  output \d_out.dcbz ;
  wire \d_out.dcbz ;
  output \d_out.hold ;
  wire \d_out.hold ;
  output \d_out.load ;
  wire \d_out.load ;
  output \d_out.nc ;
  wire \d_out.nc ;
  output \d_out.priv_mode ;
  wire \d_out.priv_mode ;
  output \d_out.reserve ;
  wire \d_out.reserve ;
  output \d_out.valid ;
  wire \d_out.valid ;
  output \d_out.virt_mode ;
  wire \d_out.virt_mode ;
  input dc_stall;
  wire dc_stall;
  output \e_out.busy ;
  wire \e_out.busy ;
  output \e_out.in_progress ;
  wire \e_out.in_progress ;
  output \e_out.interrupt ;
  wire \e_out.interrupt ;
  output \events.itlb_miss ;
  wire \events.itlb_miss ;
  output \events.load_complete ;
  wire \events.load_complete ;
  output \events.store_complete ;
  wire \events.store_complete ;
  wire flushing;
  wire in_progress;
  input [63:0] \l_in.addr1 ;
  wire [63:0] \l_in.addr1 ;
  input [63:0] \l_in.addr2 ;
  wire [63:0] \l_in.addr2 ;
  input \l_in.byte_reverse ;
  wire \l_in.byte_reverse ;
  input \l_in.ci ;
  wire \l_in.ci ;
  input [63:0] \l_in.data ;
  wire [63:0] \l_in.data ;
  input [31:0] \l_in.insn ;
  wire [31:0] \l_in.insn ;
  input [2:0] \l_in.instr_tag ;
  wire [2:0] \l_in.instr_tag ;
  input \l_in.is_32bit ;
  wire \l_in.is_32bit ;
  input [3:0] \l_in.length ;
  wire [3:0] \l_in.length ;
  input \l_in.mode_32bit ;
  wire \l_in.mode_32bit ;
  input [63:0] \l_in.msr ;
  wire [63:0] \l_in.msr ;
  input [63:0] \l_in.nia ;
  wire [63:0] \l_in.nia ;
  input [5:0] \l_in.op ;
  wire [5:0] \l_in.op ;
  input \l_in.priv_mode ;
  wire \l_in.priv_mode ;
  input \l_in.rc ;
  wire \l_in.rc ;
  input \l_in.repeat ;
  wire \l_in.repeat ;
  input \l_in.reserve ;
  wire \l_in.reserve ;
  input \l_in.second ;
  wire \l_in.second ;
  input \l_in.sign_extend ;
  wire \l_in.sign_extend ;
  input \l_in.update ;
  wire \l_in.update ;
  input \l_in.valid ;
  wire \l_in.valid ;
  input \l_in.virt_mode ;
  wire \l_in.virt_mode ;
  input [6:0] \l_in.write_reg ;
  wire [6:0] \l_in.write_reg ;
  input [4:0] \l_in.xerc ;
  wire [4:0] \l_in.xerc ;
  output [2:0] \l_out.instr_tag ;
  wire [2:0] \l_out.instr_tag ;
  output \l_out.interrupt ;
  wire \l_out.interrupt ;
  output [11:0] \l_out.intr_vec ;
  wire [11:0] \l_out.intr_vec ;
  output \l_out.rc ;
  wire \l_out.rc ;
  output [63:0] \l_out.srr0 ;
  wire [63:0] \l_out.srr0 ;
  output [15:0] \l_out.srr1 ;
  wire [15:0] \l_out.srr1 ;
  output \l_out.store_done ;
  wire \l_out.store_done ;
  output \l_out.valid ;
  wire \l_out.valid ;
  output [63:0] \l_out.write_data ;
  wire [63:0] \l_out.write_data ;
  output \l_out.write_enable ;
  wire \l_out.write_enable ;
  output [6:0] \l_out.write_reg ;
  wire [6:0] \l_out.write_reg ;
  output [4:0] \l_out.xerc ;
  wire [4:0] \l_out.xerc ;
  wire [63:0] load_dp_data;
  output [9:0] log_out;
  wire [9:0] log_out;
  input \m_in.badtree ;
  wire \m_in.badtree ;
  input \m_in.done ;
  wire \m_in.done ;
  input \m_in.err ;
  wire \m_in.err ;
  input \m_in.invalid ;
  wire \m_in.invalid ;
  input \m_in.perm_error ;
  wire \m_in.perm_error ;
  input \m_in.rc_error ;
  wire \m_in.rc_error ;
  input \m_in.segerr ;
  wire \m_in.segerr ;
  input [63:0] \m_in.sprval ;
  wire [63:0] \m_in.sprval ;
  output [63:0] \m_out.addr ;
  wire [63:0] \m_out.addr ;
  output \m_out.iside ;
  wire \m_out.iside ;
  output \m_out.load ;
  wire \m_out.load ;
  output \m_out.mtspr ;
  wire \m_out.mtspr ;
  output \m_out.priv ;
  wire \m_out.priv ;
  output [63:0] \m_out.rs ;
  wire [63:0] \m_out.rs ;
  output \m_out.slbia ;
  wire \m_out.slbia ;
  output [9:0] \m_out.sprn ;
  wire [9:0] \m_out.sprn ;
  output \m_out.tlbie ;
  wire \m_out.tlbie ;
  output \m_out.valid ;
  wire \m_out.valid ;
  wire [337:0] r1;
  wire [337:0] r1in;
  wire [373:0] r2;
  wire [373:0] r2in;
  wire [380:0] r3;
  wire [380:0] r3in;
  wire [272:0] req_in;
  input rst;
  wire rst;
  wire stage1_dcreq;
  wire stage1_dreq;
  wire stage1_issue_enable;
  wire [272:0] stage1_req;
  wire stage2_busy_next;
  wire stage3_busy_next;
  wire [63:0] store_data;
  wire [31:0] store_sp_data;
  assign _0000_ = _0290_[0] ? r1[109:102] : r1[101:94];
  assign _0001_ = _0290_[0] ? r1[141:134] : r1[133:126];
  assign _0002_ = _0292_[0] ? r1[109:102] : r1[101:94];
  assign _0003_ = _0292_[0] ? r1[141:134] : r1[133:126];
  assign _0004_ = _0294_[0] ? r1[109:102] : r1[101:94];
  assign _0005_ = _0294_[0] ? r1[141:134] : r1[133:126];
  assign _0006_ = _0296_[0] ? r1[109:102] : r1[101:94];
  assign _0007_ = _0296_[0] ? r1[141:134] : r1[133:126];
  assign _0008_ = _0298_[0] ? r1[109:102] : r1[101:94];
  assign _0009_ = _0298_[0] ? r1[141:134] : r1[133:126];
  assign _0010_ = _0300_[0] ? r1[109:102] : r1[101:94];
  assign _0011_ = _0300_[0] ? r1[141:134] : r1[133:126];
  assign _0012_ = _0302_[0] ? r1[109:102] : r1[101:94];
  assign _0013_ = _0302_[0] ? r1[141:134] : r1[133:126];
  assign _0014_ = _0304_[0] ? r1[109:102] : r1[101:94];
  assign _0015_ = _0304_[0] ? r1[141:134] : r1[133:126];
  assign _0016_ = r2[294] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0017_ = r2[294] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0018_ = r2[291] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0019_ = r2[291] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0020_ = r2[288] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0021_ = r2[288] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0022_ = r2[285] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0023_ = r2[285] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0024_ = r2[282] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0025_ = r2[282] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0026_ = r2[279] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0027_ = r2[279] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0028_ = r2[276] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0029_ = r2[276] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0030_ = r2[273] ? \d_in.data [15:8] : \d_in.data [7:0];
  assign _0031_ = r2[273] ? \d_in.data [47:40] : \d_in.data [39:32];
  assign _0032_ = _0290_[0] ? r1[125:118] : r1[117:110];
  assign _0033_ = _0290_[0] ? r1[157:150] : r1[149:142];
  assign _0034_ = _0292_[0] ? r1[125:118] : r1[117:110];
  assign _0035_ = _0292_[0] ? r1[157:150] : r1[149:142];
  assign _0036_ = _0294_[0] ? r1[125:118] : r1[117:110];
  assign _0037_ = _0294_[0] ? r1[157:150] : r1[149:142];
  assign _0038_ = _0296_[0] ? r1[125:118] : r1[117:110];
  assign _0039_ = _0296_[0] ? r1[157:150] : r1[149:142];
  assign _0040_ = _0298_[0] ? r1[125:118] : r1[117:110];
  assign _0041_ = _0298_[0] ? r1[157:150] : r1[149:142];
  assign _0042_ = _0300_[0] ? r1[125:118] : r1[117:110];
  assign _0043_ = _0300_[0] ? r1[157:150] : r1[149:142];
  assign _0044_ = _0302_[0] ? r1[125:118] : r1[117:110];
  assign _0045_ = _0302_[0] ? r1[157:150] : r1[149:142];
  assign _0046_ = _0304_[0] ? r1[125:118] : r1[117:110];
  assign _0047_ = _0304_[0] ? r1[157:150] : r1[149:142];
  assign _0048_ = r2[294] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0049_ = r2[294] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0050_ = r2[291] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0051_ = r2[291] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0052_ = r2[288] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0053_ = r2[288] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0054_ = r2[285] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0055_ = r2[285] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0056_ = r2[282] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0057_ = r2[282] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0058_ = r2[279] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0059_ = r2[279] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0060_ = r2[276] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0061_ = r2[276] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0062_ = r2[273] ? \d_in.data [31:24] : \d_in.data [23:16];
  assign _0063_ = r2[273] ? \d_in.data [63:56] : \d_in.data [55:48];
  assign _0957_ = _0290_[1] ? _0032_ : _0000_;
  assign _0958_ = _0290_[1] ? _0033_ : _0001_;
  assign _0960_ = _0292_[1] ? _0034_ : _0002_;
  assign _0961_ = _0292_[1] ? _0035_ : _0003_;
  assign _0963_ = _0294_[1] ? _0036_ : _0004_;
  assign _0964_ = _0294_[1] ? _0037_ : _0005_;
  assign _0966_ = _0296_[1] ? _0038_ : _0006_;
  assign _0967_ = _0296_[1] ? _0039_ : _0007_;
  assign _0969_ = _0298_[1] ? _0040_ : _0008_;
  assign _0970_ = _0298_[1] ? _0041_ : _0009_;
  assign _0972_ = _0300_[1] ? _0042_ : _0010_;
  assign _0973_ = _0300_[1] ? _0043_ : _0011_;
  assign _0975_ = _0302_[1] ? _0044_ : _0012_;
  assign _0976_ = _0302_[1] ? _0045_ : _0013_;
  assign _0978_ = _0304_[1] ? _0046_ : _0014_;
  assign _0979_ = _0304_[1] ? _0047_ : _0015_;
  assign _0981_ = r2[295] ? _0048_ : _0016_;
  assign _0982_ = r2[295] ? _0049_ : _0017_;
  assign _0984_ = r2[292] ? _0050_ : _0018_;
  assign _0985_ = r2[292] ? _0051_ : _0019_;
  assign _0987_ = r2[289] ? _0052_ : _0020_;
  assign _0988_ = r2[289] ? _0053_ : _0021_;
  assign _0990_ = r2[286] ? _0054_ : _0022_;
  assign _0991_ = r2[286] ? _0055_ : _0023_;
  assign _0993_ = r2[283] ? _0056_ : _0024_;
  assign _0994_ = r2[283] ? _0057_ : _0025_;
  assign _0996_ = r2[280] ? _0058_ : _0026_;
  assign _0997_ = r2[280] ? _0059_ : _0027_;
  assign _0999_ = r2[277] ? _0060_ : _0028_;
  assign _1000_ = r2[277] ? _0061_ : _0029_;
  assign _1002_ = r2[274] ? _0062_ : _0030_;
  assign _1003_ = r2[274] ? _0063_ : _0031_;
  assign _0064_ = r1in[0] & r1in[206];
  assign _0065_ = flushing | _0064_;
  assign _0066_ = ~ r3in[285];
  assign _0067_ = _0065_ & _0066_;
  assign _0068_ = rst ? 1'h0 : r1in[0];
  assign _0069_ = rst ? r1[337:1] : r1in[337:1];
  assign _0070_ = rst ? 1'h0 : r2in[0];
  assign _0071_ = rst ? r2[304:1] : r2in[304:1];
  assign _0072_ = rst ? 3'h0 : r2in[307:305];
  assign _0073_ = rst ? r2[373:308] : r2in[373:308];
  assign _0074_ = rst ? 2'h0 : r3in[1:0];
  assign _0075_ = rst ? r3[4:2] : r3in[4:2];
  assign _0076_ = rst ? 1'h0 : r3in[5];
  assign _0077_ = rst ? r3[83:6] : r3in[83:6];
  assign _0078_ = rst ? 1'h0 : r3in[84];
  assign _0079_ = rst ? r3[148:85] : r3in[148:85];
  assign _0080_ = rst ? 96'h000000000000000000000000 : r3in[244:149];
  assign _0081_ = rst ? r3[283:245] : r3in[283:245];
  assign _0082_ = rst ? 2'h1 : r3in[285:284];
  assign _0083_ = rst ? r3[380:286] : r3in[380:286];
  assign _0084_ = rst ? 1'h0 : _0067_;
  always @(posedge clk)
    _0085_ <= { _0069_, _0068_ };
  always @(posedge clk)
    _0086_ <= { _0073_, _0072_, _0071_, _0070_ };
  always @(posedge clk)
    _0087_ <= { _0083_, _0082_, _0081_, _0080_, _0079_, _0078_, _0077_, _0076_, _0075_, _0074_ };
  always @(posedge clk)
    _0088_ <= _0084_;
  always @(posedge clk)
    _0089_ <= stage1_dcreq;
  assign _0090_ = \l_in.data [62:52] > 11'h380;
  assign _0091_ = \l_in.data [62:52] >= 11'h36a;
  assign _0092_ = 5'h00 - \l_in.data [56:52];
  assign _0093_ = _0092_[1:0] == 2'h0;
  assign _0094_ = _0092_[1:0] == 2'h1;
  assign _0095_ = _0092_[1:0] == 2'h2;
  function [22:0] \19547 ;
    input [22:0] a;
    input [68:0] b;
    input [2:0] s;
    (* parallel_case *)
    casez (s)
      3'b??1:
        \19547  = b[22:0];
      3'b?1?:
        \19547  = b[45:23];
      3'b1??:
        \19547  = b[68:46];
      default:
        \19547  = a;
    endcase
  endfunction
  assign _0096_ = \19547 ({ 4'h1, \l_in.data [51:33] }, { 3'h1, \l_in.data [51:32], 2'h1, \l_in.data [51:31], 1'h1, \l_in.data [51:30] }, { _0095_, _0094_, _0093_ });
  assign _0097_ = _0092_[4:2] == 3'h0;
  assign _0098_ = _0092_[4:2] == 3'h1;
  assign _0099_ = _0092_[4:2] == 3'h2;
  assign _0100_ = _0092_[4:2] == 3'h3;
  assign _0101_ = _0092_[4:2] == 3'h4;
  function [22:0] \19576 ;
    input [22:0] a;
    input [114:0] b;
    input [4:0] s;
    (* parallel_case *)
    casez (s)
      5'b????1:
        \19576  = b[22:0];
      5'b???1?:
        \19576  = b[45:23];
      5'b??1??:
        \19576  = b[68:46];
      5'b?1???:
        \19576  = b[91:69];
      5'b1????:
        \19576  = b[114:92];
      default:
        \19576  = a;
    endcase
  endfunction
  assign _0102_ = \19576 ({ 20'h00000, _0096_[22:20] }, { 16'h0000, _0096_[22:16], 12'h000, _0096_[22:12], 8'h00, _0096_[22:8], 4'h0, _0096_[22:4], _0096_ }, { _0101_, _0100_, _0099_, _0098_, _0097_ });
  assign _0103_ = _0091_ ? _0102_ : 23'h000000;
  assign _0104_ = _0090_ ? \l_in.data [51:29] : _0103_;
  assign _0105_ = _0090_ ? { \l_in.data [62], \l_in.data [58:52] } : 8'h00;
  assign _0106_ = | r3[275:268];
  assign _0107_ = & r3[275:268];
  assign _0108_ = 11'h380 + { 3'h0, r3[275:268] };
  assign _0109_ = ~ r3[277];
  assign _0110_ = 11'h380 - { 5'h00, r3[283:278] };
  assign _0111_ = r3[282:278] + 5'h01;
  assign _0112_ = _0109_ ? 11'h000 : _0110_;
  assign _0113_ = _0109_ ? 5'h00 : _0111_;
  assign _0114_ = _0106_ ? _0108_ : _0112_;
  assign _0115_ = _0106_ ? 5'h00 : _0113_;
  assign _0116_ = _0107_ ? 11'h7ff : _0114_;
  assign _0117_ = _0107_ ? 5'h00 : _0115_;
  assign _0118_ = _0117_[1:0] == 2'h0;
  assign _0119_ = _0117_[1:0] == 2'h1;
  assign _0120_ = _0117_[1:0] == 2'h2;
  function [22:0] \19656 ;
    input [22:0] a;
    input [68:0] b;
    input [2:0] s;
    (* parallel_case *)
    casez (s)
      3'b??1:
        \19656  = b[22:0];
      3'b?1?:
        \19656  = b[45:23];
      3'b1??:
        \19656  = b[68:46];
      default:
        \19656  = a;
    endcase
  endfunction
  assign _0121_ = \19656 ({ r3[264:245], 3'h0 }, { r3[265:245], 2'h0, r3[266:245], 1'h0, r3[267:245] }, { _0120_, _0119_, _0118_ });
  assign _0122_ = _0117_[4:2] == 3'h0;
  assign _0123_ = _0117_[4:2] == 3'h1;
  assign _0124_ = _0117_[4:2] == 3'h2;
  assign _0125_ = _0117_[4:2] == 3'h3;
  assign _0126_ = _0117_[4:2] == 3'h4;
  function [22:0] \19685 ;
    input [22:0] a;
    input [114:0] b;
    input [4:0] s;
    (* parallel_case *)
    casez (s)
      5'b????1:
        \19685  = b[22:0];
      5'b???1?:
        \19685  = b[45:23];
      5'b??1??:
        \19685  = b[68:46];
      5'b?1???:
        \19685  = b[91:69];
      5'b1????:
        \19685  = b[114:92];
      default:
        \19685  = a;
    endcase
  endfunction
  assign _0127_ = \19685 ({ _0121_[2:0], 20'h00000 }, { _0121_[6:0], 16'h0000, _0121_[10:0], 12'h000, _0121_[14:0], 8'h00, _0121_[18:0], 4'h0, _0121_ }, { _0126_, _0125_, _0124_, _0123_, _0122_ });
  assign _0128_ = \l_in.addr1  + \l_in.addr2 ;
  assign _0129_ = 1'h1 & \l_in.is_32bit ;
  assign _0130_ = _0129_ ? { 32'h00000000, store_sp_data } : \l_in.data ;
  assign _0131_ = ~ \l_in.update ;
  assign _0132_ = r1[337:277] + 61'h0000000000000001;
  assign _0133_ = _0131_ ? _0132_[60:29] : r1[337:306];
  assign _0134_ = \l_in.second  ? _0133_ : _0128_[63:32];
  assign _0135_ = \l_in.mode_32bit  ? 32'd0 : _0134_;
  assign _0136_ = _0131_ ? { _0132_[28:0], r1[276:274] } : r1[305:274];
  assign _0137_ = \l_in.second  ? _0136_ : _0128_[31:0];
  assign _0138_ = _0137_[31:28] == 4'hc;
  assign _0139_ = ~ \l_in.virt_mode ;
  assign _0140_ = _0138_ & _0139_;
  assign _0141_ = _0140_ ? 1'h1 : \l_in.ci ;
  assign _0142_ = \l_in.length [2:0] - 3'h1;
  assign _0143_ = \l_in.length  == 4'h1;
  assign _0144_ = \l_in.length  == 4'h2;
  assign _0145_ = \l_in.length  == 4'h4;
  assign _0146_ = \l_in.length  == 4'h8;
  function [7:0] \19827 ;
    input [7:0] a;
    input [31:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \19827  = b[7:0];
      4'b??1?:
        \19827  = b[15:8];
      4'b?1??:
        \19827  = b[23:16];
      4'b1???:
        \19827  = b[31:24];
      default:
        \19827  = a;
    endcase
  endfunction
  assign _0147_ = \19827 (8'h00, 32'd4279173889, { _0146_, _0145_, _0144_, _0143_ });
  assign _0148_ = { 8'h00, _0147_ } << { 28'h0000000, _0137_[2:0] };
  assign _0149_ = _0148_[15:8] != 8'h00;
  assign _0150_ = _0149_ ? 1'h1 : 1'h0;
  assign _0151_ = _0142_ & _0137_[2:0];
  assign _0152_ = | _0151_;
  assign _0153_ = \l_in.reserve  & _0152_;
  assign _0154_ = ~ \l_in.second ;
  assign _0155_ = \l_in.repeat  & _0154_;
  assign _0156_ = ~ \l_in.update ;
  assign _0157_ = _0155_ & _0156_;
  assign _0158_ = _0157_ & _0137_[3];
  assign _0159_ = \l_in.op  == 6'h1f;
  assign _0160_ = ~ \l_in.byte_reverse ;
  assign _0161_ = _0159_ & _0160_;
  assign _0162_ = \l_in.reserve  | _0161_;
  assign _0163_ = _0164_ ? 1'h1 : _0153_;
  assign _0164_ = _0158_ & _0162_;
  assign _0165_ = _0158_ ? 1'h1 : _0152_;
  assign _0166_ = ~ _0165_;
  assign _0167_ = ~ _0165_;
  assign _0168_ = ~ \l_in.repeat ;
  assign _0169_ = \l_in.second  | _0168_;
  assign _0170_ = _0167_ & _0169_;
  assign _0171_ = \l_in.op  == 6'h20;
  assign _0172_ = ~ \l_in.update ;
  assign _0173_ = ~ \l_in.second ;
  assign _0174_ = _0172_ | _0173_;
  assign _0175_ = 1'h1 & \l_in.is_32bit ;
  assign _0176_ = _0179_ ? 1'h1 : 1'h0;
  assign _0177_ = _0174_ ? 1'h1 : 1'h0;
  assign _0178_ = _0174_ ? 1'h0 : 1'h1;
  assign _0179_ = _0174_ & _0175_;
  assign _0180_ = \l_in.op  == 6'h1f;
  assign _0181_ = \l_in.op  == 6'h14;
  assign _0182_ = \l_in.op  == 6'h38;
  assign _0183_ = \l_in.op  == 6'h24;
  assign _0184_ = \l_in.insn [14] | \l_in.insn [11];
  assign _0185_ = \l_in.op  == 6'h28;
  assign _0186_ = \l_in.op  == 6'h3d;
  function [0:0] \19934 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19934  = b[0:0];
      7'b?????1?:
        \19934  = b[1:1];
      7'b????1??:
        \19934  = b[2:2];
      7'b???1???:
        \19934  = b[3:3];
      7'b??1????:
        \19934  = b[4:4];
      7'b?1?????:
        \19934  = b[5:5];
      7'b1??????:
        \19934  = b[6:6];
      default:
        \19934  = a;
    endcase
  endfunction
  assign _0187_ = \19934 (1'h0, { 5'h00, _0177_, 1'h0 }, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19936 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19936  = b[0:0];
      7'b?????1?:
        \19936  = b[1:1];
      7'b????1??:
        \19936  = b[2:2];
      7'b???1???:
        \19936  = b[3:3];
      7'b??1????:
        \19936  = b[4:4];
      7'b?1?????:
        \19936  = b[5:5];
      7'b1??????:
        \19936  = b[6:6];
      default:
        \19936  = a;
    endcase
  endfunction
  assign _0188_ = \19936 (1'h0, 7'h01, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19938 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19938  = b[0:0];
      7'b?????1?:
        \19938  = b[1:1];
      7'b????1??:
        \19938  = b[2:2];
      7'b???1???:
        \19938  = b[3:3];
      7'b??1????:
        \19938  = b[4:4];
      7'b?1?????:
        \19938  = b[5:5];
      7'b1??????:
        \19938  = b[6:6];
      default:
        \19938  = a;
    endcase
  endfunction
  assign _0189_ = \19938 (1'h0, 7'h08, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19940 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19940  = b[0:0];
      7'b?????1?:
        \19940  = b[1:1];
      7'b????1??:
        \19940  = b[2:2];
      7'b???1???:
        \19940  = b[3:3];
      7'b??1????:
        \19940  = b[4:4];
      7'b?1?????:
        \19940  = b[5:5];
      7'b1??????:
        \19940  = b[6:6];
      default:
        \19940  = a;
    endcase
  endfunction
  assign _0190_ = \19940 (1'h0, 7'h04, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19942 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19942  = b[0:0];
      7'b?????1?:
        \19942  = b[1:1];
      7'b????1??:
        \19942  = b[2:2];
      7'b???1???:
        \19942  = b[3:3];
      7'b??1????:
        \19942  = b[4:4];
      7'b?1?????:
        \19942  = b[5:5];
      7'b1??????:
        \19942  = b[6:6];
      default:
        \19942  = a;
    endcase
  endfunction
  assign _0191_ = \19942 (1'h0, 7'h10, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19944 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19944  = b[0:0];
      7'b?????1?:
        \19944  = b[1:1];
      7'b????1??:
        \19944  = b[2:2];
      7'b???1???:
        \19944  = b[3:3];
      7'b??1????:
        \19944  = b[4:4];
      7'b?1?????:
        \19944  = b[5:5];
      7'b1??????:
        \19944  = b[6:6];
      default:
        \19944  = a;
    endcase
  endfunction
  assign _0192_ = \19944 (1'h0, 7'h20, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19946 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19946  = b[0:0];
      7'b?????1?:
        \19946  = b[1:1];
      7'b????1??:
        \19946  = b[2:2];
      7'b???1???:
        \19946  = b[3:3];
      7'b??1????:
        \19946  = b[4:4];
      7'b?1?????:
        \19946  = b[5:5];
      7'b1??????:
        \19946  = b[6:6];
      default:
        \19946  = a;
    endcase
  endfunction
  assign _0193_ = \19946 (1'h0, { 1'h1, _0184_, 5'h08 }, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19948 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19948  = b[0:0];
      7'b?????1?:
        \19948  = b[1:1];
      7'b????1??:
        \19948  = b[2:2];
      7'b???1???:
        \19948  = b[3:3];
      7'b??1????:
        \19948  = b[4:4];
      7'b?1?????:
        \19948  = b[5:5];
      7'b1??????:
        \19948  = b[6:6];
      default:
        \19948  = a;
    endcase
  endfunction
  assign _0194_ = \19948 (1'h0, 7'h40, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19950 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19950  = b[0:0];
      7'b?????1?:
        \19950  = b[1:1];
      7'b????1??:
        \19950  = b[2:2];
      7'b???1???:
        \19950  = b[3:3];
      7'b??1????:
        \19950  = b[4:4];
      7'b?1?????:
        \19950  = b[5:5];
      7'b1??????:
        \19950  = b[6:6];
      default:
        \19950  = a;
    endcase
  endfunction
  assign _0195_ = \19950 (1'h0, { 5'h00, _0178_, 1'h0 }, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [63:0] \19951 ;
    input [63:0] a;
    input [447:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19951  = b[63:0];
      7'b?????1?:
        \19951  = b[127:64];
      7'b????1??:
        \19951  = b[191:128];
      7'b???1???:
        \19951  = b[255:192];
      7'b??1????:
        \19951  = b[319:256];
      7'b?1?????:
        \19951  = b[383:320];
      7'b1??????:
        \19951  = b[447:384];
      default:
        \19951  = a;
    endcase
  endfunction
  assign _0196_ = \19951 ({ _0135_, _0137_ }, { \l_in.nia , _0135_, _0137_, _0135_, _0137_, \l_in.addr2 , _0135_, _0137_, _0135_, _0137_, _0135_, _0137_ }, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19952 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19952  = b[0:0];
      7'b?????1?:
        \19952  = b[1:1];
      7'b????1??:
        \19952  = b[2:2];
      7'b???1???:
        \19952  = b[3:3];
      7'b??1????:
        \19952  = b[4:4];
      7'b?1?????:
        \19952  = b[5:5];
      7'b1??????:
        \19952  = b[6:6];
      default:
        \19952  = a;
    endcase
  endfunction
  assign _0197_ = \19952 (1'h0, { 5'h00, _0176_, 1'h0 }, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19953 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19953  = b[0:0];
      7'b?????1?:
        \19953  = b[1:1];
      7'b????1??:
        \19953  = b[2:2];
      7'b???1???:
        \19953  = b[3:3];
      7'b??1????:
        \19953  = b[4:4];
      7'b?1?????:
        \19953  = b[5:5];
      7'b1??????:
        \19953  = b[6:6];
      default:
        \19953  = a;
    endcase
  endfunction
  assign _0198_ = \19953 (1'h0, { 3'h0, \l_in.insn [7], 3'h0 }, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  function [0:0] \19954 ;
    input [0:0] a;
    input [6:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \19954  = b[0:0];
      7'b?????1?:
        \19954  = b[1:1];
      7'b????1??:
        \19954  = b[2:2];
      7'b???1???:
        \19954  = b[3:3];
      7'b??1????:
        \19954  = b[4:4];
      7'b?1?????:
        \19954  = b[5:5];
      7'b1??????:
        \19954  = b[6:6];
      default:
        \19954  = a;
    endcase
  endfunction
  assign _0199_ = \19954 (_0163_, { _0163_, _0163_, _0163_, _0163_, _0141_, _0163_, _0163_ }, { _0186_, _0185_, _0183_, _0182_, _0181_, _0180_, _0171_ });
  assign _0200_ = _0187_ | _0188_;
  assign _0201_ = _0200_ | _0190_;
  assign _0202_ = \l_in.valid  & _0201_;
  assign _0203_ = ~ _0199_;
  assign _0204_ = _0202_ & _0203_;
  assign _0205_ = \l_in.length [2:0] - 3'h1;
  assign _0206_ = \l_in.byte_reverse  ? _0205_ : 3'h0;
  assign _0207_ = ~ r1[273];
  assign _0208_ = r1[1] & _0207_;
  assign _0209_ = r1[273] & \d_in.error ;
  assign _0210_ = _0208_ | _0209_;
  assign _0211_ = _0210_ | stage2_busy_next;
  assign _0212_ = r1[1] & r1[208];
  assign _0213_ = ~ r1[207];
  assign _0214_ = _0212_ & _0213_;
  assign _0215_ = _0211_ | _0214_;
  assign _0216_ = r1[0] & _0215_;
  assign _0217_ = r2[305] & \d_in.valid ;
  assign _0218_ = r2[307] | _0217_;
  assign _0219_ = r2[306] & \m_in.done ;
  assign _0220_ = _0218_ | _0219_;
  assign _0221_ = _0220_ | r3[84];
  assign _0222_ = ~ complete;
  assign _0223_ = r2[0] & _0222_;
  assign _0224_ = r1[0] | _0223_;
  assign _0225_ = r1[0] & r1[8];
  assign _0226_ = ~ _0225_;
  assign _0227_ = r3[284] & _0226_;
  assign _0228_ = r2[0] & r2[8];
  assign _0229_ = ~ _0228_;
  assign _0230_ = _0227_ & _0229_;
  assign _0231_ = ~ busy;
  assign _0232_ = flushing ? 1'h0 : req_in[1];
  assign _0233_ = \l_in.valid  & _0232_;
  assign _0234_ = \l_in.valid  ? req_in[77:14] : r1[337:274];
  assign _0235_ = _0231_ ? _0233_ : 1'h0;
  assign _0236_ = ~ r1[273];
  assign _0237_ = r1[1] & _0236_;
  assign _0238_ = r1[273] & \d_in.error ;
  assign _0239_ = ~ stage2_busy_next;
  assign _0240_ = r1[1] & r1[208];
  assign _0241_ = ~ r1[207];
  assign _0242_ = _0240_ & _0241_;
  assign _0243_ = r1[77:17] + 61'h0000000000000001;
  assign _0244_ = r1[13] ? 1'h0 : _0243_[29];
  assign _0245_ = _0231_ ? req_in[85:14] : r1[85:14];
  assign _0246_ = _0242_ ? { r1[93:86], _0243_[60:30], _0244_, _0243_[28:0], 3'h0 } : _0245_;
  assign _0247_ = _0231_ ? req_in[207] : r1[207];
  assign _0248_ = _0242_ ? 1'h1 : _0247_;
  assign _0249_ = _0254_ ? 1'h1 : _0235_;
  assign _0250_ = _0231_ ? req_in[85:14] : r1[85:14];
  assign _0251_ = _0239_ ? _0246_ : _0250_;
  assign _0252_ = _0231_ ? req_in[207] : r1[207];
  assign _0253_ = _0239_ ? _0248_ : _0252_;
  assign _0254_ = _0239_ & _0242_;
  assign _0255_ = _0231_ ? 1'h0 : r1[273];
  assign _0256_ = _0238_ ? 1'h0 : _0255_;
  assign _0257_ = _0231_ ? req_in[85:14] : r1[85:14];
  assign _0258_ = _0238_ ? _0257_ : _0251_;
  assign _0259_ = _0231_ ? req_in[207] : r1[207];
  assign _0260_ = _0238_ ? _0259_ : _0253_;
  assign _0261_ = _0238_ ? _0235_ : _0249_;
  assign _0262_ = _0231_ ? 1'h0 : r1[273];
  assign _0263_ = _0237_ ? _0262_ : _0256_;
  assign _0264_ = _0231_ ? req_in[85:14] : r1[85:14];
  assign _0265_ = _0237_ ? _0264_ : _0258_;
  assign _0266_ = _0231_ ? req_in[207] : r1[207];
  assign _0267_ = _0237_ ? _0266_ : _0260_;
  assign _0268_ = _0237_ ? 1'h1 : _0261_;
  assign _0269_ = _0231_ ? 1'h0 : r1[273];
  assign _0270_ = r1[0] ? _0263_ : _0269_;
  assign _0271_ = _0231_ ? _0234_ : r1[337:274];
  assign _0272_ = _0231_ ? req_in[85:14] : r1[85:14];
  assign _0273_ = r1[0] ? _0265_ : _0272_;
  assign _0274_ = _0231_ ? req_in[207] : r1[207];
  assign _0275_ = r1[0] ? _0267_ : _0274_;
  assign _0276_ = _0231_ ? req_in[272:208] : r1[272:208];
  assign _0277_ = _0231_ ? req_in[206:86] : r1[206:86];
  assign _0278_ = r1[0] ? _0268_ : _0235_;
  assign _0279_ = _0231_ ? req_in[0] : r1[0];
  assign _0280_ = r3in[285] ? 1'h0 : _0279_;
  assign _0281_ = _0231_ ? { req_in[13:2], _0232_ } : r1[13:1];
  assign _0282_ = r3in[285] ? 1'h0 : _0278_;
  assign _0283_ = _0282_ & stage1_issue_enable;
  assign _0284_ = ~ \d_in.error ;
  assign _0285_ = _0283_ & _0284_;
  assign _0286_ = ~ dc_stall;
  assign _0287_ = _0285_ & _0286_;
  assign _0288_ = _0282_ ? _0287_ : _0270_;
  assign _0289_ = 3'h0 - r1[276:274];
  assign _0290_ = _0289_ ^ r1[179:177];
  assign _0291_ = 3'h1 - r1[276:274];
  assign _0292_ = _0291_ ^ r1[179:177];
  assign _0293_ = 3'h2 - r1[276:274];
  assign _0294_ = _0293_ ^ r1[179:177];
  assign _0295_ = 3'h3 - r1[276:274];
  assign _0296_ = _0295_ ^ r1[179:177];
  assign _0297_ = 3'h4 - r1[276:274];
  assign _0298_ = _0297_ ^ r1[179:177];
  assign _0299_ = 3'h5 - r1[276:274];
  assign _0300_ = _0299_ ^ r1[179:177];
  assign _0301_ = 3'h6 - r1[276:274];
  assign _0302_ = _0301_ ^ r1[179:177];
  assign _0303_ = 3'h7 - r1[276:274];
  assign _0304_ = _0303_ ^ r1[179:177];
  assign _0305_ = ~ stage3_busy_next;
  assign _0306_ = ~ r1[0];
  assign _0307_ = _0306_ | r1[273];
  assign _0308_ = ~ r1[1];
  assign _0309_ = _0307_ | _0308_;
  assign _0310_ = _0305_ & _0309_;
  assign _0311_ = r1[0] & r1[1];
  assign _0312_ = ~ r1[194];
  assign _0313_ = _0311_ & _0312_;
  assign _0314_ = ~ r1[207];
  assign _0315_ = r1[208] & _0314_;
  assign _0316_ = ~ _0315_;
  assign _0317_ = _0313_ & _0316_;
  assign _0318_ = r1[0] & r1[8];
  assign _0319_ = r1[12] | r1[6];
  assign _0320_ = ~ r1[8];
  assign _0321_ = r1[7] & _0320_;
  assign _0322_ = _0319_ | _0321_;
  assign _0323_ = _0322_ | r1[10];
  assign _0324_ = _0323_ | r1[11];
  assign _0325_ = r1[0] & _0324_;
  assign _0326_ = r1[11] | r1[3];
  assign _0327_ = r1[194] ? 2'h2 : 2'h3;
  assign _0328_ = _0326_ ? 2'h1 : _0327_;
  assign _0329_ = r1[6] ? 2'h0 : _0328_;
  assign _0330_ = 3'h0 ^ r1[179:177];
  assign _0331_ = { 1'h0, _0330_ } + { 1'h0, r1[276:274] };
  assign _0332_ = 3'h1 ^ r1[179:177];
  assign _0333_ = { 1'h0, _0332_ } + { 1'h0, r1[276:274] };
  assign _0334_ = 3'h2 ^ r1[179:177];
  assign _0335_ = { 1'h0, _0334_ } + { 1'h0, r1[276:274] };
  assign _0336_ = 3'h3 ^ r1[179:177];
  assign _0337_ = { 1'h0, _0336_ } + { 1'h0, r1[276:274] };
  assign _0338_ = 3'h4 ^ r1[179:177];
  assign _0339_ = { 1'h0, _0338_ } + { 1'h0, r1[276:274] };
  assign _0340_ = 3'h5 ^ r1[179:177];
  assign _0341_ = { 1'h0, _0340_ } + { 1'h0, r1[276:274] };
  assign _0342_ = 3'h6 ^ r1[179:177];
  assign _0343_ = { 1'h0, _0342_ } + { 1'h0, r1[276:274] };
  assign _0344_ = 3'h7 ^ r1[179:177];
  assign _0345_ = { 1'h0, _0344_ } + { 1'h0, r1[276:274] };
  assign _0346_ = ~ stage3_busy_next;
  assign _0347_ = _0346_ ? 1'h0 : r2[0];
  assign _0348_ = _0346_ ? 2'h0 : r2[306:305];
  assign _0349_ = _0310_ ? r1[0] : _0347_;
  assign _0350_ = _0310_ ? { _0345_[3], _0343_[3], _0341_[3], _0339_[3], _0337_[3], _0335_[3], _0333_[3], _0331_, _0333_[2:0], _0335_[2:0], _0337_[2:0], _0339_[2:0], _0341_[2:0], _0343_[2:0], _0345_[2:0], r1[272:158], store_data, r1[93:1] } : r2[304:1];
  assign _0351_ = _0310_ ? { _0318_, _0317_ } : _0348_;
  assign _0352_ = _0310_ ? { r1[337:274], _0329_, _0325_ } : r2[373:307];
  assign _0353_ = r1[0] & stage3_busy_next;
  assign _0354_ = r3in[285] ? 1'h0 : _0349_;
  assign _0355_ = r2[207] & r2[176];
  assign _0356_ = r2[171] & r3[148];
  assign _0357_ = r2[170] & r3[116];
  assign _0358_ = _0356_ | _0357_;
  assign _0359_ = r2[169] & r3[100];
  assign _0360_ = _0358_ | _0359_;
  assign _0361_ = r2[168] & r3[92];
  assign _0362_ = _0360_ | _0361_;
  assign _0363_ = r2[171] & _1004_[7];
  assign _0364_ = r2[170] & _0992_[7];
  assign _0365_ = _0363_ | _0364_;
  assign _0366_ = r2[169] & _0986_[7];
  assign _0367_ = _0365_ | _0366_;
  assign _0368_ = r2[168] & _0983_[7];
  assign _0369_ = _0367_ | _0368_;
  assign _0370_ = _0355_ ? _0362_ : _0369_;
  assign _0371_ = $signed(32'd0) < $signed({ 28'h0000000, r2[171:168] });
  assign _0372_ = ~ r2[297];
  assign _0373_ = r2[207] ? { 1'h1, _0372_ } : 2'h2;
  assign _0374_ = _0371_ ? _0373_ : 2'h0;
  assign _0375_ = $signed(32'd1) < $signed({ 28'h0000000, r2[171:168] });
  assign _0376_ = ~ r2[298];
  assign _0377_ = r2[207] ? { 1'h1, _0376_ } : 2'h2;
  assign _0378_ = _0375_ ? _0377_ : 2'h0;
  assign _0379_ = $signed(32'd2) < $signed({ 28'h0000000, r2[171:168] });
  assign _0380_ = ~ r2[299];
  assign _0381_ = r2[207] ? { 1'h1, _0380_ } : 2'h2;
  assign _0382_ = _0379_ ? _0381_ : 2'h0;
  assign _0383_ = $signed(32'd3) < $signed({ 28'h0000000, r2[171:168] });
  assign _0384_ = ~ r2[300];
  assign _0385_ = r2[207] ? { 1'h1, _0384_ } : 2'h2;
  assign _0386_ = _0383_ ? _0385_ : 2'h0;
  assign _0387_ = $signed(32'd4) < $signed({ 28'h0000000, r2[171:168] });
  assign _0388_ = ~ r2[301];
  assign _0389_ = r2[207] ? { 1'h1, _0388_ } : 2'h2;
  assign _0390_ = _0387_ ? _0389_ : 2'h0;
  assign _0391_ = $signed(32'd5) < $signed({ 28'h0000000, r2[171:168] });
  assign _0392_ = ~ r2[302];
  assign _0393_ = r2[207] ? { 1'h1, _0392_ } : 2'h2;
  assign _0394_ = _0391_ ? _0393_ : 2'h0;
  assign _0395_ = $signed(32'd6) < $signed({ 28'h0000000, r2[171:168] });
  assign _0396_ = ~ r2[303];
  assign _0397_ = r2[207] ? { 1'h1, _0396_ } : 2'h2;
  assign _0398_ = _0395_ ? _0397_ : 2'h0;
  assign _0399_ = $signed(32'd7) < $signed({ 28'h0000000, r2[171:168] });
  assign _0400_ = ~ r2[304];
  assign _0401_ = r2[207] ? { 1'h1, _0400_ } : 2'h2;
  assign _0402_ = _0399_ ? _0401_ : 2'h0;
  assign _0403_ = _0374_ == 2'h3;
  assign _0404_ = _0374_ == 2'h2;
  assign _0405_ = _0370_ & r2[180];
  assign _0406_ = _0370_ & r2[180];
  assign _0407_ = _0370_ & r2[180];
  assign _0408_ = _0370_ & r2[180];
  assign _0409_ = _0370_ & r2[180];
  assign _0410_ = _0370_ & r2[180];
  assign _0411_ = _0370_ & r2[180];
  assign _0412_ = _0370_ & r2[180];
  function [7:0] \20827 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \20827  = b[7:0];
      2'b1?:
        \20827  = b[15:8];
      default:
        \20827  = a;
    endcase
  endfunction
  assign _0413_ = \20827 ({ _0405_, _0406_, _0407_, _0408_, _0409_, _0410_, _0411_, _0412_ }, { _0983_, r3[92:85] }, { _0404_, _0403_ });
  assign _0414_ = _0378_ == 2'h3;
  assign _0415_ = _0378_ == 2'h2;
  assign _0416_ = _0370_ & r2[180];
  assign _0417_ = _0370_ & r2[180];
  assign _0418_ = _0370_ & r2[180];
  assign _0419_ = _0370_ & r2[180];
  assign _0420_ = _0370_ & r2[180];
  assign _0421_ = _0370_ & r2[180];
  assign _0422_ = _0370_ & r2[180];
  assign _0423_ = _0370_ & r2[180];
  function [7:0] \20865 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \20865  = b[7:0];
      2'b1?:
        \20865  = b[15:8];
      default:
        \20865  = a;
    endcase
  endfunction
  assign _0424_ = \20865 ({ _0416_, _0417_, _0418_, _0419_, _0420_, _0421_, _0422_, _0423_ }, { _0986_, r3[100:93] }, { _0415_, _0414_ });
  assign _0425_ = _0382_ == 2'h3;
  assign _0426_ = _0382_ == 2'h2;
  assign _0427_ = _0370_ & r2[180];
  assign _0428_ = _0370_ & r2[180];
  assign _0429_ = _0370_ & r2[180];
  assign _0430_ = _0370_ & r2[180];
  assign _0431_ = _0370_ & r2[180];
  assign _0432_ = _0370_ & r2[180];
  assign _0433_ = _0370_ & r2[180];
  assign _0434_ = _0370_ & r2[180];
  function [7:0] \20903 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \20903  = b[7:0];
      2'b1?:
        \20903  = b[15:8];
      default:
        \20903  = a;
    endcase
  endfunction
  assign _0435_ = \20903 ({ _0427_, _0428_, _0429_, _0430_, _0431_, _0432_, _0433_, _0434_ }, { _0989_, r3[108:101] }, { _0426_, _0425_ });
  assign _0436_ = _0386_ == 2'h3;
  assign _0437_ = _0386_ == 2'h2;
  assign _0438_ = _0370_ & r2[180];
  assign _0439_ = _0370_ & r2[180];
  assign _0440_ = _0370_ & r2[180];
  assign _0441_ = _0370_ & r2[180];
  assign _0442_ = _0370_ & r2[180];
  assign _0443_ = _0370_ & r2[180];
  assign _0444_ = _0370_ & r2[180];
  assign _0445_ = _0370_ & r2[180];
  function [7:0] \20941 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \20941  = b[7:0];
      2'b1?:
        \20941  = b[15:8];
      default:
        \20941  = a;
    endcase
  endfunction
  assign _0446_ = \20941 ({ _0438_, _0439_, _0440_, _0441_, _0442_, _0443_, _0444_, _0445_ }, { _0992_, r3[116:109] }, { _0437_, _0436_ });
  assign _0447_ = _0390_ == 2'h3;
  assign _0448_ = _0390_ == 2'h2;
  assign _0449_ = _0370_ & r2[180];
  assign _0450_ = _0370_ & r2[180];
  assign _0451_ = _0370_ & r2[180];
  assign _0452_ = _0370_ & r2[180];
  assign _0453_ = _0370_ & r2[180];
  assign _0454_ = _0370_ & r2[180];
  assign _0455_ = _0370_ & r2[180];
  assign _0456_ = _0370_ & r2[180];
  function [7:0] \20979 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \20979  = b[7:0];
      2'b1?:
        \20979  = b[15:8];
      default:
        \20979  = a;
    endcase
  endfunction
  assign _0457_ = \20979 ({ _0449_, _0450_, _0451_, _0452_, _0453_, _0454_, _0455_, _0456_ }, { _0995_, r3[124:117] }, { _0448_, _0447_ });
  assign _0458_ = _0394_ == 2'h3;
  assign _0459_ = _0394_ == 2'h2;
  assign _0460_ = _0370_ & r2[180];
  assign _0461_ = _0370_ & r2[180];
  assign _0462_ = _0370_ & r2[180];
  assign _0463_ = _0370_ & r2[180];
  assign _0464_ = _0370_ & r2[180];
  assign _0465_ = _0370_ & r2[180];
  assign _0466_ = _0370_ & r2[180];
  assign _0467_ = _0370_ & r2[180];
  function [7:0] \21017 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \21017  = b[7:0];
      2'b1?:
        \21017  = b[15:8];
      default:
        \21017  = a;
    endcase
  endfunction
  assign _0468_ = \21017 ({ _0460_, _0461_, _0462_, _0463_, _0464_, _0465_, _0466_, _0467_ }, { _0998_, r3[132:125] }, { _0459_, _0458_ });
  assign _0469_ = _0398_ == 2'h3;
  assign _0470_ = _0398_ == 2'h2;
  assign _0471_ = _0370_ & r2[180];
  assign _0472_ = _0370_ & r2[180];
  assign _0473_ = _0370_ & r2[180];
  assign _0474_ = _0370_ & r2[180];
  assign _0475_ = _0370_ & r2[180];
  assign _0476_ = _0370_ & r2[180];
  assign _0477_ = _0370_ & r2[180];
  assign _0478_ = _0370_ & r2[180];
  function [7:0] \21055 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \21055  = b[7:0];
      2'b1?:
        \21055  = b[15:8];
      default:
        \21055  = a;
    endcase
  endfunction
  assign _0479_ = \21055 ({ _0471_, _0472_, _0473_, _0474_, _0475_, _0476_, _0477_, _0478_ }, { _1001_, r3[140:133] }, { _0470_, _0469_ });
  assign _0480_ = _0402_ == 2'h3;
  assign _0481_ = _0402_ == 2'h2;
  assign _0482_ = _0370_ & r2[180];
  assign _0483_ = _0370_ & r2[180];
  assign _0484_ = _0370_ & r2[180];
  assign _0485_ = _0370_ & r2[180];
  assign _0486_ = _0370_ & r2[180];
  assign _0487_ = _0370_ & r2[180];
  assign _0488_ = _0370_ & r2[180];
  assign _0489_ = _0370_ & r2[180];
  function [7:0] \21093 ;
    input [7:0] a;
    input [15:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \21093  = b[7:0];
      2'b1?:
        \21093  = b[15:8];
      default:
        \21093  = a;
    endcase
  endfunction
  assign _0490_ = \21093 ({ _0482_, _0483_, _0484_, _0485_, _0486_, _0487_, _0488_, _0489_ }, { _1004_, r3[148:141] }, { _0481_, _0480_ });
  assign _0491_ = | { _0435_[6:0], _0424_, _0413_ };
  assign _0492_ = - $signed({ _0413_[0], _0413_[1], _0413_[2], _0413_[3], _0413_[4], _0413_[5], _0413_[6], _0413_[7], _0424_[0], _0424_[1], _0424_[2], _0424_[3], _0424_[4], _0424_[5], _0424_[6], _0424_[7], _0435_[0], _0435_[1], _0435_[2], _0435_[3], _0435_[4], _0435_[5], _0435_[6] });
  assign _0493_ = _0492_ & { _0413_[0], _0413_[1], _0413_[2], _0413_[3], _0413_[4], _0413_[5], _0413_[6], _0413_[7], _0424_[0], _0424_[1], _0424_[2], _0424_[3], _0424_[4], _0424_[5], _0424_[6], _0424_[7], _0435_[0], _0435_[1], _0435_[2], _0435_[3], _0435_[4], _0435_[5], _0435_[6] };
  assign _0494_ = _0492_ | { _0413_[0], _0413_[1], _0413_[2], _0413_[3], _0413_[4], _0413_[5], _0413_[6], _0413_[7], _0424_[0], _0424_[1], _0424_[2], _0424_[3], _0424_[4], _0424_[5], _0424_[6], _0424_[7], _0435_[0], _0435_[1], _0435_[2], _0435_[3], _0435_[4], _0435_[5], _0435_[6] };
  assign _0495_ = ~ _0494_[0];
  assign _0496_ = _0494_[1] & _0495_;
  assign _0497_ = 1'h0 | _0496_;
  assign _0498_ = ~ _0494_[2];
  assign _0499_ = _0494_[3] & _0498_;
  assign _0500_ = _0497_ | _0499_;
  assign _0501_ = ~ _0494_[4];
  assign _0502_ = _0494_[5] & _0501_;
  assign _0503_ = _0500_ | _0502_;
  assign _0504_ = ~ _0494_[6];
  assign _0505_ = _0494_[7] & _0504_;
  assign _0506_ = _0503_ | _0505_;
  assign _0507_ = ~ _0494_[8];
  assign _0508_ = _0494_[9] & _0507_;
  assign _0509_ = _0506_ | _0508_;
  assign _0510_ = ~ _0494_[10];
  assign _0511_ = _0494_[11] & _0510_;
  assign _0512_ = _0509_ | _0511_;
  assign _0513_ = ~ _0494_[12];
  assign _0514_ = _0494_[13] & _0513_;
  assign _0515_ = _0512_ | _0514_;
  assign _0516_ = ~ _0494_[14];
  assign _0517_ = _0494_[15] & _0516_;
  assign _0518_ = _0515_ | _0517_;
  assign _0519_ = ~ _0494_[16];
  assign _0520_ = _0494_[17] & _0519_;
  assign _0521_ = _0518_ | _0520_;
  assign _0522_ = ~ _0494_[18];
  assign _0523_ = _0494_[19] & _0522_;
  assign _0524_ = _0521_ | _0523_;
  assign _0525_ = ~ _0494_[20];
  assign _0526_ = _0494_[21] & _0525_;
  assign _0527_ = _0524_ | _0526_;
  assign _0528_ = ~ _0494_[22];
  assign _0529_ = _0494_[22] & _0528_;
  assign _0530_ = _0527_ | _0529_;
  assign _0531_ = ~ _0494_[22];
  assign _0532_ = _0494_[22] & _0531_;
  assign _0533_ = _0530_ | _0532_;
  assign _0534_ = ~ _0494_[22];
  assign _0535_ = _0494_[22] & _0534_;
  assign _0536_ = _0533_ | _0535_;
  assign _0537_ = ~ _0494_[22];
  assign _0538_ = _0494_[22] & _0537_;
  assign _0539_ = _0536_ | _0538_;
  assign _0540_ = ~ _0494_[22];
  assign _0541_ = _0494_[22] & _0540_;
  assign _0542_ = _0539_ | _0541_;
  assign _0543_ = ~ _0494_[22];
  assign _0544_ = _0494_[22] & _0543_;
  assign _0545_ = _0542_ | _0544_;
  assign _0546_ = ~ _0494_[22];
  assign _0547_ = _0494_[22] & _0546_;
  assign _0548_ = _0545_ | _0547_;
  assign _0549_ = ~ _0494_[22];
  assign _0550_ = _0494_[22] & _0549_;
  assign _0551_ = _0548_ | _0550_;
  assign _0552_ = ~ _0494_[22];
  assign _0553_ = _0494_[22] & _0552_;
  assign _0554_ = _0551_ | _0553_;
  assign _0555_ = ~ _0494_[22];
  assign _0556_ = _0494_[22] & _0555_;
  assign _0557_ = _0554_ | _0556_;
  assign _0558_ = ~ _0494_[22];
  assign _0559_ = _0494_[22] & _0558_;
  assign _0560_ = _0557_ | _0559_;
  assign _0561_ = ~ _0494_[22];
  assign _0562_ = _0494_[22] & _0561_;
  assign _0563_ = _0560_ | _0562_;
  assign _0564_ = ~ _0494_[22];
  assign _0565_ = _0494_[22] & _0564_;
  assign _0566_ = _0563_ | _0565_;
  assign _0567_ = ~ _0494_[22];
  assign _0568_ = _0494_[22] & _0567_;
  assign _0569_ = _0566_ | _0568_;
  assign _0570_ = ~ _0494_[22];
  assign _0571_ = _0494_[22] & _0570_;
  assign _0572_ = _0569_ | _0571_;
  assign _0573_ = ~ _0494_[22];
  assign _0574_ = _0494_[22] & _0573_;
  assign _0575_ = _0572_ | _0574_;
  assign _0576_ = ~ _0494_[22];
  assign _0577_ = _0494_[22] & _0576_;
  assign _0578_ = _0575_ | _0577_;
  assign _0579_ = ~ _0494_[22];
  assign _0580_ = _0494_[22] & _0579_;
  assign _0581_ = _0578_ | _0580_;
  assign _0582_ = ~ _0494_[22];
  assign _0583_ = _0494_[22] & _0582_;
  assign _0584_ = _0581_ | _0583_;
  assign _0585_ = ~ _0494_[22];
  assign _0586_ = _0494_[22] & _0585_;
  assign _0587_ = _0584_ | _0586_;
  assign _0588_ = ~ _0494_[22];
  assign _0589_ = _0494_[22] & _0588_;
  assign _0590_ = _0587_ | _0589_;
  assign _0591_ = ~ _0494_[1];
  assign _0592_ = _0494_[3] & _0591_;
  assign _0593_ = 1'h0 | _0592_;
  assign _0594_ = ~ _0494_[5];
  assign _0595_ = _0494_[7] & _0594_;
  assign _0596_ = _0593_ | _0595_;
  assign _0597_ = ~ _0494_[9];
  assign _0598_ = _0494_[11] & _0597_;
  assign _0599_ = _0596_ | _0598_;
  assign _0600_ = ~ _0494_[13];
  assign _0601_ = _0494_[15] & _0600_;
  assign _0602_ = _0599_ | _0601_;
  assign _0603_ = ~ _0494_[17];
  assign _0604_ = _0494_[19] & _0603_;
  assign _0605_ = _0602_ | _0604_;
  assign _0606_ = ~ _0494_[21];
  assign _0607_ = _0494_[22] & _0606_;
  assign _0608_ = _0605_ | _0607_;
  assign _0609_ = ~ _0494_[22];
  assign _0610_ = _0494_[22] & _0609_;
  assign _0611_ = _0608_ | _0610_;
  assign _0612_ = ~ _0494_[22];
  assign _0613_ = _0494_[22] & _0612_;
  assign _0614_ = _0611_ | _0613_;
  assign _0615_ = ~ _0494_[22];
  assign _0616_ = _0494_[22] & _0615_;
  assign _0617_ = _0614_ | _0616_;
  assign _0618_ = ~ _0494_[22];
  assign _0619_ = _0494_[22] & _0618_;
  assign _0620_ = _0617_ | _0619_;
  assign _0621_ = ~ _0494_[22];
  assign _0622_ = _0494_[22] & _0621_;
  assign _0623_ = _0620_ | _0622_;
  assign _0624_ = ~ _0494_[22];
  assign _0625_ = _0494_[22] & _0624_;
  assign _0626_ = _0623_ | _0625_;
  assign _0627_ = ~ _0494_[22];
  assign _0628_ = _0494_[22] & _0627_;
  assign _0629_ = _0626_ | _0628_;
  assign _0630_ = ~ _0494_[22];
  assign _0631_ = _0494_[22] & _0630_;
  assign _0632_ = _0629_ | _0631_;
  assign _0633_ = ~ _0494_[22];
  assign _0634_ = _0494_[22] & _0633_;
  assign _0635_ = _0632_ | _0634_;
  assign _0636_ = ~ _0494_[22];
  assign _0637_ = _0494_[22] & _0636_;
  assign _0638_ = _0635_ | _0637_;
  assign _0639_ = ~ _0494_[3];
  assign _0640_ = _0494_[7] & _0639_;
  assign _0641_ = 1'h0 | _0640_;
  assign _0642_ = ~ _0494_[11];
  assign _0643_ = _0494_[15] & _0642_;
  assign _0644_ = _0641_ | _0643_;
  assign _0645_ = ~ _0494_[19];
  assign _0646_ = _0494_[22] & _0645_;
  assign _0647_ = _0644_ | _0646_;
  assign _0648_ = ~ _0494_[22];
  assign _0649_ = _0494_[22] & _0648_;
  assign _0650_ = _0647_ | _0649_;
  assign _0651_ = ~ _0494_[22];
  assign _0652_ = _0494_[22] & _0651_;
  assign _0653_ = _0650_ | _0652_;
  assign _0654_ = ~ _0494_[22];
  assign _0655_ = _0494_[22] & _0654_;
  assign _0656_ = _0653_ | _0655_;
  assign _0657_ = ~ _0494_[22];
  assign _0658_ = _0494_[22] & _0657_;
  assign _0659_ = _0656_ | _0658_;
  assign _0660_ = ~ _0494_[22];
  assign _0661_ = _0494_[22] & _0660_;
  assign _0662_ = _0659_ | _0661_;
  assign _0663_ = ~ _0494_[7];
  assign _0664_ = _0494_[15] & _0663_;
  assign _0665_ = 1'h0 | _0664_;
  assign _0666_ = ~ _0494_[22];
  assign _0667_ = _0494_[22] & _0666_;
  assign _0668_ = _0665_ | _0667_;
  assign _0669_ = ~ _0494_[22];
  assign _0670_ = _0494_[22] & _0669_;
  assign _0671_ = _0668_ | _0670_;
  assign _0672_ = ~ _0494_[22];
  assign _0673_ = _0494_[22] & _0672_;
  assign _0674_ = _0671_ | _0673_;
  assign _0675_ = ~ _0494_[15];
  assign _0676_ = _0494_[22] & _0675_;
  assign _0677_ = 1'h0 | _0676_;
  assign _0678_ = ~ _0494_[22];
  assign _0679_ = _0494_[22] & _0678_;
  assign _0680_ = _0677_ | _0679_;
  assign _0681_ = ~ _0494_[22];
  assign _0682_ = _0494_[22] & _0681_;
  assign _0683_ = 1'h0 | _0682_;
  assign _0684_ = | _0493_[1];
  assign _0685_ = 1'h0 | _0684_;
  assign _0686_ = | _0493_[3];
  assign _0687_ = _0685_ | _0686_;
  assign _0688_ = | _0493_[5];
  assign _0689_ = _0687_ | _0688_;
  assign _0690_ = | _0493_[7];
  assign _0691_ = _0689_ | _0690_;
  assign _0692_ = | _0493_[9];
  assign _0693_ = _0691_ | _0692_;
  assign _0694_ = | _0493_[11];
  assign _0695_ = _0693_ | _0694_;
  assign _0696_ = | _0493_[13];
  assign _0697_ = _0695_ | _0696_;
  assign _0698_ = | _0493_[15];
  assign _0699_ = _0697_ | _0698_;
  assign _0700_ = | _0493_[17];
  assign _0701_ = _0699_ | _0700_;
  assign _0702_ = | _0493_[19];
  assign _0703_ = _0701_ | _0702_;
  assign _0704_ = | _0493_[21];
  assign _0705_ = _0703_ | _0704_;
  assign _0706_ = | 1'h0;
  assign _0707_ = _0705_ | _0706_;
  assign _0708_ = | 1'h0;
  assign _0709_ = _0707_ | _0708_;
  assign _0710_ = | 1'h0;
  assign _0711_ = _0709_ | _0710_;
  assign _0712_ = | 1'h0;
  assign _0713_ = _0711_ | _0712_;
  assign _0714_ = | 1'h0;
  assign _0715_ = _0713_ | _0714_;
  assign _0716_ = | 1'h0;
  assign _0717_ = _0715_ | _0716_;
  assign _0718_ = | 1'h0;
  assign _0719_ = _0717_ | _0718_;
  assign _0720_ = | 1'h0;
  assign _0721_ = _0719_ | _0720_;
  assign _0722_ = | 1'h0;
  assign _0723_ = _0721_ | _0722_;
  assign _0724_ = | 1'h0;
  assign _0725_ = _0723_ | _0724_;
  assign _0726_ = | 1'h0;
  assign _0727_ = _0725_ | _0726_;
  assign _0728_ = | 1'h0;
  assign _0729_ = _0727_ | _0728_;
  assign _0730_ = | 1'h0;
  assign _0731_ = _0729_ | _0730_;
  assign _0732_ = | 1'h0;
  assign _0733_ = _0731_ | _0732_;
  assign _0734_ = | 1'h0;
  assign _0735_ = _0733_ | _0734_;
  assign _0736_ = | 1'h0;
  assign _0737_ = _0735_ | _0736_;
  assign _0738_ = | 1'h0;
  assign _0739_ = _0737_ | _0738_;
  assign _0740_ = | 1'h0;
  assign _0741_ = _0739_ | _0740_;
  assign _0742_ = | 1'h0;
  assign _0743_ = _0741_ | _0742_;
  assign _0744_ = | 1'h0;
  assign _0745_ = _0743_ | _0744_;
  assign _0746_ = | 1'h0;
  assign _0747_ = _0745_ | _0746_;
  assign _0748_ = | _0493_[3:2];
  assign _0749_ = 1'h0 | _0748_;
  assign _0750_ = | _0493_[7:6];
  assign _0751_ = _0749_ | _0750_;
  assign _0752_ = | _0493_[11:10];
  assign _0753_ = _0751_ | _0752_;
  assign _0754_ = | _0493_[15:14];
  assign _0755_ = _0753_ | _0754_;
  assign _0756_ = | _0493_[19:18];
  assign _0757_ = _0755_ | _0756_;
  assign _0758_ = | { 1'h0, _0493_[22] };
  assign _0759_ = _0757_ | _0758_;
  assign _0760_ = | 2'h0;
  assign _0761_ = _0759_ | _0760_;
  assign _0762_ = | 2'h0;
  assign _0763_ = _0761_ | _0762_;
  assign _0764_ = | 2'h0;
  assign _0765_ = _0763_ | _0764_;
  assign _0766_ = | 2'h0;
  assign _0767_ = _0765_ | _0766_;
  assign _0768_ = | 2'h0;
  assign _0769_ = _0767_ | _0768_;
  assign _0770_ = | 2'h0;
  assign _0771_ = _0769_ | _0770_;
  assign _0772_ = | 2'h0;
  assign _0773_ = _0771_ | _0772_;
  assign _0774_ = | 2'h0;
  assign _0775_ = _0773_ | _0774_;
  assign _0776_ = | 2'h0;
  assign _0777_ = _0775_ | _0776_;
  assign _0778_ = | 2'h0;
  assign _0779_ = _0777_ | _0778_;
  assign _0780_ = | _0493_[7:4];
  assign _0781_ = 1'h0 | _0780_;
  assign _0782_ = | _0493_[15:12];
  assign _0783_ = _0781_ | _0782_;
  assign _0784_ = | { 1'h0, _0493_[22:20] };
  assign _0785_ = _0783_ | _0784_;
  assign _0786_ = | 4'h0;
  assign _0787_ = _0785_ | _0786_;
  assign _0788_ = | 4'h0;
  assign _0789_ = _0787_ | _0788_;
  assign _0790_ = | 4'h0;
  assign _0791_ = _0789_ | _0790_;
  assign _0792_ = | 4'h0;
  assign _0793_ = _0791_ | _0792_;
  assign _0794_ = | 4'h0;
  assign _0795_ = _0793_ | _0794_;
  assign _0796_ = | _0493_[15:8];
  assign _0797_ = 1'h0 | _0796_;
  assign _0798_ = | 8'h00;
  assign _0799_ = _0797_ | _0798_;
  assign _0800_ = | 8'h00;
  assign _0801_ = _0799_ | _0800_;
  assign _0802_ = | 8'h00;
  assign _0803_ = _0801_ | _0802_;
  assign _0804_ = | { 9'h000, _0493_[22:16] };
  assign _0805_ = 1'h0 | _0804_;
  assign _0806_ = | 16'h0000;
  assign _0807_ = _0805_ | _0806_;
  assign _0808_ = | 32'd0;
  assign _0809_ = 1'h0 | _0808_;
  assign _0810_ = \d_in.valid  & r2[2];
  assign _0811_ = _0810_ ? { _1004_, _1001_, _0998_, _0995_, _0992_, _0989_, _0986_, _0983_ } : r3[148:85];
  assign _0812_ = ~ r2[203];
  assign _0813_ = ~ r2[200];
  assign _0814_ = _0812_ & _0813_;
  assign _0815_ = ~ r2[195];
  assign _0816_ = _0815_ ? { 32'h00000000, r3[244:213] } : r3[212:149];
  assign _0817_ = _0814_ ? _0816_ : \m_in.sprval ;
  assign _0818_ = r2[6] ? 1'h1 : 1'h0;
  assign _0819_ = r2[6] ? _0817_ : 64'h0000000000000000;
  assign _0820_ = r2[206] ? 1'h1 : 1'h0;
  assign _0821_ = r2[10] ? 1'h1 : _0818_;
  assign _0822_ = r2[11] ? 1'h1 : 1'h0;
  assign _0823_ = r2[0] ? _0821_ : 1'h0;
  assign _0824_ = r2[0] ? _0822_ : 1'h0;
  assign _0825_ = r2[0] ? _0820_ : 1'h0;
  assign _0826_ = r2[0] ? _0819_ : 64'h0000000000000000;
  assign _0827_ = ~ r2[208];
  assign _0828_ = _0827_ | r2[207];
  assign _0829_ = ~ r2[194];
  assign _0830_ = r2[2] & _0829_;
  assign _0831_ = 1'h1 & r2[194];
  assign _0832_ = r2[181] & r2[3];
  assign _0833_ = _0841_ ? 2'h3 : r3[1:0];
  assign _0834_ = _0842_ ? 1'h1 : 1'h0;
  assign _0835_ = _0831_ ? _0824_ : _0832_;
  assign _0836_ = _0828_ & _0831_;
  assign _0837_ = _0828_ & _0831_;
  assign _0838_ = _0843_ ? _0830_ : _0823_;
  assign _0839_ = _0844_ ? _0835_ : _0824_;
  assign _0840_ = _0828_ ? 1'h0 : 1'h1;
  assign _0841_ = \d_in.valid  & _0836_;
  assign _0842_ = \d_in.valid  & _0837_;
  assign _0843_ = \d_in.valid  & _0828_;
  assign _0844_ = \d_in.valid  & _0828_;
  assign _0845_ = \d_in.valid  ? _0840_ : 1'h0;
  assign _0846_ = ~ r2[2];
  assign _0847_ = \d_in.cache_paradox  ? _0833_ : 2'h1;
  assign _0848_ = \d_in.cache_paradox  ? r3[284] : 1'h0;
  assign _0849_ = \d_in.cache_paradox  ? 1'h0 : 1'h1;
  assign _0850_ = _0856_ ? 1'h1 : _0825_;
  assign _0851_ = \d_in.cache_paradox  ? _0846_ : 1'h0;
  assign _0852_ = \d_in.cache_paradox  ? \d_in.cache_paradox  : 1'h0;
  assign _0853_ = \d_in.error  ? _0847_ : _0833_;
  assign _0854_ = \d_in.error  ? _0848_ : r3[284];
  assign _0855_ = \d_in.error  ? _0849_ : 1'h0;
  assign _0856_ = \d_in.error  & \d_in.cache_paradox ;
  assign _0857_ = \d_in.error  ? _0851_ : 1'h0;
  assign _0858_ = \d_in.error  ? _0852_ : 1'h0;
  assign _0859_ = ~ r2[7];
  assign _0860_ = r2[9] ? 2'h1 : 2'h2;
  assign _0861_ = _0873_ ? 1'h1 : 1'h0;
  assign _0862_ = ~ r2[195];
  assign _0863_ = _0862_ ? r3[212:149] : r2[157:94];
  assign _0864_ = _0862_ ? r2[125:94] : r3[244:213];
  assign _0865_ = r2[7] ? { _0864_, _0863_ } : r3[244:149];
  assign _0866_ = _0871_ ? _0860_ : _0853_;
  assign _0867_ = r2[8] ? r3[244:149] : _0865_;
  assign _0868_ = r2[8] & r2[9];
  assign _0869_ = _0874_ ? _0859_ : _0855_;
  assign _0870_ = r2[8] ? r2[7] : 1'h0;
  assign _0871_ = r2[0] & r2[8];
  assign _0872_ = r2[0] ? _0867_ : r3[244:149];
  assign _0873_ = r2[0] & _0868_;
  assign _0874_ = r2[0] & r2[8];
  assign _0875_ = r2[0] ? _0870_ : 1'h0;
  assign _0876_ = r3[1:0] == 2'h0;
  assign _0877_ = ~ r2[9];
  assign _0878_ = _0881_ ? 2'h0 : r3[1:0];
  assign _0879_ = _0882_ ? 1'h1 : r3[284];
  assign _0880_ = _0877_ ? 1'h1 : 1'h0;
  assign _0881_ = \m_in.done  & _0877_;
  assign _0882_ = \m_in.done  & _0877_;
  assign _0883_ = \m_in.done  ? _0880_ : 1'h0;
  assign _0884_ = r2[3] | r2[5];
  assign _0885_ = \m_in.err  ? 1'h1 : _0825_;
  assign _0886_ = \m_in.err  ? { \m_in.badtree , \m_in.rc_error  } : 2'h0;
  assign _0887_ = \m_in.err  ? _0884_ : 1'h0;
  assign _0888_ = \m_in.err  ? \m_in.perm_error  : 1'h0;
  assign _0889_ = \m_in.err  ? \m_in.invalid  : 1'h0;
  assign _0890_ = r3[1:0] == 2'h1;
  assign _0891_ = r3[1:0] == 2'h2;
  assign _0892_ = r3[1:0] == 2'h3;
  function [1:0] \21976 ;
    input [1:0] a;
    input [7:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \21976  = b[1:0];
      4'b??1?:
        \21976  = b[3:2];
      4'b?1??:
        \21976  = b[5:4];
      4'b1???:
        \21976  = b[7:6];
      default:
        \21976  = a;
    endcase
  endfunction
  assign _0893_ = \21976 (2'hx, { r3[1:0], r3[1:0], _0878_, _0866_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \21978 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \21978  = b[0:0];
      4'b??1?:
        \21978  = b[1:1];
      4'b?1??:
        \21978  = b[2:2];
      4'b1???:
        \21978  = b[3:3];
      default:
        \21978  = a;
    endcase
  endfunction
  assign _0894_ = \21978 (1'hx, { 3'h0, _0834_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [95:0] \21980 ;
    input [95:0] a;
    input [383:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \21980  = b[95:0];
      4'b??1?:
        \21980  = b[191:96];
      4'b?1??:
        \21980  = b[287:192];
      4'b1???:
        \21980  = b[383:288];
      default:
        \21980  = a;
    endcase
  endfunction
  assign _0895_ = \21980 (96'hxxxxxxxxxxxxxxxxxxxxxxxx, { r3[244:149], r3[244:149], r3[244:149], _0872_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \21983 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \21983  = b[0:0];
      4'b??1?:
        \21983  = b[1:1];
      4'b?1??:
        \21983  = b[2:2];
      4'b1???:
        \21983  = b[3:3];
      default:
        \21983  = a;
    endcase
  endfunction
  assign _0896_ = \21983 (1'hx, { r3[284], r3[284], _0879_, _0854_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \21986 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \21986  = b[0:0];
      4'b??1?:
        \21986  = b[1:1];
      4'b?1??:
        \21986  = b[2:2];
      4'b1???:
        \21986  = b[3:3];
      default:
        \21986  = a;
    endcase
  endfunction
  assign _0897_ = \21986 (1'hx, { 3'h0, _0861_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \21992 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \21992  = b[0:0];
      4'b??1?:
        \21992  = b[1:1];
      4'b?1??:
        \21992  = b[2:2];
      4'b1???:
        \21992  = b[3:3];
      default:
        \21992  = a;
    endcase
  endfunction
  assign _0898_ = \21992 (1'hx, { 2'h0, _0883_, 1'h0 }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \21996 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \21996  = b[0:0];
      4'b??1?:
        \21996  = b[1:1];
      4'b?1??:
        \21996  = b[2:2];
      4'b1???:
        \21996  = b[3:3];
      default:
        \21996  = a;
    endcase
  endfunction
  assign _0899_ = \21996 (1'hx, { 3'h0, _0869_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22000 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22000  = b[0:0];
      4'b??1?:
        \22000  = b[1:1];
      4'b?1??:
        \22000  = b[2:2];
      4'b1???:
        \22000  = b[3:3];
      default:
        \22000  = a;
    endcase
  endfunction
  assign _0900_ = \22000 (1'hx, { 3'h0, _0875_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22004 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22004  = b[0:0];
      4'b??1?:
        \22004  = b[1:1];
      4'b?1??:
        \22004  = b[2:2];
      4'b1???:
        \22004  = b[3:3];
      default:
        \22004  = a;
    endcase
  endfunction
  assign _0901_ = \22004 (1'hx, { 1'h1, _0823_, _0823_, _0838_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22006 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22006  = b[0:0];
      4'b??1?:
        \22006  = b[1:1];
      4'b?1??:
        \22006  = b[2:2];
      4'b1???:
        \22006  = b[3:3];
      default:
        \22006  = a;
    endcase
  endfunction
  assign _0902_ = \22006 (1'hx, { _0824_, _0824_, _0824_, _0839_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22009 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22009  = b[0:0];
      4'b??1?:
        \22009  = b[1:1];
      4'b?1??:
        \22009  = b[2:2];
      4'b1???:
        \22009  = b[3:3];
      default:
        \22009  = a;
    endcase
  endfunction
  assign _0903_ = \22009 (1'hx, { 3'h0, _0845_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22012 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22012  = b[0:0];
      4'b??1?:
        \22012  = b[1:1];
      4'b?1??:
        \22012  = b[2:2];
      4'b1???:
        \22012  = b[3:3];
      default:
        \22012  = a;
    endcase
  endfunction
  assign _0904_ = \22012 (1'hx, { _0825_, _0825_, _0885_, _0850_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [1:0] \22015 ;
    input [1:0] a;
    input [7:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22015  = b[1:0];
      4'b??1?:
        \22015  = b[3:2];
      4'b?1??:
        \22015  = b[5:4];
      4'b1???:
        \22015  = b[7:6];
      default:
        \22015  = a;
    endcase
  endfunction
  assign _0905_ = \22015 (2'hx, { 4'h0, _0886_, 2'h0 }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22018 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22018  = b[0:0];
      4'b??1?:
        \22018  = b[1:1];
      4'b?1??:
        \22018  = b[2:2];
      4'b1???:
        \22018  = b[3:3];
      default:
        \22018  = a;
    endcase
  endfunction
  assign _0906_ = \22018 (1'hx, { 2'h0, _0887_, _0857_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22021 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22021  = b[0:0];
      4'b??1?:
        \22021  = b[1:1];
      4'b?1??:
        \22021  = b[2:2];
      4'b1???:
        \22021  = b[3:3];
      default:
        \22021  = a;
    endcase
  endfunction
  assign _0907_ = \22021 (1'hx, { 2'h0, _0888_, 1'h0 }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22024 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22024  = b[0:0];
      4'b??1?:
        \22024  = b[1:1];
      4'b?1??:
        \22024  = b[2:2];
      4'b1???:
        \22024  = b[3:3];
      default:
        \22024  = a;
    endcase
  endfunction
  assign _0908_ = \22024 (1'hx, { 3'h0, _0858_ }, { _0892_, _0891_, _0890_, _0876_ });
  function [0:0] \22027 ;
    input [0:0] a;
    input [3:0] b;
    input [3:0] s;
    (* parallel_case *)
    casez (s)
      4'b???1:
        \22027  = b[0:0];
      4'b??1?:
        \22027  = b[1:1];
      4'b?1??:
        \22027  = b[2:2];
      4'b1???:
        \22027  = b[3:3];
      default:
        \22027  = a;
    endcase
  endfunction
  assign _0909_ = \22027 (1'hx, { 2'h0, _0889_, 1'h0 }, { _0892_, _0891_, _0890_, _0876_ });
  assign _0910_ = complete | _0904_;
  assign _0911_ = _0910_ ? 2'h0 : _0893_;
  assign _0912_ = _0910_ ? 1'h1 : _0896_;
  assign _0913_ = r2[2] & complete;
  assign _0914_ = r2[3] | r2[5];
  assign _0915_ = _0914_ & complete;
  assign _0916_ = ~ r2[9];
  assign _0917_ = ~ \m_in.segerr ;
  assign _0918_ = _0917_ ? { 1'h0, _0909_, 1'h0, _0908_, _0907_, 1'h0, _0906_, 5'h00, _0905_, 18'h00000 } : _0895_[95:64];
  assign _0919_ = _0917_ ? 12'h300 : 12'h380;
  assign _0920_ = ~ \m_in.segerr ;
  assign _0921_ = _0920_ ? 12'h400 : 12'h480;
  assign _0922_ = _0920_ ? { \m_in.badtree , \m_in.rc_error  } : 2'h0;
  assign _0923_ = _0920_ ? \m_in.perm_error  : 1'h0;
  assign _0924_ = _0920_ ? \m_in.invalid  : 1'h0;
  assign _0925_ = _0916_ ? { _0918_, r2[77:14] } : _0895_;
  assign _0926_ = _0916_ ? _0919_ : _0921_;
  assign _0927_ = _0916_ ? 2'h0 : _0922_;
  assign _0928_ = _0916_ ? 1'h0 : _0923_;
  assign _0929_ = _0916_ ? 1'h0 : _0924_;
  assign _0930_ = r2[206] ? r2[77:14] : _0925_[63:0];
  assign _0931_ = r2[206] ? _0895_[95:64] : _0925_[95:64];
  assign _0932_ = r2[206] ? 12'h600 : _0926_;
  assign _0933_ = r2[206] ? 2'h0 : _0927_;
  assign _0934_ = r2[206] ? 1'h0 : _0928_;
  assign _0935_ = r2[206] ? 1'h0 : _0929_;
  assign _0936_ = _0904_ ? { _0931_, _0930_ } : _0895_;
  assign _0937_ = _0904_ ? { r2[272:209], _0932_ } : r3[361:286];
  assign _0938_ = _0904_ ? _0933_ : 2'h0;
  assign _0939_ = _0904_ ? _0934_ : 1'h0;
  assign _0940_ = _0904_ ? _0935_ : 1'h0;
  assign _0941_ = r2[309:308] == 2'h0;
  assign _0942_ = r2[309:308] == 2'h1;
  assign _0943_ = r2[309:308] == 2'h2;
  function [63:0] \22137 ;
    input [63:0] a;
    input [191:0] b;
    input [2:0] s;
    (* parallel_case *)
    casez (s)
      3'b??1:
        \22137  = b[63:0];
      3'b?1?:
        \22137  = b[127:64];
      3'b1??:
        \22137  = b[191:128];
      default:
        \22137  = a;
    endcase
  endfunction
  assign _0944_ = \22137 ({ _0490_, _0479_, _0468_, _0457_, _0446_, _0435_, _0424_, _0413_ }, { load_dp_data, r2[373:310], _0826_ }, { _0943_, _0942_, _0941_ });
  assign _0945_ = stage1_issue_enable ? stage1_dcreq : _0898_;
  assign _0946_ = stage1_issue_enable ? { stage1_req[77:14], stage1_req[193:192], stage1_req[189:187], stage1_req[191], stage1_req[5], stage1_req[2] } : { r2[77:14], r2[193:192], r2[189:187], r2[191], r2[5], r2[2] };
  assign _0947_ = stage1_issue_enable ? stage1_req[85:78] : r2[85:78];
  assign _0948_ = stage1_dreq ? store_data : r2[157:94];
  assign _0949_ = r2[0] & r2[194];
  assign _0950_ = _0949_ & \d_in.valid ;
  assign _0951_ = _0901_ | _0902_;
  assign _0952_ = r2[190] & complete;
  assign _0953_ = complete | _0903_;
  assign _0954_ = _0953_ | _0904_;
  assign _0955_ = ~ _0954_;
  assign _0956_ = r2[0] & _0955_;
  assign _0959_ = _0290_[2] ? _0958_ : _0957_;
  assign _0962_ = _0292_[2] ? _0961_ : _0960_;
  assign _0965_ = _0294_[2] ? _0964_ : _0963_;
  assign _0968_ = _0296_[2] ? _0967_ : _0966_;
  assign _0971_ = _0298_[2] ? _0970_ : _0969_;
  assign _0974_ = _0300_[2] ? _0973_ : _0972_;
  assign _0977_ = _0302_[2] ? _0976_ : _0975_;
  assign _0980_ = _0304_[2] ? _0979_ : _0978_;
  assign _0983_ = r2[296] ? _0982_ : _0981_;
  assign _0986_ = r2[293] ? _0985_ : _0984_;
  assign _0989_ = r2[290] ? _0988_ : _0987_;
  assign _0992_ = r2[287] ? _0991_ : _0990_;
  assign _0995_ = r2[284] ? _0994_ : _0993_;
  assign _0998_ = r2[281] ? _0997_ : _0996_;
  assign _1001_ = r2[278] ? _1000_ : _0999_;
  assign _1004_ = r2[275] ? _1003_ : _1002_;
  assign req_in = { \l_in.nia , _0150_, 1'h0, _0199_, _0198_, \l_in.insn [15:11], \l_in.insn [20:16], _0197_, \l_in.priv_mode , \l_in.virt_mode , _0141_, \l_in.rc , _0170_, _0166_, \l_in.reserve , \l_in.xerc , \l_in.update , \l_in.sign_extend , _0206_, \l_in.byte_reverse , \l_in.length , \l_in.length , \l_in.write_reg , \l_in.instr_tag , _0130_, _0148_, _0196_, \l_in.mode_32bit , 1'h0, _0195_, 1'h0, _0194_, _0193_, _0192_, _0191_, _0190_, _0189_, _0188_, _0187_, _0204_, \l_in.valid  };
  assign r1 = _0085_;
  assign r1in = { _0271_, _0288_, _0276_, _0275_, _0277_, _0273_, _0281_, _0280_ };
  assign r2 = _0086_;
  assign r2in = { _0352_, _0351_, _0350_, _0354_ };
  assign r3 = _0087_;
  assign r3in = { _0897_, _0915_, _0913_, 1'h0, _0940_, 1'h0, _0939_, 8'h00, _0938_, 2'h0, _0937_, _0904_, _0912_, _0683_, _0680_, _0674_, _0662_, _0779_, _0747_, _0491_, _0446_, _0435_, _0424_, _0413_, _0936_, _0811_, _0894_, r3[83:2], _0911_ };
  assign busy = _0216_;
  assign complete = _0221_;
  assign in_progress = _0224_;
  assign flushing = _0088_;
  assign store_sp_data = { \l_in.data [63], _0105_, _0104_ };
  assign load_dp_data = { r3[276], _0116_, _0127_, 29'h00000000 };
  assign store_data = { _0980_, _0977_, _0974_, _0971_, _0968_, _0965_, _0962_, _0959_ };
  assign stage1_issue_enable = _0230_;
  assign stage1_req = { _0276_, _0275_, _0277_, _0273_, _0281_, _0280_ };
  assign stage1_dcreq = _0287_;
  assign stage1_dreq = _0089_;
  assign stage2_busy_next = _0353_;
  assign stage3_busy_next = _0956_;
  assign \e_out.busy  = busy;
  assign \e_out.in_progress  = in_progress;
  assign \e_out.interrupt  = r3[285];
  assign \l_out.valid  = complete;
  assign \l_out.instr_tag  = r2[160:158];
  assign \l_out.write_enable  = _0951_;
  assign \l_out.write_reg  = r2[167:161];
  assign \l_out.write_data  = _0944_;
  assign \l_out.xerc  = r2[186:182];
  assign \l_out.rc  = _0952_;
  assign \l_out.store_done  = \d_in.store_done ;
  assign \l_out.interrupt  = r3[285];
  assign \l_out.intr_vec  = r3[297:286];
  assign \l_out.srr0  = r3[361:298];
  assign \l_out.srr1  = r3[377:362];
  assign \d_out.valid  = _0945_;
  assign \d_out.hold  = _0950_;
  assign \d_out.load  = _0946_[0];
  assign \d_out.dcbz  = _0946_[1];
  assign \d_out.nc  = _0946_[2];
  assign \d_out.reserve  = _0946_[3];
  assign \d_out.atomic  = _0946_[4];
  assign \d_out.atomic_last  = _0946_[5];
  assign \d_out.virt_mode  = _0946_[6];
  assign \d_out.priv_mode  = _0946_[7];
  assign \d_out.addr  = _0946_[71:8];
  assign \d_out.data  = _0948_;
  assign \d_out.byte_sel  = _0947_;
  assign \m_out.valid  = _0899_;
  assign \m_out.tlbie  = r2[4];
  assign \m_out.slbia  = r2[205];
  assign \m_out.mtspr  = _0900_;
  assign \m_out.iside  = r2[9];
  assign \m_out.load  = r2[2];
  assign \m_out.priv  = r2[193];
  assign \m_out.sprn  = r2[204:195];
  assign \m_out.addr  = r2[77:14];
  assign \m_out.rs  = r2[157:94];
  assign \events.load_complete  = r3[378];
  assign \events.store_complete  = r3[379];
  assign \events.itlb_miss  = r3[380];
  assign log_out = 10'hzzz;
endmodule