module lsu_bypass
(
  clk_i,
  rst_ni,
  flush_i,
  lsu_req_i,
  lus_req_valid_i,
  pop_ld_i,
  pop_st_i,
  lsu_ctrl_o,
  ready_o
);

  input [150:0] lsu_req_i;
  output [150:0] lsu_ctrl_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input lus_req_valid_i;
  input pop_ld_i;
  input pop_st_i;
  output ready_o;
  wire [150:0] lsu_ctrl_o;
  wire ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,read_pointer_n,write_pointer_n,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413;
  wire [301:0] mem_n;
  wire [1:0] status_cnt_n;
  reg N41,N17;
  reg [301:0] mem_q;
  reg [1:0] status_cnt_q;
  assign N206 = (N43)? mem_q[150] : 
                (N0)? mem_q[301] : 1'b0;
  assign N0 = N41;
  assign N207 = (N43)? mem_q[149] : 
                (N0)? mem_q[300] : 1'b0;
  assign N208 = (N43)? mem_q[148] : 
                (N0)? mem_q[299] : 1'b0;
  assign N209 = (N43)? mem_q[147] : 
                (N0)? mem_q[298] : 1'b0;
  assign N210 = (N43)? mem_q[146] : 
                (N0)? mem_q[297] : 1'b0;
  assign N211 = (N43)? mem_q[145] : 
                (N0)? mem_q[296] : 1'b0;
  assign N212 = (N43)? mem_q[144] : 
                (N0)? mem_q[295] : 1'b0;
  assign N213 = (N43)? mem_q[143] : 
                (N0)? mem_q[294] : 1'b0;
  assign N214 = (N43)? mem_q[142] : 
                (N0)? mem_q[293] : 1'b0;
  assign N215 = (N43)? mem_q[141] : 
                (N0)? mem_q[292] : 1'b0;
  assign N216 = (N43)? mem_q[140] : 
                (N0)? mem_q[291] : 1'b0;
  assign N217 = (N43)? mem_q[139] : 
                (N0)? mem_q[290] : 1'b0;
  assign N218 = (N43)? mem_q[138] : 
                (N0)? mem_q[289] : 1'b0;
  assign N219 = (N43)? mem_q[137] : 
                (N0)? mem_q[288] : 1'b0;
  assign N220 = (N43)? mem_q[136] : 
                (N0)? mem_q[287] : 1'b0;
  assign N221 = (N43)? mem_q[135] : 
                (N0)? mem_q[286] : 1'b0;
  assign N222 = (N43)? mem_q[134] : 
                (N0)? mem_q[285] : 1'b0;
  assign N223 = (N43)? mem_q[133] : 
                (N0)? mem_q[284] : 1'b0;
  assign N224 = (N43)? mem_q[132] : 
                (N0)? mem_q[283] : 1'b0;
  assign N225 = (N43)? mem_q[131] : 
                (N0)? mem_q[282] : 1'b0;
  assign N226 = (N43)? mem_q[130] : 
                (N0)? mem_q[281] : 1'b0;
  assign N227 = (N43)? mem_q[129] : 
                (N0)? mem_q[280] : 1'b0;
  assign N228 = (N43)? mem_q[128] : 
                (N0)? mem_q[279] : 1'b0;
  assign N229 = (N43)? mem_q[127] : 
                (N0)? mem_q[278] : 1'b0;
  assign N230 = (N43)? mem_q[126] : 
                (N0)? mem_q[277] : 1'b0;
  assign N231 = (N43)? mem_q[125] : 
                (N0)? mem_q[276] : 1'b0;
  assign N232 = (N43)? mem_q[124] : 
                (N0)? mem_q[275] : 1'b0;
  assign N233 = (N43)? mem_q[123] : 
                (N0)? mem_q[274] : 1'b0;
  assign N234 = (N43)? mem_q[122] : 
                (N0)? mem_q[273] : 1'b0;
  assign N235 = (N43)? mem_q[121] : 
                (N0)? mem_q[272] : 1'b0;
  assign N236 = (N43)? mem_q[120] : 
                (N0)? mem_q[271] : 1'b0;
  assign N237 = (N43)? mem_q[119] : 
                (N0)? mem_q[270] : 1'b0;
  assign N238 = (N43)? mem_q[118] : 
                (N0)? mem_q[269] : 1'b0;
  assign N239 = (N43)? mem_q[117] : 
                (N0)? mem_q[268] : 1'b0;
  assign N240 = (N43)? mem_q[116] : 
                (N0)? mem_q[267] : 1'b0;
  assign N241 = (N43)? mem_q[115] : 
                (N0)? mem_q[266] : 1'b0;
  assign N242 = (N43)? mem_q[114] : 
                (N0)? mem_q[265] : 1'b0;
  assign N243 = (N43)? mem_q[113] : 
                (N0)? mem_q[264] : 1'b0;
  assign N244 = (N43)? mem_q[112] : 
                (N0)? mem_q[263] : 1'b0;
  assign N245 = (N43)? mem_q[111] : 
                (N0)? mem_q[262] : 1'b0;
  assign N246 = (N43)? mem_q[110] : 
                (N0)? mem_q[261] : 1'b0;
  assign N247 = (N43)? mem_q[109] : 
                (N0)? mem_q[260] : 1'b0;
  assign N248 = (N43)? mem_q[108] : 
                (N0)? mem_q[259] : 1'b0;
  assign N249 = (N43)? mem_q[107] : 
                (N0)? mem_q[258] : 1'b0;
  assign N250 = (N43)? mem_q[106] : 
                (N0)? mem_q[257] : 1'b0;
  assign N251 = (N43)? mem_q[105] : 
                (N0)? mem_q[256] : 1'b0;
  assign N252 = (N43)? mem_q[104] : 
                (N0)? mem_q[255] : 1'b0;
  assign N253 = (N43)? mem_q[103] : 
                (N0)? mem_q[254] : 1'b0;
  assign N254 = (N43)? mem_q[102] : 
                (N0)? mem_q[253] : 1'b0;
  assign N255 = (N43)? mem_q[101] : 
                (N0)? mem_q[252] : 1'b0;
  assign N256 = (N43)? mem_q[100] : 
                (N0)? mem_q[251] : 1'b0;
  assign N257 = (N43)? mem_q[99] : 
                (N0)? mem_q[250] : 1'b0;
  assign N258 = (N43)? mem_q[98] : 
                (N0)? mem_q[249] : 1'b0;
  assign N259 = (N43)? mem_q[97] : 
                (N0)? mem_q[248] : 1'b0;
  assign N260 = (N43)? mem_q[96] : 
                (N0)? mem_q[247] : 1'b0;
  assign N261 = (N43)? mem_q[95] : 
                (N0)? mem_q[246] : 1'b0;
  assign N262 = (N43)? mem_q[94] : 
                (N0)? mem_q[245] : 1'b0;
  assign N263 = (N43)? mem_q[93] : 
                (N0)? mem_q[244] : 1'b0;
  assign N264 = (N43)? mem_q[92] : 
                (N0)? mem_q[243] : 1'b0;
  assign N265 = (N43)? mem_q[91] : 
                (N0)? mem_q[242] : 1'b0;
  assign N266 = (N43)? mem_q[90] : 
                (N0)? mem_q[241] : 1'b0;
  assign N267 = (N43)? mem_q[89] : 
                (N0)? mem_q[240] : 1'b0;
  assign N268 = (N43)? mem_q[88] : 
                (N0)? mem_q[239] : 1'b0;
  assign N269 = (N43)? mem_q[87] : 
                (N0)? mem_q[238] : 1'b0;
  assign N270 = (N43)? mem_q[86] : 
                (N0)? mem_q[237] : 1'b0;
  assign N271 = (N43)? mem_q[85] : 
                (N0)? mem_q[236] : 1'b0;
  assign N272 = (N43)? mem_q[84] : 
                (N0)? mem_q[235] : 1'b0;
  assign N273 = (N43)? mem_q[83] : 
                (N0)? mem_q[234] : 1'b0;
  assign N274 = (N43)? mem_q[82] : 
                (N0)? mem_q[233] : 1'b0;
  assign N275 = (N43)? mem_q[81] : 
                (N0)? mem_q[232] : 1'b0;
  assign N276 = (N43)? mem_q[80] : 
                (N0)? mem_q[231] : 1'b0;
  assign N277 = (N43)? mem_q[79] : 
                (N0)? mem_q[230] : 1'b0;
  assign N278 = (N43)? mem_q[78] : 
                (N0)? mem_q[229] : 1'b0;
  assign N279 = (N43)? mem_q[77] : 
                (N0)? mem_q[228] : 1'b0;
  assign N280 = (N43)? mem_q[76] : 
                (N0)? mem_q[227] : 1'b0;
  assign N281 = (N43)? mem_q[75] : 
                (N0)? mem_q[226] : 1'b0;
  assign N282 = (N43)? mem_q[74] : 
                (N0)? mem_q[225] : 1'b0;
  assign N283 = (N43)? mem_q[73] : 
                (N0)? mem_q[224] : 1'b0;
  assign N284 = (N43)? mem_q[72] : 
                (N0)? mem_q[223] : 1'b0;
  assign N285 = (N43)? mem_q[71] : 
                (N0)? mem_q[222] : 1'b0;
  assign N286 = (N43)? mem_q[70] : 
                (N0)? mem_q[221] : 1'b0;
  assign N287 = (N43)? mem_q[69] : 
                (N0)? mem_q[220] : 1'b0;
  assign N288 = (N43)? mem_q[68] : 
                (N0)? mem_q[219] : 1'b0;
  assign N289 = (N43)? mem_q[67] : 
                (N0)? mem_q[218] : 1'b0;
  assign N290 = (N43)? mem_q[66] : 
                (N0)? mem_q[217] : 1'b0;
  assign N291 = (N43)? mem_q[65] : 
                (N0)? mem_q[216] : 1'b0;
  assign N292 = (N43)? mem_q[64] : 
                (N0)? mem_q[215] : 1'b0;
  assign N293 = (N43)? mem_q[63] : 
                (N0)? mem_q[214] : 1'b0;
  assign N294 = (N43)? mem_q[62] : 
                (N0)? mem_q[213] : 1'b0;
  assign N295 = (N43)? mem_q[61] : 
                (N0)? mem_q[212] : 1'b0;
  assign N296 = (N43)? mem_q[60] : 
                (N0)? mem_q[211] : 1'b0;
  assign N297 = (N43)? mem_q[59] : 
                (N0)? mem_q[210] : 1'b0;
  assign N298 = (N43)? mem_q[58] : 
                (N0)? mem_q[209] : 1'b0;
  assign N299 = (N43)? mem_q[57] : 
                (N0)? mem_q[208] : 1'b0;
  assign N300 = (N43)? mem_q[56] : 
                (N0)? mem_q[207] : 1'b0;
  assign N301 = (N43)? mem_q[55] : 
                (N0)? mem_q[206] : 1'b0;
  assign N302 = (N43)? mem_q[54] : 
                (N0)? mem_q[205] : 1'b0;
  assign N303 = (N43)? mem_q[53] : 
                (N0)? mem_q[204] : 1'b0;
  assign N304 = (N43)? mem_q[52] : 
                (N0)? mem_q[203] : 1'b0;
  assign N305 = (N43)? mem_q[51] : 
                (N0)? mem_q[202] : 1'b0;
  assign N306 = (N43)? mem_q[50] : 
                (N0)? mem_q[201] : 1'b0;
  assign N307 = (N43)? mem_q[49] : 
                (N0)? mem_q[200] : 1'b0;
  assign N308 = (N43)? mem_q[48] : 
                (N0)? mem_q[199] : 1'b0;
  assign N309 = (N43)? mem_q[47] : 
                (N0)? mem_q[198] : 1'b0;
  assign N310 = (N43)? mem_q[46] : 
                (N0)? mem_q[197] : 1'b0;
  assign N311 = (N43)? mem_q[45] : 
                (N0)? mem_q[196] : 1'b0;
  assign N312 = (N43)? mem_q[44] : 
                (N0)? mem_q[195] : 1'b0;
  assign N313 = (N43)? mem_q[43] : 
                (N0)? mem_q[194] : 1'b0;
  assign N314 = (N43)? mem_q[42] : 
                (N0)? mem_q[193] : 1'b0;
  assign N315 = (N43)? mem_q[41] : 
                (N0)? mem_q[192] : 1'b0;
  assign N316 = (N43)? mem_q[40] : 
                (N0)? mem_q[191] : 1'b0;
  assign N317 = (N43)? mem_q[39] : 
                (N0)? mem_q[190] : 1'b0;
  assign N318 = (N43)? mem_q[38] : 
                (N0)? mem_q[189] : 1'b0;
  assign N319 = (N43)? mem_q[37] : 
                (N0)? mem_q[188] : 1'b0;
  assign N320 = (N43)? mem_q[36] : 
                (N0)? mem_q[187] : 1'b0;
  assign N321 = (N43)? mem_q[35] : 
                (N0)? mem_q[186] : 1'b0;
  assign N322 = (N43)? mem_q[34] : 
                (N0)? mem_q[185] : 1'b0;
  assign N323 = (N43)? mem_q[33] : 
                (N0)? mem_q[184] : 1'b0;
  assign N324 = (N43)? mem_q[32] : 
                (N0)? mem_q[183] : 1'b0;
  assign N325 = (N43)? mem_q[31] : 
                (N0)? mem_q[182] : 1'b0;
  assign N326 = (N43)? mem_q[30] : 
                (N0)? mem_q[181] : 1'b0;
  assign N327 = (N43)? mem_q[29] : 
                (N0)? mem_q[180] : 1'b0;
  assign N328 = (N43)? mem_q[28] : 
                (N0)? mem_q[179] : 1'b0;
  assign N329 = (N43)? mem_q[27] : 
                (N0)? mem_q[178] : 1'b0;
  assign N330 = (N43)? mem_q[26] : 
                (N0)? mem_q[177] : 1'b0;
  assign N331 = (N43)? mem_q[25] : 
                (N0)? mem_q[176] : 1'b0;
  assign N332 = (N43)? mem_q[24] : 
                (N0)? mem_q[175] : 1'b0;
  assign N333 = (N43)? mem_q[23] : 
                (N0)? mem_q[174] : 1'b0;
  assign N334 = (N43)? mem_q[22] : 
                (N0)? mem_q[173] : 1'b0;
  assign N335 = (N43)? mem_q[21] : 
                (N0)? mem_q[172] : 1'b0;
  assign N336 = (N43)? mem_q[20] : 
                (N0)? mem_q[171] : 1'b0;
  assign N337 = (N43)? mem_q[19] : 
                (N0)? mem_q[170] : 1'b0;
  assign N338 = (N43)? mem_q[18] : 
                (N0)? mem_q[169] : 1'b0;
  assign N339 = (N43)? mem_q[17] : 
                (N0)? mem_q[168] : 1'b0;
  assign N340 = (N43)? mem_q[16] : 
                (N0)? mem_q[167] : 1'b0;
  assign N341 = (N43)? mem_q[15] : 
                (N0)? mem_q[166] : 1'b0;
  assign N342 = (N43)? mem_q[14] : 
                (N0)? mem_q[165] : 1'b0;
  assign N343 = (N43)? mem_q[13] : 
                (N0)? mem_q[164] : 1'b0;
  assign N344 = (N43)? mem_q[12] : 
                (N0)? mem_q[163] : 1'b0;
  assign N345 = (N43)? mem_q[11] : 
                (N0)? mem_q[162] : 1'b0;
  assign N346 = (N43)? mem_q[10] : 
                (N0)? mem_q[161] : 1'b0;
  assign N347 = (N43)? mem_q[9] : 
                (N0)? mem_q[160] : 1'b0;
  assign N348 = (N43)? mem_q[8] : 
                (N0)? mem_q[159] : 1'b0;
  assign N349 = (N43)? mem_q[7] : 
                (N0)? mem_q[158] : 1'b0;
  assign N350 = (N43)? mem_q[6] : 
                (N0)? mem_q[157] : 1'b0;
  assign N351 = (N43)? mem_q[5] : 
                (N0)? mem_q[156] : 1'b0;
  assign N352 = (N43)? mem_q[4] : 
                (N0)? mem_q[155] : 1'b0;
  assign N353 = (N43)? mem_q[3] : 
                (N0)? mem_q[154] : 1'b0;
  assign N354 = (N43)? mem_q[2] : 
                (N0)? mem_q[153] : 1'b0;
  assign N355 = (N43)? mem_q[1] : 
                (N0)? mem_q[152] : 1'b0;
  assign N356 = (N43)? mem_q[0] : 
                (N0)? mem_q[151] : 1'b0;

  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      N41 <= 1'b0;
    end else if(1'b1) begin
      N41 <= read_pointer_n;
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[301] <= 1'b0;
    end else if(1'b1) begin
      mem_q[301] <= mem_n[301];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[300] <= 1'b0;
    end else if(N364) begin
      mem_q[300] <= mem_n[300];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[299] <= 1'b0;
    end else if(N371) begin
      mem_q[299] <= mem_n[299];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[298] <= 1'b0;
    end else if(N378) begin
      mem_q[298] <= mem_n[298];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[297] <= 1'b0;
    end else if(N382) begin
      mem_q[297] <= mem_n[297];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[296] <= 1'b0;
    end else if(N382) begin
      mem_q[296] <= mem_n[296];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[295] <= 1'b0;
    end else if(N382) begin
      mem_q[295] <= mem_n[295];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[294] <= 1'b0;
    end else if(N382) begin
      mem_q[294] <= mem_n[294];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[293] <= 1'b0;
    end else if(N382) begin
      mem_q[293] <= mem_n[293];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[292] <= 1'b0;
    end else if(N382) begin
      mem_q[292] <= mem_n[292];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[291] <= 1'b0;
    end else if(N382) begin
      mem_q[291] <= mem_n[291];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[290] <= 1'b0;
    end else if(N382) begin
      mem_q[290] <= mem_n[290];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[289] <= 1'b0;
    end else if(N382) begin
      mem_q[289] <= mem_n[289];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[288] <= 1'b0;
    end else if(N382) begin
      mem_q[288] <= mem_n[288];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[287] <= 1'b0;
    end else if(N382) begin
      mem_q[287] <= mem_n[287];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[286] <= 1'b0;
    end else if(N382) begin
      mem_q[286] <= mem_n[286];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[285] <= 1'b0;
    end else if(N382) begin
      mem_q[285] <= mem_n[285];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[284] <= 1'b0;
    end else if(N382) begin
      mem_q[284] <= mem_n[284];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[283] <= 1'b0;
    end else if(N382) begin
      mem_q[283] <= mem_n[283];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[282] <= 1'b0;
    end else if(N382) begin
      mem_q[282] <= mem_n[282];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[281] <= 1'b0;
    end else if(N382) begin
      mem_q[281] <= mem_n[281];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[280] <= 1'b0;
    end else if(N382) begin
      mem_q[280] <= mem_n[280];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[279] <= 1'b0;
    end else if(N382) begin
      mem_q[279] <= mem_n[279];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[278] <= 1'b0;
    end else if(N382) begin
      mem_q[278] <= mem_n[278];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[277] <= 1'b0;
    end else if(N382) begin
      mem_q[277] <= mem_n[277];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[276] <= 1'b0;
    end else if(N382) begin
      mem_q[276] <= mem_n[276];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[275] <= 1'b0;
    end else if(N382) begin
      mem_q[275] <= mem_n[275];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[274] <= 1'b0;
    end else if(N382) begin
      mem_q[274] <= mem_n[274];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[273] <= 1'b0;
    end else if(N382) begin
      mem_q[273] <= mem_n[273];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[272] <= 1'b0;
    end else if(N382) begin
      mem_q[272] <= mem_n[272];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[271] <= 1'b0;
    end else if(N382) begin
      mem_q[271] <= mem_n[271];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[270] <= 1'b0;
    end else if(N382) begin
      mem_q[270] <= mem_n[270];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[269] <= 1'b0;
    end else if(N382) begin
      mem_q[269] <= mem_n[269];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[268] <= 1'b0;
    end else if(N382) begin
      mem_q[268] <= mem_n[268];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[267] <= 1'b0;
    end else if(N382) begin
      mem_q[267] <= mem_n[267];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[266] <= 1'b0;
    end else if(N382) begin
      mem_q[266] <= mem_n[266];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[265] <= 1'b0;
    end else if(N382) begin
      mem_q[265] <= mem_n[265];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[264] <= 1'b0;
    end else if(N382) begin
      mem_q[264] <= mem_n[264];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[263] <= 1'b0;
    end else if(N382) begin
      mem_q[263] <= mem_n[263];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[262] <= 1'b0;
    end else if(N382) begin
      mem_q[262] <= mem_n[262];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[261] <= 1'b0;
    end else if(N382) begin
      mem_q[261] <= mem_n[261];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[260] <= 1'b0;
    end else if(N382) begin
      mem_q[260] <= mem_n[260];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[259] <= 1'b0;
    end else if(N382) begin
      mem_q[259] <= mem_n[259];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[258] <= 1'b0;
    end else if(N382) begin
      mem_q[258] <= mem_n[258];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[257] <= 1'b0;
    end else if(N382) begin
      mem_q[257] <= mem_n[257];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[256] <= 1'b0;
    end else if(N382) begin
      mem_q[256] <= mem_n[256];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[255] <= 1'b0;
    end else if(N382) begin
      mem_q[255] <= mem_n[255];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[254] <= 1'b0;
    end else if(N382) begin
      mem_q[254] <= mem_n[254];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[253] <= 1'b0;
    end else if(N382) begin
      mem_q[253] <= mem_n[253];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[252] <= 1'b0;
    end else if(N382) begin
      mem_q[252] <= mem_n[252];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[251] <= 1'b0;
    end else if(N382) begin
      mem_q[251] <= mem_n[251];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[250] <= 1'b0;
    end else if(N382) begin
      mem_q[250] <= mem_n[250];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[249] <= 1'b0;
    end else if(N382) begin
      mem_q[249] <= mem_n[249];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[248] <= 1'b0;
    end else if(N385) begin
      mem_q[248] <= mem_n[248];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[247] <= 1'b0;
    end else if(N387) begin
      mem_q[247] <= mem_n[247];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[246] <= 1'b0;
    end else if(N387) begin
      mem_q[246] <= mem_n[246];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[245] <= 1'b0;
    end else if(N387) begin
      mem_q[245] <= mem_n[245];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[244] <= 1'b0;
    end else if(N387) begin
      mem_q[244] <= mem_n[244];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[243] <= 1'b0;
    end else if(N387) begin
      mem_q[243] <= mem_n[243];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[242] <= 1'b0;
    end else if(N387) begin
      mem_q[242] <= mem_n[242];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[241] <= 1'b0;
    end else if(N387) begin
      mem_q[241] <= mem_n[241];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[240] <= 1'b0;
    end else if(N387) begin
      mem_q[240] <= mem_n[240];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[239] <= 1'b0;
    end else if(N387) begin
      mem_q[239] <= mem_n[239];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[238] <= 1'b0;
    end else if(N387) begin
      mem_q[238] <= mem_n[238];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[237] <= 1'b0;
    end else if(N387) begin
      mem_q[237] <= mem_n[237];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[236] <= 1'b0;
    end else if(N387) begin
      mem_q[236] <= mem_n[236];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[235] <= 1'b0;
    end else if(N387) begin
      mem_q[235] <= mem_n[235];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[234] <= 1'b0;
    end else if(N387) begin
      mem_q[234] <= mem_n[234];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[233] <= 1'b0;
    end else if(N387) begin
      mem_q[233] <= mem_n[233];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[232] <= 1'b0;
    end else if(N387) begin
      mem_q[232] <= mem_n[232];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[231] <= 1'b0;
    end else if(N387) begin
      mem_q[231] <= mem_n[231];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[230] <= 1'b0;
    end else if(N387) begin
      mem_q[230] <= mem_n[230];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[229] <= 1'b0;
    end else if(N387) begin
      mem_q[229] <= mem_n[229];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[228] <= 1'b0;
    end else if(N387) begin
      mem_q[228] <= mem_n[228];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[227] <= 1'b0;
    end else if(N387) begin
      mem_q[227] <= mem_n[227];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[226] <= 1'b0;
    end else if(N387) begin
      mem_q[226] <= mem_n[226];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[225] <= 1'b0;
    end else if(N387) begin
      mem_q[225] <= mem_n[225];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[224] <= 1'b0;
    end else if(N387) begin
      mem_q[224] <= mem_n[224];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[223] <= 1'b0;
    end else if(N387) begin
      mem_q[223] <= mem_n[223];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[222] <= 1'b0;
    end else if(N387) begin
      mem_q[222] <= mem_n[222];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[221] <= 1'b0;
    end else if(N387) begin
      mem_q[221] <= mem_n[221];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[220] <= 1'b0;
    end else if(N387) begin
      mem_q[220] <= mem_n[220];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[219] <= 1'b0;
    end else if(N387) begin
      mem_q[219] <= mem_n[219];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[218] <= 1'b0;
    end else if(N387) begin
      mem_q[218] <= mem_n[218];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[217] <= 1'b0;
    end else if(N387) begin
      mem_q[217] <= mem_n[217];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[216] <= 1'b0;
    end else if(N387) begin
      mem_q[216] <= mem_n[216];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[215] <= 1'b0;
    end else if(N387) begin
      mem_q[215] <= mem_n[215];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[214] <= 1'b0;
    end else if(N387) begin
      mem_q[214] <= mem_n[214];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[213] <= 1'b0;
    end else if(N387) begin
      mem_q[213] <= mem_n[213];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[212] <= 1'b0;
    end else if(N387) begin
      mem_q[212] <= mem_n[212];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[211] <= 1'b0;
    end else if(N387) begin
      mem_q[211] <= mem_n[211];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[210] <= 1'b0;
    end else if(N387) begin
      mem_q[210] <= mem_n[210];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[209] <= 1'b0;
    end else if(N387) begin
      mem_q[209] <= mem_n[209];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[208] <= 1'b0;
    end else if(N387) begin
      mem_q[208] <= mem_n[208];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[207] <= 1'b0;
    end else if(N387) begin
      mem_q[207] <= mem_n[207];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[206] <= 1'b0;
    end else if(N387) begin
      mem_q[206] <= mem_n[206];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[205] <= 1'b0;
    end else if(N387) begin
      mem_q[205] <= mem_n[205];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[204] <= 1'b0;
    end else if(N387) begin
      mem_q[204] <= mem_n[204];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[203] <= 1'b0;
    end else if(N387) begin
      mem_q[203] <= mem_n[203];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[202] <= 1'b0;
    end else if(N387) begin
      mem_q[202] <= mem_n[202];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[201] <= 1'b0;
    end else if(N387) begin
      mem_q[201] <= mem_n[201];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[200] <= 1'b0;
    end else if(N387) begin
      mem_q[200] <= mem_n[200];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[199] <= 1'b0;
    end else if(N387) begin
      mem_q[199] <= mem_n[199];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[198] <= 1'b0;
    end else if(N391) begin
      mem_q[198] <= mem_n[198];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[197] <= 1'b0;
    end else if(N391) begin
      mem_q[197] <= mem_n[197];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[196] <= 1'b0;
    end else if(N391) begin
      mem_q[196] <= mem_n[196];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[195] <= 1'b0;
    end else if(N391) begin
      mem_q[195] <= mem_n[195];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[194] <= 1'b0;
    end else if(N391) begin
      mem_q[194] <= mem_n[194];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[193] <= 1'b0;
    end else if(N391) begin
      mem_q[193] <= mem_n[193];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[192] <= 1'b0;
    end else if(N391) begin
      mem_q[192] <= mem_n[192];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[191] <= 1'b0;
    end else if(N391) begin
      mem_q[191] <= mem_n[191];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[190] <= 1'b0;
    end else if(N391) begin
      mem_q[190] <= mem_n[190];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[189] <= 1'b0;
    end else if(N391) begin
      mem_q[189] <= mem_n[189];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[188] <= 1'b0;
    end else if(N391) begin
      mem_q[188] <= mem_n[188];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[187] <= 1'b0;
    end else if(N391) begin
      mem_q[187] <= mem_n[187];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[186] <= 1'b0;
    end else if(N391) begin
      mem_q[186] <= mem_n[186];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[185] <= 1'b0;
    end else if(N391) begin
      mem_q[185] <= mem_n[185];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[184] <= 1'b0;
    end else if(N391) begin
      mem_q[184] <= mem_n[184];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[183] <= 1'b0;
    end else if(N391) begin
      mem_q[183] <= mem_n[183];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[182] <= 1'b0;
    end else if(N391) begin
      mem_q[182] <= mem_n[182];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[181] <= 1'b0;
    end else if(N391) begin
      mem_q[181] <= mem_n[181];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[180] <= 1'b0;
    end else if(N391) begin
      mem_q[180] <= mem_n[180];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[179] <= 1'b0;
    end else if(N391) begin
      mem_q[179] <= mem_n[179];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[178] <= 1'b0;
    end else if(N391) begin
      mem_q[178] <= mem_n[178];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[177] <= 1'b0;
    end else if(N391) begin
      mem_q[177] <= mem_n[177];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[176] <= 1'b0;
    end else if(N391) begin
      mem_q[176] <= mem_n[176];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[175] <= 1'b0;
    end else if(N391) begin
      mem_q[175] <= mem_n[175];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[174] <= 1'b0;
    end else if(N391) begin
      mem_q[174] <= mem_n[174];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[173] <= 1'b0;
    end else if(N391) begin
      mem_q[173] <= mem_n[173];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[172] <= 1'b0;
    end else if(N391) begin
      mem_q[172] <= mem_n[172];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[171] <= 1'b0;
    end else if(N391) begin
      mem_q[171] <= mem_n[171];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[170] <= 1'b0;
    end else if(N391) begin
      mem_q[170] <= mem_n[170];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[169] <= 1'b0;
    end else if(N391) begin
      mem_q[169] <= mem_n[169];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[168] <= 1'b0;
    end else if(N391) begin
      mem_q[168] <= mem_n[168];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[167] <= 1'b0;
    end else if(N391) begin
      mem_q[167] <= mem_n[167];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[166] <= 1'b0;
    end else if(N391) begin
      mem_q[166] <= mem_n[166];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[165] <= 1'b0;
    end else if(N391) begin
      mem_q[165] <= mem_n[165];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[164] <= 1'b0;
    end else if(N391) begin
      mem_q[164] <= mem_n[164];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[163] <= 1'b0;
    end else if(N391) begin
      mem_q[163] <= mem_n[163];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[162] <= 1'b0;
    end else if(N391) begin
      mem_q[162] <= mem_n[162];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[161] <= 1'b0;
    end else if(N391) begin
      mem_q[161] <= mem_n[161];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[160] <= 1'b0;
    end else if(N391) begin
      mem_q[160] <= mem_n[160];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[159] <= 1'b0;
    end else if(N391) begin
      mem_q[159] <= mem_n[159];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[158] <= 1'b0;
    end else if(N391) begin
      mem_q[158] <= mem_n[158];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[157] <= 1'b0;
    end else if(N391) begin
      mem_q[157] <= mem_n[157];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[156] <= 1'b0;
    end else if(N391) begin
      mem_q[156] <= mem_n[156];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[155] <= 1'b0;
    end else if(N391) begin
      mem_q[155] <= mem_n[155];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[154] <= 1'b0;
    end else if(N391) begin
      mem_q[154] <= mem_n[154];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[153] <= 1'b0;
    end else if(N391) begin
      mem_q[153] <= mem_n[153];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[152] <= 1'b0;
    end else if(N391) begin
      mem_q[152] <= mem_n[152];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[151] <= 1'b0;
    end else if(N391) begin
      mem_q[151] <= mem_n[151];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[150] <= 1'b0;
    end else if(1'b1) begin
      mem_q[150] <= mem_n[150];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[149] <= 1'b0;
    end else if(N394) begin
      mem_q[149] <= mem_n[149];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[148] <= 1'b0;
    end else if(N397) begin
      mem_q[148] <= mem_n[148];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[147] <= 1'b0;
    end else if(N400) begin
      mem_q[147] <= mem_n[147];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[146] <= 1'b0;
    end else if(N400) begin
      mem_q[146] <= mem_n[146];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[145] <= 1'b0;
    end else if(N400) begin
      mem_q[145] <= mem_n[145];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[144] <= 1'b0;
    end else if(N400) begin
      mem_q[144] <= mem_n[144];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[143] <= 1'b0;
    end else if(N400) begin
      mem_q[143] <= mem_n[143];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[142] <= 1'b0;
    end else if(N400) begin
      mem_q[142] <= mem_n[142];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[141] <= 1'b0;
    end else if(N400) begin
      mem_q[141] <= mem_n[141];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[140] <= 1'b0;
    end else if(N400) begin
      mem_q[140] <= mem_n[140];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[139] <= 1'b0;
    end else if(N400) begin
      mem_q[139] <= mem_n[139];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[138] <= 1'b0;
    end else if(N400) begin
      mem_q[138] <= mem_n[138];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[137] <= 1'b0;
    end else if(N400) begin
      mem_q[137] <= mem_n[137];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[136] <= 1'b0;
    end else if(N400) begin
      mem_q[136] <= mem_n[136];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[135] <= 1'b0;
    end else if(N400) begin
      mem_q[135] <= mem_n[135];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[134] <= 1'b0;
    end else if(N400) begin
      mem_q[134] <= mem_n[134];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[133] <= 1'b0;
    end else if(N400) begin
      mem_q[133] <= mem_n[133];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[132] <= 1'b0;
    end else if(N400) begin
      mem_q[132] <= mem_n[132];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[131] <= 1'b0;
    end else if(N400) begin
      mem_q[131] <= mem_n[131];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[130] <= 1'b0;
    end else if(N400) begin
      mem_q[130] <= mem_n[130];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[129] <= 1'b0;
    end else if(N400) begin
      mem_q[129] <= mem_n[129];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[128] <= 1'b0;
    end else if(N400) begin
      mem_q[128] <= mem_n[128];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[127] <= 1'b0;
    end else if(N400) begin
      mem_q[127] <= mem_n[127];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[126] <= 1'b0;
    end else if(N400) begin
      mem_q[126] <= mem_n[126];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[125] <= 1'b0;
    end else if(N400) begin
      mem_q[125] <= mem_n[125];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[124] <= 1'b0;
    end else if(N400) begin
      mem_q[124] <= mem_n[124];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[123] <= 1'b0;
    end else if(N400) begin
      mem_q[123] <= mem_n[123];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[122] <= 1'b0;
    end else if(N400) begin
      mem_q[122] <= mem_n[122];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[121] <= 1'b0;
    end else if(N400) begin
      mem_q[121] <= mem_n[121];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[120] <= 1'b0;
    end else if(N400) begin
      mem_q[120] <= mem_n[120];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[119] <= 1'b0;
    end else if(N400) begin
      mem_q[119] <= mem_n[119];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[118] <= 1'b0;
    end else if(N400) begin
      mem_q[118] <= mem_n[118];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[117] <= 1'b0;
    end else if(N400) begin
      mem_q[117] <= mem_n[117];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[116] <= 1'b0;
    end else if(N400) begin
      mem_q[116] <= mem_n[116];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[115] <= 1'b0;
    end else if(N400) begin
      mem_q[115] <= mem_n[115];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[114] <= 1'b0;
    end else if(N400) begin
      mem_q[114] <= mem_n[114];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[113] <= 1'b0;
    end else if(N400) begin
      mem_q[113] <= mem_n[113];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[112] <= 1'b0;
    end else if(N400) begin
      mem_q[112] <= mem_n[112];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[111] <= 1'b0;
    end else if(N400) begin
      mem_q[111] <= mem_n[111];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[110] <= 1'b0;
    end else if(N400) begin
      mem_q[110] <= mem_n[110];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[109] <= 1'b0;
    end else if(N400) begin
      mem_q[109] <= mem_n[109];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[108] <= 1'b0;
    end else if(N400) begin
      mem_q[108] <= mem_n[108];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[107] <= 1'b0;
    end else if(N400) begin
      mem_q[107] <= mem_n[107];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[106] <= 1'b0;
    end else if(N400) begin
      mem_q[106] <= mem_n[106];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[105] <= 1'b0;
    end else if(N400) begin
      mem_q[105] <= mem_n[105];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[104] <= 1'b0;
    end else if(N400) begin
      mem_q[104] <= mem_n[104];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[103] <= 1'b0;
    end else if(N400) begin
      mem_q[103] <= mem_n[103];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[102] <= 1'b0;
    end else if(N400) begin
      mem_q[102] <= mem_n[102];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[101] <= 1'b0;
    end else if(N400) begin
      mem_q[101] <= mem_n[101];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[100] <= 1'b0;
    end else if(N400) begin
      mem_q[100] <= mem_n[100];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[99] <= 1'b0;
    end else if(N400) begin
      mem_q[99] <= mem_n[99];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[98] <= 1'b0;
    end else if(N404) begin
      mem_q[98] <= mem_n[98];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[97] <= 1'b0;
    end else if(N404) begin
      mem_q[97] <= mem_n[97];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[96] <= 1'b0;
    end else if(N404) begin
      mem_q[96] <= mem_n[96];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[95] <= 1'b0;
    end else if(N404) begin
      mem_q[95] <= mem_n[95];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[94] <= 1'b0;
    end else if(N404) begin
      mem_q[94] <= mem_n[94];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[93] <= 1'b0;
    end else if(N404) begin
      mem_q[93] <= mem_n[93];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[92] <= 1'b0;
    end else if(N404) begin
      mem_q[92] <= mem_n[92];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[91] <= 1'b0;
    end else if(N404) begin
      mem_q[91] <= mem_n[91];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[90] <= 1'b0;
    end else if(N404) begin
      mem_q[90] <= mem_n[90];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[89] <= 1'b0;
    end else if(N404) begin
      mem_q[89] <= mem_n[89];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[88] <= 1'b0;
    end else if(N404) begin
      mem_q[88] <= mem_n[88];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[87] <= 1'b0;
    end else if(N404) begin
      mem_q[87] <= mem_n[87];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[86] <= 1'b0;
    end else if(N404) begin
      mem_q[86] <= mem_n[86];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[85] <= 1'b0;
    end else if(N404) begin
      mem_q[85] <= mem_n[85];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[84] <= 1'b0;
    end else if(N404) begin
      mem_q[84] <= mem_n[84];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[83] <= 1'b0;
    end else if(N404) begin
      mem_q[83] <= mem_n[83];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[82] <= 1'b0;
    end else if(N404) begin
      mem_q[82] <= mem_n[82];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[81] <= 1'b0;
    end else if(N404) begin
      mem_q[81] <= mem_n[81];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[80] <= 1'b0;
    end else if(N404) begin
      mem_q[80] <= mem_n[80];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[79] <= 1'b0;
    end else if(N404) begin
      mem_q[79] <= mem_n[79];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[78] <= 1'b0;
    end else if(N404) begin
      mem_q[78] <= mem_n[78];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[77] <= 1'b0;
    end else if(N404) begin
      mem_q[77] <= mem_n[77];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[76] <= 1'b0;
    end else if(N404) begin
      mem_q[76] <= mem_n[76];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[75] <= 1'b0;
    end else if(N404) begin
      mem_q[75] <= mem_n[75];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[74] <= 1'b0;
    end else if(N404) begin
      mem_q[74] <= mem_n[74];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[73] <= 1'b0;
    end else if(N404) begin
      mem_q[73] <= mem_n[73];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[72] <= 1'b0;
    end else if(N404) begin
      mem_q[72] <= mem_n[72];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[71] <= 1'b0;
    end else if(N404) begin
      mem_q[71] <= mem_n[71];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[70] <= 1'b0;
    end else if(N404) begin
      mem_q[70] <= mem_n[70];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[69] <= 1'b0;
    end else if(N404) begin
      mem_q[69] <= mem_n[69];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[68] <= 1'b0;
    end else if(N404) begin
      mem_q[68] <= mem_n[68];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[67] <= 1'b0;
    end else if(N404) begin
      mem_q[67] <= mem_n[67];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[66] <= 1'b0;
    end else if(N404) begin
      mem_q[66] <= mem_n[66];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[65] <= 1'b0;
    end else if(N404) begin
      mem_q[65] <= mem_n[65];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[64] <= 1'b0;
    end else if(N404) begin
      mem_q[64] <= mem_n[64];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[63] <= 1'b0;
    end else if(N404) begin
      mem_q[63] <= mem_n[63];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[62] <= 1'b0;
    end else if(N404) begin
      mem_q[62] <= mem_n[62];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[61] <= 1'b0;
    end else if(N404) begin
      mem_q[61] <= mem_n[61];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[60] <= 1'b0;
    end else if(N404) begin
      mem_q[60] <= mem_n[60];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[59] <= 1'b0;
    end else if(N404) begin
      mem_q[59] <= mem_n[59];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[58] <= 1'b0;
    end else if(N404) begin
      mem_q[58] <= mem_n[58];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[57] <= 1'b0;
    end else if(N404) begin
      mem_q[57] <= mem_n[57];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[56] <= 1'b0;
    end else if(N404) begin
      mem_q[56] <= mem_n[56];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[55] <= 1'b0;
    end else if(N404) begin
      mem_q[55] <= mem_n[55];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[54] <= 1'b0;
    end else if(N404) begin
      mem_q[54] <= mem_n[54];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[53] <= 1'b0;
    end else if(N404) begin
      mem_q[53] <= mem_n[53];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[52] <= 1'b0;
    end else if(N404) begin
      mem_q[52] <= mem_n[52];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[51] <= 1'b0;
    end else if(N404) begin
      mem_q[51] <= mem_n[51];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[50] <= 1'b0;
    end else if(N404) begin
      mem_q[50] <= mem_n[50];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[49] <= 1'b0;
    end else if(N407) begin
      mem_q[49] <= mem_n[49];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[48] <= 1'b0;
    end else if(N410) begin
      mem_q[48] <= mem_n[48];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[47] <= 1'b0;
    end else if(N410) begin
      mem_q[47] <= mem_n[47];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[46] <= 1'b0;
    end else if(N410) begin
      mem_q[46] <= mem_n[46];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[45] <= 1'b0;
    end else if(N410) begin
      mem_q[45] <= mem_n[45];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[44] <= 1'b0;
    end else if(N410) begin
      mem_q[44] <= mem_n[44];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[43] <= 1'b0;
    end else if(N410) begin
      mem_q[43] <= mem_n[43];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[42] <= 1'b0;
    end else if(N410) begin
      mem_q[42] <= mem_n[42];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[41] <= 1'b0;
    end else if(N410) begin
      mem_q[41] <= mem_n[41];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[40] <= 1'b0;
    end else if(N410) begin
      mem_q[40] <= mem_n[40];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[39] <= 1'b0;
    end else if(N410) begin
      mem_q[39] <= mem_n[39];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[38] <= 1'b0;
    end else if(N410) begin
      mem_q[38] <= mem_n[38];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[37] <= 1'b0;
    end else if(N410) begin
      mem_q[37] <= mem_n[37];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[36] <= 1'b0;
    end else if(N410) begin
      mem_q[36] <= mem_n[36];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[35] <= 1'b0;
    end else if(N410) begin
      mem_q[35] <= mem_n[35];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[34] <= 1'b0;
    end else if(N410) begin
      mem_q[34] <= mem_n[34];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[33] <= 1'b0;
    end else if(N410) begin
      mem_q[33] <= mem_n[33];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[32] <= 1'b0;
    end else if(N410) begin
      mem_q[32] <= mem_n[32];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[31] <= 1'b0;
    end else if(N410) begin
      mem_q[31] <= mem_n[31];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[30] <= 1'b0;
    end else if(N410) begin
      mem_q[30] <= mem_n[30];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[29] <= 1'b0;
    end else if(N410) begin
      mem_q[29] <= mem_n[29];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[28] <= 1'b0;
    end else if(N410) begin
      mem_q[28] <= mem_n[28];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[27] <= 1'b0;
    end else if(N410) begin
      mem_q[27] <= mem_n[27];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[26] <= 1'b0;
    end else if(N410) begin
      mem_q[26] <= mem_n[26];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[25] <= 1'b0;
    end else if(N410) begin
      mem_q[25] <= mem_n[25];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[24] <= 1'b0;
    end else if(N410) begin
      mem_q[24] <= mem_n[24];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[23] <= 1'b0;
    end else if(N410) begin
      mem_q[23] <= mem_n[23];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[22] <= 1'b0;
    end else if(N410) begin
      mem_q[22] <= mem_n[22];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[21] <= 1'b0;
    end else if(N410) begin
      mem_q[21] <= mem_n[21];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[20] <= 1'b0;
    end else if(N410) begin
      mem_q[20] <= mem_n[20];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[19] <= 1'b0;
    end else if(N410) begin
      mem_q[19] <= mem_n[19];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[18] <= 1'b0;
    end else if(N410) begin
      mem_q[18] <= mem_n[18];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[17] <= 1'b0;
    end else if(N410) begin
      mem_q[17] <= mem_n[17];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[16] <= 1'b0;
    end else if(N410) begin
      mem_q[16] <= mem_n[16];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[15] <= 1'b0;
    end else if(N410) begin
      mem_q[15] <= mem_n[15];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[14] <= 1'b0;
    end else if(N410) begin
      mem_q[14] <= mem_n[14];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[13] <= 1'b0;
    end else if(N410) begin
      mem_q[13] <= mem_n[13];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[12] <= 1'b0;
    end else if(N410) begin
      mem_q[12] <= mem_n[12];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[11] <= 1'b0;
    end else if(N410) begin
      mem_q[11] <= mem_n[11];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[10] <= 1'b0;
    end else if(N410) begin
      mem_q[10] <= mem_n[10];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[9] <= 1'b0;
    end else if(N410) begin
      mem_q[9] <= mem_n[9];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[8] <= 1'b0;
    end else if(N410) begin
      mem_q[8] <= mem_n[8];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[7] <= 1'b0;
    end else if(N410) begin
      mem_q[7] <= mem_n[7];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[6] <= 1'b0;
    end else if(N410) begin
      mem_q[6] <= mem_n[6];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[5] <= 1'b0;
    end else if(N410) begin
      mem_q[5] <= mem_n[5];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[4] <= 1'b0;
    end else if(N410) begin
      mem_q[4] <= mem_n[4];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[3] <= 1'b0;
    end else if(N410) begin
      mem_q[3] <= mem_n[3];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[2] <= 1'b0;
    end else if(N410) begin
      mem_q[2] <= mem_n[2];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[1] <= 1'b0;
    end else if(N410) begin
      mem_q[1] <= mem_n[1];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      mem_q[0] <= 1'b0;
    end else if(N410) begin
      mem_q[0] <= mem_n[0];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      status_cnt_q[1] <= 1'b0;
    end else if(1'b1) begin
      status_cnt_q[1] <= status_cnt_n[1];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      status_cnt_q[0] <= 1'b0;
    end else if(1'b1) begin
      status_cnt_q[0] <= status_cnt_n[0];
    end 
  end


  always @(posedge clk_i or posedge N357) begin
    if(N357) begin
      N17 <= 1'b0;
    end else if(N412) begin
      N17 <= write_pointer_n;
    end 
  end

  assign N413 = status_cnt_q[0] | status_cnt_q[1];
  assign ready_o = ~N413;
  assign N32 = N41 ^ 1'b1;
  assign N21 = N17 ^ 1'b1;
  assign { N23, N22 } = status_cnt_q + 1'b1;
  assign N45 = N35 ^ 1'b1;
  assign { N37, N36 } = { N27, N26 } - pop_ld_i;
  assign { N50, N49 } = { N37, N36 } - pop_st_i;
  assign N16 = ~N17;
  assign N40 = ~N41;
  assign N18 = (N1)? lsu_req_i[150] : 
               (N2)? mem_q[150] : 1'b0;
  assign N1 = N16;
  assign N2 = N17;
  assign N20 = (N2)? lsu_req_i[150] : 
               (N19)? mem_q[301] : 1'b0;
  assign { N25, N24 } = (N3)? { N20, N18 } : 
                        (N4)? { mem_q[301:301], mem_q[150:150] } : 1'b0;
  assign N3 = lus_req_valid_i;
  assign N4 = N15;
  assign { N27, N26 } = (N3)? { N23, N22 } : 
                        (N4)? status_cnt_q : 1'b0;
  assign N30 = (N5)? 1'b0 : 
               (N0)? N24 : 1'b0;
  assign N5 = N40;
  assign N31 = (N0)? 1'b0 : 
               (N43)? N25 : 1'b0;
  assign { N34, N33 } = (N6)? { N31, N30 } : 
                        (N7)? { N25, N24 } : 1'b0;
  assign N6 = pop_ld_i;
  assign N7 = N28;
  assign N35 = (N6)? N32 : 
               (N7)? N41 : 1'b0;
  assign N42 = (N5)? 1'b0 : 
               (N0)? N33 : 1'b0;
  assign N44 = (N0)? 1'b0 : 
               (N43)? N34 : 1'b0;
  assign { N47, N46 } = (N8)? { N44, N42 } : 
                        (N9)? { N34, N33 } : 1'b0;
  assign N8 = pop_st_i;
  assign N9 = N38;
  assign N48 = (N8)? N45 : 
               (N9)? N35 : 1'b0;
  assign { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53 } = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               (N52)? { N47, N46, lsu_req_i[149:0] } : 1'b0;
  assign N10 = N51;
  assign status_cnt_n = (N11)? { 1'b0, 1'b0 } : 
                        (N12)? { N50, N49 } : 1'b0;
  assign N11 = flush_i;
  assign N12 = N205;
  assign write_pointer_n = (N11)? 1'b0 : 
                           (N12)? N21 : 1'b0;
  assign read_pointer_n = (N11)? 1'b0 : 
                          (N12)? N48 : 1'b0;
  assign mem_n = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N12)? { N204, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53 } : 1'b0;
  assign lsu_ctrl_o = (N13)? lsu_req_i : 
                      (N14)? { N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356 } : 1'b0;
  assign N13 = ready_o;
  assign N14 = N413;
  assign N15 = ~lus_req_valid_i;
  assign N19 = ~N17;
  assign N28 = ~pop_ld_i;
  assign N29 = pop_ld_i;
  assign N38 = ~pop_st_i;
  assign N39 = pop_st_i;
  assign N43 = ~N41;
  assign N51 = pop_st_i & pop_ld_i;
  assign N52 = ~N51;
  assign N205 = ~flush_i;
  assign N357 = ~rst_ni;
  assign N358 = N52 & N205;
  assign N359 = lus_req_valid_i & N358;
  assign N360 = N19 & N359;
  assign N361 = N52 & N205;
  assign N362 = N15 & N361;
  assign N363 = N360 | N362;
  assign N364 = ~N363;
  assign N365 = N52 & N205;
  assign N366 = lus_req_valid_i & N365;
  assign N367 = N19 & N366;
  assign N368 = N52 & N205;
  assign N369 = N15 & N368;
  assign N370 = N367 | N369;
  assign N371 = ~N370;
  assign N372 = N52 & N205;
  assign N373 = lus_req_valid_i & N372;
  assign N374 = N19 & N373;
  assign N375 = N52 & N205;
  assign N376 = N15 & N375;
  assign N377 = N374 | N376;
  assign N378 = ~N377;
  assign N379 = lus_req_valid_i & N375;
  assign N380 = N19 & N379;
  assign N381 = N380 | N376;
  assign N382 = ~N381;
  assign N383 = N15 & N372;
  assign N384 = N380 | N383;
  assign N385 = ~N384;
  assign N386 = N374 | N383;
  assign N387 = ~N386;
  assign N388 = lus_req_valid_i & N368;
  assign N389 = N19 & N388;
  assign N390 = N389 | N369;
  assign N391 = ~N390;
  assign N392 = N17 & N388;
  assign N393 = N392 | N369;
  assign N394 = ~N393;
  assign N395 = N15 & N365;
  assign N396 = N392 | N395;
  assign N397 = ~N396;
  assign N398 = N17 & N366;
  assign N399 = N398 | N395;
  assign N400 = ~N399;
  assign N401 = lus_req_valid_i & N361;
  assign N402 = N17 & N401;
  assign N403 = N402 | N362;
  assign N404 = ~N403;
  assign N405 = N15 & N358;
  assign N406 = N402 | N405;
  assign N407 = ~N406;
  assign N408 = N17 & N359;
  assign N409 = N408 | N405;
  assign N410 = ~N409;
  assign N411 = N15 & N205;
  assign N412 = ~N411;

endmodule