module bsg_cache_sbuf_queue_width_p115
(
  clk_i,
  data_i,
  el0_en_i,
  el1_en_i,
  mux0_sel_i,
  mux1_sel_i,
  el0_snoop_o,
  el1_snoop_o,
  data_o
);

  input [114:0] data_i;
  output [114:0] el0_snoop_o;
  output [114:0] el1_snoop_o;
  output [114:0] data_o;
  input clk_i;
  input el0_en_i;
  input el1_en_i;
  input mux0_sel_i;
  input mux1_sel_i;
  wire [114:0] el0_snoop_o,el1_snoop_o,data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120;
  reg el0_snoop_o_114_sv2v_reg,el0_snoop_o_113_sv2v_reg,el0_snoop_o_112_sv2v_reg,
  el0_snoop_o_111_sv2v_reg,el0_snoop_o_110_sv2v_reg,el0_snoop_o_109_sv2v_reg,
  el0_snoop_o_108_sv2v_reg,el0_snoop_o_107_sv2v_reg,el0_snoop_o_106_sv2v_reg,
  el0_snoop_o_105_sv2v_reg,el0_snoop_o_104_sv2v_reg,el0_snoop_o_103_sv2v_reg,
  el0_snoop_o_102_sv2v_reg,el0_snoop_o_101_sv2v_reg,el0_snoop_o_100_sv2v_reg,el0_snoop_o_99_sv2v_reg,
  el0_snoop_o_98_sv2v_reg,el0_snoop_o_97_sv2v_reg,el0_snoop_o_96_sv2v_reg,
  el0_snoop_o_95_sv2v_reg,el0_snoop_o_94_sv2v_reg,el0_snoop_o_93_sv2v_reg,
  el0_snoop_o_92_sv2v_reg,el0_snoop_o_91_sv2v_reg,el0_snoop_o_90_sv2v_reg,el0_snoop_o_89_sv2v_reg,
  el0_snoop_o_88_sv2v_reg,el0_snoop_o_87_sv2v_reg,el0_snoop_o_86_sv2v_reg,
  el0_snoop_o_85_sv2v_reg,el0_snoop_o_84_sv2v_reg,el0_snoop_o_83_sv2v_reg,
  el0_snoop_o_82_sv2v_reg,el0_snoop_o_81_sv2v_reg,el0_snoop_o_80_sv2v_reg,el0_snoop_o_79_sv2v_reg,
  el0_snoop_o_78_sv2v_reg,el0_snoop_o_77_sv2v_reg,el0_snoop_o_76_sv2v_reg,
  el0_snoop_o_75_sv2v_reg,el0_snoop_o_74_sv2v_reg,el0_snoop_o_73_sv2v_reg,
  el0_snoop_o_72_sv2v_reg,el0_snoop_o_71_sv2v_reg,el0_snoop_o_70_sv2v_reg,el0_snoop_o_69_sv2v_reg,
  el0_snoop_o_68_sv2v_reg,el0_snoop_o_67_sv2v_reg,el0_snoop_o_66_sv2v_reg,
  el0_snoop_o_65_sv2v_reg,el0_snoop_o_64_sv2v_reg,el0_snoop_o_63_sv2v_reg,
  el0_snoop_o_62_sv2v_reg,el0_snoop_o_61_sv2v_reg,el0_snoop_o_60_sv2v_reg,el0_snoop_o_59_sv2v_reg,
  el0_snoop_o_58_sv2v_reg,el0_snoop_o_57_sv2v_reg,el0_snoop_o_56_sv2v_reg,
  el0_snoop_o_55_sv2v_reg,el0_snoop_o_54_sv2v_reg,el0_snoop_o_53_sv2v_reg,
  el0_snoop_o_52_sv2v_reg,el0_snoop_o_51_sv2v_reg,el0_snoop_o_50_sv2v_reg,el0_snoop_o_49_sv2v_reg,
  el0_snoop_o_48_sv2v_reg,el0_snoop_o_47_sv2v_reg,el0_snoop_o_46_sv2v_reg,
  el0_snoop_o_45_sv2v_reg,el0_snoop_o_44_sv2v_reg,el0_snoop_o_43_sv2v_reg,
  el0_snoop_o_42_sv2v_reg,el0_snoop_o_41_sv2v_reg,el0_snoop_o_40_sv2v_reg,el0_snoop_o_39_sv2v_reg,
  el0_snoop_o_38_sv2v_reg,el0_snoop_o_37_sv2v_reg,el0_snoop_o_36_sv2v_reg,
  el0_snoop_o_35_sv2v_reg,el0_snoop_o_34_sv2v_reg,el0_snoop_o_33_sv2v_reg,
  el0_snoop_o_32_sv2v_reg,el0_snoop_o_31_sv2v_reg,el0_snoop_o_30_sv2v_reg,el0_snoop_o_29_sv2v_reg,
  el0_snoop_o_28_sv2v_reg,el0_snoop_o_27_sv2v_reg,el0_snoop_o_26_sv2v_reg,
  el0_snoop_o_25_sv2v_reg,el0_snoop_o_24_sv2v_reg,el0_snoop_o_23_sv2v_reg,
  el0_snoop_o_22_sv2v_reg,el0_snoop_o_21_sv2v_reg,el0_snoop_o_20_sv2v_reg,el0_snoop_o_19_sv2v_reg,
  el0_snoop_o_18_sv2v_reg,el0_snoop_o_17_sv2v_reg,el0_snoop_o_16_sv2v_reg,
  el0_snoop_o_15_sv2v_reg,el0_snoop_o_14_sv2v_reg,el0_snoop_o_13_sv2v_reg,
  el0_snoop_o_12_sv2v_reg,el0_snoop_o_11_sv2v_reg,el0_snoop_o_10_sv2v_reg,el0_snoop_o_9_sv2v_reg,
  el0_snoop_o_8_sv2v_reg,el0_snoop_o_7_sv2v_reg,el0_snoop_o_6_sv2v_reg,
  el0_snoop_o_5_sv2v_reg,el0_snoop_o_4_sv2v_reg,el0_snoop_o_3_sv2v_reg,el0_snoop_o_2_sv2v_reg,
  el0_snoop_o_1_sv2v_reg,el0_snoop_o_0_sv2v_reg,el1_snoop_o_114_sv2v_reg,
  el1_snoop_o_113_sv2v_reg,el1_snoop_o_112_sv2v_reg,el1_snoop_o_111_sv2v_reg,
  el1_snoop_o_110_sv2v_reg,el1_snoop_o_109_sv2v_reg,el1_snoop_o_108_sv2v_reg,
  el1_snoop_o_107_sv2v_reg,el1_snoop_o_106_sv2v_reg,el1_snoop_o_105_sv2v_reg,el1_snoop_o_104_sv2v_reg,
  el1_snoop_o_103_sv2v_reg,el1_snoop_o_102_sv2v_reg,el1_snoop_o_101_sv2v_reg,
  el1_snoop_o_100_sv2v_reg,el1_snoop_o_99_sv2v_reg,el1_snoop_o_98_sv2v_reg,
  el1_snoop_o_97_sv2v_reg,el1_snoop_o_96_sv2v_reg,el1_snoop_o_95_sv2v_reg,
  el1_snoop_o_94_sv2v_reg,el1_snoop_o_93_sv2v_reg,el1_snoop_o_92_sv2v_reg,el1_snoop_o_91_sv2v_reg,
  el1_snoop_o_90_sv2v_reg,el1_snoop_o_89_sv2v_reg,el1_snoop_o_88_sv2v_reg,
  el1_snoop_o_87_sv2v_reg,el1_snoop_o_86_sv2v_reg,el1_snoop_o_85_sv2v_reg,
  el1_snoop_o_84_sv2v_reg,el1_snoop_o_83_sv2v_reg,el1_snoop_o_82_sv2v_reg,el1_snoop_o_81_sv2v_reg,
  el1_snoop_o_80_sv2v_reg,el1_snoop_o_79_sv2v_reg,el1_snoop_o_78_sv2v_reg,
  el1_snoop_o_77_sv2v_reg,el1_snoop_o_76_sv2v_reg,el1_snoop_o_75_sv2v_reg,
  el1_snoop_o_74_sv2v_reg,el1_snoop_o_73_sv2v_reg,el1_snoop_o_72_sv2v_reg,el1_snoop_o_71_sv2v_reg,
  el1_snoop_o_70_sv2v_reg,el1_snoop_o_69_sv2v_reg,el1_snoop_o_68_sv2v_reg,
  el1_snoop_o_67_sv2v_reg,el1_snoop_o_66_sv2v_reg,el1_snoop_o_65_sv2v_reg,
  el1_snoop_o_64_sv2v_reg,el1_snoop_o_63_sv2v_reg,el1_snoop_o_62_sv2v_reg,el1_snoop_o_61_sv2v_reg,
  el1_snoop_o_60_sv2v_reg,el1_snoop_o_59_sv2v_reg,el1_snoop_o_58_sv2v_reg,
  el1_snoop_o_57_sv2v_reg,el1_snoop_o_56_sv2v_reg,el1_snoop_o_55_sv2v_reg,
  el1_snoop_o_54_sv2v_reg,el1_snoop_o_53_sv2v_reg,el1_snoop_o_52_sv2v_reg,el1_snoop_o_51_sv2v_reg,
  el1_snoop_o_50_sv2v_reg,el1_snoop_o_49_sv2v_reg,el1_snoop_o_48_sv2v_reg,
  el1_snoop_o_47_sv2v_reg,el1_snoop_o_46_sv2v_reg,el1_snoop_o_45_sv2v_reg,
  el1_snoop_o_44_sv2v_reg,el1_snoop_o_43_sv2v_reg,el1_snoop_o_42_sv2v_reg,el1_snoop_o_41_sv2v_reg,
  el1_snoop_o_40_sv2v_reg,el1_snoop_o_39_sv2v_reg,el1_snoop_o_38_sv2v_reg,
  el1_snoop_o_37_sv2v_reg,el1_snoop_o_36_sv2v_reg,el1_snoop_o_35_sv2v_reg,
  el1_snoop_o_34_sv2v_reg,el1_snoop_o_33_sv2v_reg,el1_snoop_o_32_sv2v_reg,el1_snoop_o_31_sv2v_reg,
  el1_snoop_o_30_sv2v_reg,el1_snoop_o_29_sv2v_reg,el1_snoop_o_28_sv2v_reg,
  el1_snoop_o_27_sv2v_reg,el1_snoop_o_26_sv2v_reg,el1_snoop_o_25_sv2v_reg,
  el1_snoop_o_24_sv2v_reg,el1_snoop_o_23_sv2v_reg,el1_snoop_o_22_sv2v_reg,el1_snoop_o_21_sv2v_reg,
  el1_snoop_o_20_sv2v_reg,el1_snoop_o_19_sv2v_reg,el1_snoop_o_18_sv2v_reg,
  el1_snoop_o_17_sv2v_reg,el1_snoop_o_16_sv2v_reg,el1_snoop_o_15_sv2v_reg,
  el1_snoop_o_14_sv2v_reg,el1_snoop_o_13_sv2v_reg,el1_snoop_o_12_sv2v_reg,el1_snoop_o_11_sv2v_reg,
  el1_snoop_o_10_sv2v_reg,el1_snoop_o_9_sv2v_reg,el1_snoop_o_8_sv2v_reg,
  el1_snoop_o_7_sv2v_reg,el1_snoop_o_6_sv2v_reg,el1_snoop_o_5_sv2v_reg,el1_snoop_o_4_sv2v_reg,
  el1_snoop_o_3_sv2v_reg,el1_snoop_o_2_sv2v_reg,el1_snoop_o_1_sv2v_reg,
  el1_snoop_o_0_sv2v_reg;
  assign el0_snoop_o[114] = el0_snoop_o_114_sv2v_reg;
  assign el0_snoop_o[113] = el0_snoop_o_113_sv2v_reg;
  assign el0_snoop_o[112] = el0_snoop_o_112_sv2v_reg;
  assign el0_snoop_o[111] = el0_snoop_o_111_sv2v_reg;
  assign el0_snoop_o[110] = el0_snoop_o_110_sv2v_reg;
  assign el0_snoop_o[109] = el0_snoop_o_109_sv2v_reg;
  assign el0_snoop_o[108] = el0_snoop_o_108_sv2v_reg;
  assign el0_snoop_o[107] = el0_snoop_o_107_sv2v_reg;
  assign el0_snoop_o[106] = el0_snoop_o_106_sv2v_reg;
  assign el0_snoop_o[105] = el0_snoop_o_105_sv2v_reg;
  assign el0_snoop_o[104] = el0_snoop_o_104_sv2v_reg;
  assign el0_snoop_o[103] = el0_snoop_o_103_sv2v_reg;
  assign el0_snoop_o[102] = el0_snoop_o_102_sv2v_reg;
  assign el0_snoop_o[101] = el0_snoop_o_101_sv2v_reg;
  assign el0_snoop_o[100] = el0_snoop_o_100_sv2v_reg;
  assign el0_snoop_o[99] = el0_snoop_o_99_sv2v_reg;
  assign el0_snoop_o[98] = el0_snoop_o_98_sv2v_reg;
  assign el0_snoop_o[97] = el0_snoop_o_97_sv2v_reg;
  assign el0_snoop_o[96] = el0_snoop_o_96_sv2v_reg;
  assign el0_snoop_o[95] = el0_snoop_o_95_sv2v_reg;
  assign el0_snoop_o[94] = el0_snoop_o_94_sv2v_reg;
  assign el0_snoop_o[93] = el0_snoop_o_93_sv2v_reg;
  assign el0_snoop_o[92] = el0_snoop_o_92_sv2v_reg;
  assign el0_snoop_o[91] = el0_snoop_o_91_sv2v_reg;
  assign el0_snoop_o[90] = el0_snoop_o_90_sv2v_reg;
  assign el0_snoop_o[89] = el0_snoop_o_89_sv2v_reg;
  assign el0_snoop_o[88] = el0_snoop_o_88_sv2v_reg;
  assign el0_snoop_o[87] = el0_snoop_o_87_sv2v_reg;
  assign el0_snoop_o[86] = el0_snoop_o_86_sv2v_reg;
  assign el0_snoop_o[85] = el0_snoop_o_85_sv2v_reg;
  assign el0_snoop_o[84] = el0_snoop_o_84_sv2v_reg;
  assign el0_snoop_o[83] = el0_snoop_o_83_sv2v_reg;
  assign el0_snoop_o[82] = el0_snoop_o_82_sv2v_reg;
  assign el0_snoop_o[81] = el0_snoop_o_81_sv2v_reg;
  assign el0_snoop_o[80] = el0_snoop_o_80_sv2v_reg;
  assign el0_snoop_o[79] = el0_snoop_o_79_sv2v_reg;
  assign el0_snoop_o[78] = el0_snoop_o_78_sv2v_reg;
  assign el0_snoop_o[77] = el0_snoop_o_77_sv2v_reg;
  assign el0_snoop_o[76] = el0_snoop_o_76_sv2v_reg;
  assign el0_snoop_o[75] = el0_snoop_o_75_sv2v_reg;
  assign el0_snoop_o[74] = el0_snoop_o_74_sv2v_reg;
  assign el0_snoop_o[73] = el0_snoop_o_73_sv2v_reg;
  assign el0_snoop_o[72] = el0_snoop_o_72_sv2v_reg;
  assign el0_snoop_o[71] = el0_snoop_o_71_sv2v_reg;
  assign el0_snoop_o[70] = el0_snoop_o_70_sv2v_reg;
  assign el0_snoop_o[69] = el0_snoop_o_69_sv2v_reg;
  assign el0_snoop_o[68] = el0_snoop_o_68_sv2v_reg;
  assign el0_snoop_o[67] = el0_snoop_o_67_sv2v_reg;
  assign el0_snoop_o[66] = el0_snoop_o_66_sv2v_reg;
  assign el0_snoop_o[65] = el0_snoop_o_65_sv2v_reg;
  assign el0_snoop_o[64] = el0_snoop_o_64_sv2v_reg;
  assign el0_snoop_o[63] = el0_snoop_o_63_sv2v_reg;
  assign el0_snoop_o[62] = el0_snoop_o_62_sv2v_reg;
  assign el0_snoop_o[61] = el0_snoop_o_61_sv2v_reg;
  assign el0_snoop_o[60] = el0_snoop_o_60_sv2v_reg;
  assign el0_snoop_o[59] = el0_snoop_o_59_sv2v_reg;
  assign el0_snoop_o[58] = el0_snoop_o_58_sv2v_reg;
  assign el0_snoop_o[57] = el0_snoop_o_57_sv2v_reg;
  assign el0_snoop_o[56] = el0_snoop_o_56_sv2v_reg;
  assign el0_snoop_o[55] = el0_snoop_o_55_sv2v_reg;
  assign el0_snoop_o[54] = el0_snoop_o_54_sv2v_reg;
  assign el0_snoop_o[53] = el0_snoop_o_53_sv2v_reg;
  assign el0_snoop_o[52] = el0_snoop_o_52_sv2v_reg;
  assign el0_snoop_o[51] = el0_snoop_o_51_sv2v_reg;
  assign el0_snoop_o[50] = el0_snoop_o_50_sv2v_reg;
  assign el0_snoop_o[49] = el0_snoop_o_49_sv2v_reg;
  assign el0_snoop_o[48] = el0_snoop_o_48_sv2v_reg;
  assign el0_snoop_o[47] = el0_snoop_o_47_sv2v_reg;
  assign el0_snoop_o[46] = el0_snoop_o_46_sv2v_reg;
  assign el0_snoop_o[45] = el0_snoop_o_45_sv2v_reg;
  assign el0_snoop_o[44] = el0_snoop_o_44_sv2v_reg;
  assign el0_snoop_o[43] = el0_snoop_o_43_sv2v_reg;
  assign el0_snoop_o[42] = el0_snoop_o_42_sv2v_reg;
  assign el0_snoop_o[41] = el0_snoop_o_41_sv2v_reg;
  assign el0_snoop_o[40] = el0_snoop_o_40_sv2v_reg;
  assign el0_snoop_o[39] = el0_snoop_o_39_sv2v_reg;
  assign el0_snoop_o[38] = el0_snoop_o_38_sv2v_reg;
  assign el0_snoop_o[37] = el0_snoop_o_37_sv2v_reg;
  assign el0_snoop_o[36] = el0_snoop_o_36_sv2v_reg;
  assign el0_snoop_o[35] = el0_snoop_o_35_sv2v_reg;
  assign el0_snoop_o[34] = el0_snoop_o_34_sv2v_reg;
  assign el0_snoop_o[33] = el0_snoop_o_33_sv2v_reg;
  assign el0_snoop_o[32] = el0_snoop_o_32_sv2v_reg;
  assign el0_snoop_o[31] = el0_snoop_o_31_sv2v_reg;
  assign el0_snoop_o[30] = el0_snoop_o_30_sv2v_reg;
  assign el0_snoop_o[29] = el0_snoop_o_29_sv2v_reg;
  assign el0_snoop_o[28] = el0_snoop_o_28_sv2v_reg;
  assign el0_snoop_o[27] = el0_snoop_o_27_sv2v_reg;
  assign el0_snoop_o[26] = el0_snoop_o_26_sv2v_reg;
  assign el0_snoop_o[25] = el0_snoop_o_25_sv2v_reg;
  assign el0_snoop_o[24] = el0_snoop_o_24_sv2v_reg;
  assign el0_snoop_o[23] = el0_snoop_o_23_sv2v_reg;
  assign el0_snoop_o[22] = el0_snoop_o_22_sv2v_reg;
  assign el0_snoop_o[21] = el0_snoop_o_21_sv2v_reg;
  assign el0_snoop_o[20] = el0_snoop_o_20_sv2v_reg;
  assign el0_snoop_o[19] = el0_snoop_o_19_sv2v_reg;
  assign el0_snoop_o[18] = el0_snoop_o_18_sv2v_reg;
  assign el0_snoop_o[17] = el0_snoop_o_17_sv2v_reg;
  assign el0_snoop_o[16] = el0_snoop_o_16_sv2v_reg;
  assign el0_snoop_o[15] = el0_snoop_o_15_sv2v_reg;
  assign el0_snoop_o[14] = el0_snoop_o_14_sv2v_reg;
  assign el0_snoop_o[13] = el0_snoop_o_13_sv2v_reg;
  assign el0_snoop_o[12] = el0_snoop_o_12_sv2v_reg;
  assign el0_snoop_o[11] = el0_snoop_o_11_sv2v_reg;
  assign el0_snoop_o[10] = el0_snoop_o_10_sv2v_reg;
  assign el0_snoop_o[9] = el0_snoop_o_9_sv2v_reg;
  assign el0_snoop_o[8] = el0_snoop_o_8_sv2v_reg;
  assign el0_snoop_o[7] = el0_snoop_o_7_sv2v_reg;
  assign el0_snoop_o[6] = el0_snoop_o_6_sv2v_reg;
  assign el0_snoop_o[5] = el0_snoop_o_5_sv2v_reg;
  assign el0_snoop_o[4] = el0_snoop_o_4_sv2v_reg;
  assign el0_snoop_o[3] = el0_snoop_o_3_sv2v_reg;
  assign el0_snoop_o[2] = el0_snoop_o_2_sv2v_reg;
  assign el0_snoop_o[1] = el0_snoop_o_1_sv2v_reg;
  assign el0_snoop_o[0] = el0_snoop_o_0_sv2v_reg;
  assign el1_snoop_o[114] = el1_snoop_o_114_sv2v_reg;
  assign el1_snoop_o[113] = el1_snoop_o_113_sv2v_reg;
  assign el1_snoop_o[112] = el1_snoop_o_112_sv2v_reg;
  assign el1_snoop_o[111] = el1_snoop_o_111_sv2v_reg;
  assign el1_snoop_o[110] = el1_snoop_o_110_sv2v_reg;
  assign el1_snoop_o[109] = el1_snoop_o_109_sv2v_reg;
  assign el1_snoop_o[108] = el1_snoop_o_108_sv2v_reg;
  assign el1_snoop_o[107] = el1_snoop_o_107_sv2v_reg;
  assign el1_snoop_o[106] = el1_snoop_o_106_sv2v_reg;
  assign el1_snoop_o[105] = el1_snoop_o_105_sv2v_reg;
  assign el1_snoop_o[104] = el1_snoop_o_104_sv2v_reg;
  assign el1_snoop_o[103] = el1_snoop_o_103_sv2v_reg;
  assign el1_snoop_o[102] = el1_snoop_o_102_sv2v_reg;
  assign el1_snoop_o[101] = el1_snoop_o_101_sv2v_reg;
  assign el1_snoop_o[100] = el1_snoop_o_100_sv2v_reg;
  assign el1_snoop_o[99] = el1_snoop_o_99_sv2v_reg;
  assign el1_snoop_o[98] = el1_snoop_o_98_sv2v_reg;
  assign el1_snoop_o[97] = el1_snoop_o_97_sv2v_reg;
  assign el1_snoop_o[96] = el1_snoop_o_96_sv2v_reg;
  assign el1_snoop_o[95] = el1_snoop_o_95_sv2v_reg;
  assign el1_snoop_o[94] = el1_snoop_o_94_sv2v_reg;
  assign el1_snoop_o[93] = el1_snoop_o_93_sv2v_reg;
  assign el1_snoop_o[92] = el1_snoop_o_92_sv2v_reg;
  assign el1_snoop_o[91] = el1_snoop_o_91_sv2v_reg;
  assign el1_snoop_o[90] = el1_snoop_o_90_sv2v_reg;
  assign el1_snoop_o[89] = el1_snoop_o_89_sv2v_reg;
  assign el1_snoop_o[88] = el1_snoop_o_88_sv2v_reg;
  assign el1_snoop_o[87] = el1_snoop_o_87_sv2v_reg;
  assign el1_snoop_o[86] = el1_snoop_o_86_sv2v_reg;
  assign el1_snoop_o[85] = el1_snoop_o_85_sv2v_reg;
  assign el1_snoop_o[84] = el1_snoop_o_84_sv2v_reg;
  assign el1_snoop_o[83] = el1_snoop_o_83_sv2v_reg;
  assign el1_snoop_o[82] = el1_snoop_o_82_sv2v_reg;
  assign el1_snoop_o[81] = el1_snoop_o_81_sv2v_reg;
  assign el1_snoop_o[80] = el1_snoop_o_80_sv2v_reg;
  assign el1_snoop_o[79] = el1_snoop_o_79_sv2v_reg;
  assign el1_snoop_o[78] = el1_snoop_o_78_sv2v_reg;
  assign el1_snoop_o[77] = el1_snoop_o_77_sv2v_reg;
  assign el1_snoop_o[76] = el1_snoop_o_76_sv2v_reg;
  assign el1_snoop_o[75] = el1_snoop_o_75_sv2v_reg;
  assign el1_snoop_o[74] = el1_snoop_o_74_sv2v_reg;
  assign el1_snoop_o[73] = el1_snoop_o_73_sv2v_reg;
  assign el1_snoop_o[72] = el1_snoop_o_72_sv2v_reg;
  assign el1_snoop_o[71] = el1_snoop_o_71_sv2v_reg;
  assign el1_snoop_o[70] = el1_snoop_o_70_sv2v_reg;
  assign el1_snoop_o[69] = el1_snoop_o_69_sv2v_reg;
  assign el1_snoop_o[68] = el1_snoop_o_68_sv2v_reg;
  assign el1_snoop_o[67] = el1_snoop_o_67_sv2v_reg;
  assign el1_snoop_o[66] = el1_snoop_o_66_sv2v_reg;
  assign el1_snoop_o[65] = el1_snoop_o_65_sv2v_reg;
  assign el1_snoop_o[64] = el1_snoop_o_64_sv2v_reg;
  assign el1_snoop_o[63] = el1_snoop_o_63_sv2v_reg;
  assign el1_snoop_o[62] = el1_snoop_o_62_sv2v_reg;
  assign el1_snoop_o[61] = el1_snoop_o_61_sv2v_reg;
  assign el1_snoop_o[60] = el1_snoop_o_60_sv2v_reg;
  assign el1_snoop_o[59] = el1_snoop_o_59_sv2v_reg;
  assign el1_snoop_o[58] = el1_snoop_o_58_sv2v_reg;
  assign el1_snoop_o[57] = el1_snoop_o_57_sv2v_reg;
  assign el1_snoop_o[56] = el1_snoop_o_56_sv2v_reg;
  assign el1_snoop_o[55] = el1_snoop_o_55_sv2v_reg;
  assign el1_snoop_o[54] = el1_snoop_o_54_sv2v_reg;
  assign el1_snoop_o[53] = el1_snoop_o_53_sv2v_reg;
  assign el1_snoop_o[52] = el1_snoop_o_52_sv2v_reg;
  assign el1_snoop_o[51] = el1_snoop_o_51_sv2v_reg;
  assign el1_snoop_o[50] = el1_snoop_o_50_sv2v_reg;
  assign el1_snoop_o[49] = el1_snoop_o_49_sv2v_reg;
  assign el1_snoop_o[48] = el1_snoop_o_48_sv2v_reg;
  assign el1_snoop_o[47] = el1_snoop_o_47_sv2v_reg;
  assign el1_snoop_o[46] = el1_snoop_o_46_sv2v_reg;
  assign el1_snoop_o[45] = el1_snoop_o_45_sv2v_reg;
  assign el1_snoop_o[44] = el1_snoop_o_44_sv2v_reg;
  assign el1_snoop_o[43] = el1_snoop_o_43_sv2v_reg;
  assign el1_snoop_o[42] = el1_snoop_o_42_sv2v_reg;
  assign el1_snoop_o[41] = el1_snoop_o_41_sv2v_reg;
  assign el1_snoop_o[40] = el1_snoop_o_40_sv2v_reg;
  assign el1_snoop_o[39] = el1_snoop_o_39_sv2v_reg;
  assign el1_snoop_o[38] = el1_snoop_o_38_sv2v_reg;
  assign el1_snoop_o[37] = el1_snoop_o_37_sv2v_reg;
  assign el1_snoop_o[36] = el1_snoop_o_36_sv2v_reg;
  assign el1_snoop_o[35] = el1_snoop_o_35_sv2v_reg;
  assign el1_snoop_o[34] = el1_snoop_o_34_sv2v_reg;
  assign el1_snoop_o[33] = el1_snoop_o_33_sv2v_reg;
  assign el1_snoop_o[32] = el1_snoop_o_32_sv2v_reg;
  assign el1_snoop_o[31] = el1_snoop_o_31_sv2v_reg;
  assign el1_snoop_o[30] = el1_snoop_o_30_sv2v_reg;
  assign el1_snoop_o[29] = el1_snoop_o_29_sv2v_reg;
  assign el1_snoop_o[28] = el1_snoop_o_28_sv2v_reg;
  assign el1_snoop_o[27] = el1_snoop_o_27_sv2v_reg;
  assign el1_snoop_o[26] = el1_snoop_o_26_sv2v_reg;
  assign el1_snoop_o[25] = el1_snoop_o_25_sv2v_reg;
  assign el1_snoop_o[24] = el1_snoop_o_24_sv2v_reg;
  assign el1_snoop_o[23] = el1_snoop_o_23_sv2v_reg;
  assign el1_snoop_o[22] = el1_snoop_o_22_sv2v_reg;
  assign el1_snoop_o[21] = el1_snoop_o_21_sv2v_reg;
  assign el1_snoop_o[20] = el1_snoop_o_20_sv2v_reg;
  assign el1_snoop_o[19] = el1_snoop_o_19_sv2v_reg;
  assign el1_snoop_o[18] = el1_snoop_o_18_sv2v_reg;
  assign el1_snoop_o[17] = el1_snoop_o_17_sv2v_reg;
  assign el1_snoop_o[16] = el1_snoop_o_16_sv2v_reg;
  assign el1_snoop_o[15] = el1_snoop_o_15_sv2v_reg;
  assign el1_snoop_o[14] = el1_snoop_o_14_sv2v_reg;
  assign el1_snoop_o[13] = el1_snoop_o_13_sv2v_reg;
  assign el1_snoop_o[12] = el1_snoop_o_12_sv2v_reg;
  assign el1_snoop_o[11] = el1_snoop_o_11_sv2v_reg;
  assign el1_snoop_o[10] = el1_snoop_o_10_sv2v_reg;
  assign el1_snoop_o[9] = el1_snoop_o_9_sv2v_reg;
  assign el1_snoop_o[8] = el1_snoop_o_8_sv2v_reg;
  assign el1_snoop_o[7] = el1_snoop_o_7_sv2v_reg;
  assign el1_snoop_o[6] = el1_snoop_o_6_sv2v_reg;
  assign el1_snoop_o[5] = el1_snoop_o_5_sv2v_reg;
  assign el1_snoop_o[4] = el1_snoop_o_4_sv2v_reg;
  assign el1_snoop_o[3] = el1_snoop_o_3_sv2v_reg;
  assign el1_snoop_o[2] = el1_snoop_o_2_sv2v_reg;
  assign el1_snoop_o[1] = el1_snoop_o_1_sv2v_reg;
  assign el1_snoop_o[0] = el1_snoop_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_114_sv2v_reg <= data_i[114];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_113_sv2v_reg <= data_i[113];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_112_sv2v_reg <= data_i[112];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_111_sv2v_reg <= data_i[111];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_110_sv2v_reg <= data_i[110];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_109_sv2v_reg <= data_i[109];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_108_sv2v_reg <= data_i[108];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_107_sv2v_reg <= data_i[107];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_106_sv2v_reg <= data_i[106];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_105_sv2v_reg <= data_i[105];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_104_sv2v_reg <= data_i[104];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_103_sv2v_reg <= data_i[103];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_102_sv2v_reg <= data_i[102];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_101_sv2v_reg <= data_i[101];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_100_sv2v_reg <= data_i[100];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_99_sv2v_reg <= data_i[99];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_98_sv2v_reg <= data_i[98];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_97_sv2v_reg <= data_i[97];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_96_sv2v_reg <= data_i[96];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_95_sv2v_reg <= data_i[95];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_94_sv2v_reg <= data_i[94];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_93_sv2v_reg <= data_i[93];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_92_sv2v_reg <= data_i[92];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_91_sv2v_reg <= data_i[91];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_90_sv2v_reg <= data_i[90];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_89_sv2v_reg <= data_i[89];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_88_sv2v_reg <= data_i[88];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_87_sv2v_reg <= data_i[87];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_86_sv2v_reg <= data_i[86];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_85_sv2v_reg <= data_i[85];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_84_sv2v_reg <= data_i[84];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_83_sv2v_reg <= data_i[83];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_82_sv2v_reg <= data_i[82];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_81_sv2v_reg <= data_i[81];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_80_sv2v_reg <= data_i[80];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_79_sv2v_reg <= data_i[79];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_78_sv2v_reg <= data_i[78];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_77_sv2v_reg <= data_i[77];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_76_sv2v_reg <= data_i[76];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_75_sv2v_reg <= data_i[75];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_74_sv2v_reg <= data_i[74];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_73_sv2v_reg <= data_i[73];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_72_sv2v_reg <= data_i[72];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_71_sv2v_reg <= data_i[71];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_70_sv2v_reg <= data_i[70];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_69_sv2v_reg <= data_i[69];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_68_sv2v_reg <= data_i[68];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_67_sv2v_reg <= data_i[67];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_66_sv2v_reg <= data_i[66];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_65_sv2v_reg <= data_i[65];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_64_sv2v_reg <= data_i[64];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_63_sv2v_reg <= data_i[63];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_62_sv2v_reg <= data_i[62];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_61_sv2v_reg <= data_i[61];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_60_sv2v_reg <= data_i[60];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_59_sv2v_reg <= data_i[59];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_58_sv2v_reg <= data_i[58];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_57_sv2v_reg <= data_i[57];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_56_sv2v_reg <= data_i[56];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_55_sv2v_reg <= data_i[55];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_54_sv2v_reg <= data_i[54];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_53_sv2v_reg <= data_i[53];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_52_sv2v_reg <= data_i[52];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_51_sv2v_reg <= data_i[51];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_50_sv2v_reg <= data_i[50];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_49_sv2v_reg <= data_i[49];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_48_sv2v_reg <= data_i[48];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_47_sv2v_reg <= data_i[47];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_46_sv2v_reg <= data_i[46];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_45_sv2v_reg <= data_i[45];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_44_sv2v_reg <= data_i[44];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_43_sv2v_reg <= data_i[43];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_42_sv2v_reg <= data_i[42];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_41_sv2v_reg <= data_i[41];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_40_sv2v_reg <= data_i[40];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_39_sv2v_reg <= data_i[39];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_38_sv2v_reg <= data_i[38];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_37_sv2v_reg <= data_i[37];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_36_sv2v_reg <= data_i[36];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_35_sv2v_reg <= data_i[35];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_34_sv2v_reg <= data_i[34];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_33_sv2v_reg <= data_i[33];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_32_sv2v_reg <= data_i[32];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_31_sv2v_reg <= data_i[31];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_30_sv2v_reg <= data_i[30];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_29_sv2v_reg <= data_i[29];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_28_sv2v_reg <= data_i[28];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_27_sv2v_reg <= data_i[27];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_26_sv2v_reg <= data_i[26];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_25_sv2v_reg <= data_i[25];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_24_sv2v_reg <= data_i[24];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_23_sv2v_reg <= data_i[23];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_22_sv2v_reg <= data_i[22];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_21_sv2v_reg <= data_i[21];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_20_sv2v_reg <= data_i[20];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_19_sv2v_reg <= data_i[19];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_18_sv2v_reg <= data_i[18];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_17_sv2v_reg <= data_i[17];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_16_sv2v_reg <= data_i[16];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_15_sv2v_reg <= data_i[15];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_14_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_13_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_12_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_11_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_10_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_9_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_8_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_7_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_6_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_5_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_4_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_3_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_2_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_1_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(el0_en_i) begin
      el0_snoop_o_0_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_114_sv2v_reg <= N119;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_113_sv2v_reg <= N118;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_112_sv2v_reg <= N117;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_111_sv2v_reg <= N116;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_110_sv2v_reg <= N115;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_109_sv2v_reg <= N114;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_108_sv2v_reg <= N113;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_107_sv2v_reg <= N112;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_106_sv2v_reg <= N111;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_105_sv2v_reg <= N110;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_104_sv2v_reg <= N109;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_103_sv2v_reg <= N108;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_102_sv2v_reg <= N107;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_101_sv2v_reg <= N106;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_100_sv2v_reg <= N105;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_99_sv2v_reg <= N104;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_98_sv2v_reg <= N103;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_97_sv2v_reg <= N102;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_96_sv2v_reg <= N101;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_95_sv2v_reg <= N100;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_94_sv2v_reg <= N99;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_93_sv2v_reg <= N98;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_92_sv2v_reg <= N97;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_91_sv2v_reg <= N96;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_90_sv2v_reg <= N95;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_89_sv2v_reg <= N94;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_88_sv2v_reg <= N93;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_87_sv2v_reg <= N92;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_86_sv2v_reg <= N91;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_85_sv2v_reg <= N90;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_84_sv2v_reg <= N89;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_83_sv2v_reg <= N88;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_82_sv2v_reg <= N87;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_81_sv2v_reg <= N86;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_80_sv2v_reg <= N85;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_79_sv2v_reg <= N84;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_78_sv2v_reg <= N83;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_77_sv2v_reg <= N82;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_76_sv2v_reg <= N81;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_75_sv2v_reg <= N80;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_74_sv2v_reg <= N79;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_73_sv2v_reg <= N78;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_72_sv2v_reg <= N77;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_71_sv2v_reg <= N76;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_70_sv2v_reg <= N75;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_69_sv2v_reg <= N74;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_68_sv2v_reg <= N73;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_67_sv2v_reg <= N72;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_66_sv2v_reg <= N71;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_65_sv2v_reg <= N70;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_64_sv2v_reg <= N69;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_63_sv2v_reg <= N68;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_62_sv2v_reg <= N67;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_61_sv2v_reg <= N66;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_60_sv2v_reg <= N65;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_59_sv2v_reg <= N64;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_58_sv2v_reg <= N63;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_57_sv2v_reg <= N62;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_56_sv2v_reg <= N61;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_55_sv2v_reg <= N60;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_54_sv2v_reg <= N59;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_53_sv2v_reg <= N58;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_52_sv2v_reg <= N57;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_51_sv2v_reg <= N56;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_50_sv2v_reg <= N55;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_49_sv2v_reg <= N54;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_48_sv2v_reg <= N53;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_47_sv2v_reg <= N52;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_46_sv2v_reg <= N51;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_45_sv2v_reg <= N50;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_44_sv2v_reg <= N49;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_43_sv2v_reg <= N48;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_42_sv2v_reg <= N47;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_41_sv2v_reg <= N46;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_40_sv2v_reg <= N45;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_39_sv2v_reg <= N44;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_38_sv2v_reg <= N43;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_37_sv2v_reg <= N42;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_36_sv2v_reg <= N41;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_35_sv2v_reg <= N40;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_34_sv2v_reg <= N39;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_33_sv2v_reg <= N38;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_32_sv2v_reg <= N37;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_31_sv2v_reg <= N36;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_30_sv2v_reg <= N35;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_29_sv2v_reg <= N34;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_28_sv2v_reg <= N33;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_27_sv2v_reg <= N32;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_26_sv2v_reg <= N31;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_25_sv2v_reg <= N30;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_24_sv2v_reg <= N29;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_23_sv2v_reg <= N28;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_22_sv2v_reg <= N27;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_21_sv2v_reg <= N26;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_20_sv2v_reg <= N25;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_19_sv2v_reg <= N24;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_18_sv2v_reg <= N23;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_17_sv2v_reg <= N22;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_16_sv2v_reg <= N21;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_15_sv2v_reg <= N20;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_14_sv2v_reg <= N19;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_13_sv2v_reg <= N18;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_12_sv2v_reg <= N17;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_11_sv2v_reg <= N16;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_10_sv2v_reg <= N15;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_9_sv2v_reg <= N14;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_8_sv2v_reg <= N13;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_7_sv2v_reg <= N12;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_6_sv2v_reg <= N11;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_5_sv2v_reg <= N10;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_4_sv2v_reg <= N9;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_3_sv2v_reg <= N8;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_2_sv2v_reg <= N7;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_1_sv2v_reg <= N6;
    end 
  end


  always @(posedge clk_i) begin
    if(el1_en_i) begin
      el1_snoop_o_0_sv2v_reg <= N5;
    end 
  end

  assign { N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 } = (N0)? el0_snoop_o : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N1)? data_i : 1'b0;
  assign N0 = mux0_sel_i;
  assign N1 = N4;
  assign data_o = (N2)? el1_snoop_o : 
                  (N3)? data_i : 1'b0;
  assign N2 = mux1_sel_i;
  assign N3 = N120;
  assign N4 = ~mux0_sel_i;
  assign N120 = ~mux1_sel_i;

endmodule