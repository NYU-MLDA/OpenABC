module rvmaskandmatch
(
  mask,
  data,
  masken,
  match
);

  input [31:0] mask;
  input [31:0] data;
  input masken;
  output match;
  wire match,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,masken_or_fullmask,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683;
  wire [31:0] matchvec;
  assign N0 = mask[0] ^ data[0];
  assign N63 = ~N0;
  assign N1 = mask[1] ^ data[1];
  assign N66 = ~N1;
  assign N2 = mask[2] ^ data[2];
  assign N69 = ~N2;
  assign N3 = mask[3] ^ data[3];
  assign N72 = ~N3;
  assign N4 = mask[4] ^ data[4];
  assign N75 = ~N4;
  assign N5 = mask[5] ^ data[5];
  assign N78 = ~N5;
  assign N6 = mask[6] ^ data[6];
  assign N81 = ~N6;
  assign N7 = mask[7] ^ data[7];
  assign N84 = ~N7;
  assign N8 = mask[8] ^ data[8];
  assign N87 = ~N8;
  assign N9 = mask[9] ^ data[9];
  assign N90 = ~N9;
  assign N10 = mask[10] ^ data[10];
  assign N93 = ~N10;
  assign N11 = mask[11] ^ data[11];
  assign N96 = ~N11;
  assign N12 = mask[12] ^ data[12];
  assign N99 = ~N12;
  assign N13 = mask[13] ^ data[13];
  assign N102 = ~N13;
  assign N14 = mask[14] ^ data[14];
  assign N105 = ~N14;
  assign N15 = mask[15] ^ data[15];
  assign N108 = ~N15;
  assign N16 = mask[16] ^ data[16];
  assign N111 = ~N16;
  assign N17 = mask[17] ^ data[17];
  assign N114 = ~N17;
  assign N18 = mask[18] ^ data[18];
  assign N117 = ~N18;
  assign N19 = mask[19] ^ data[19];
  assign N120 = ~N19;
  assign N20 = mask[20] ^ data[20];
  assign N123 = ~N20;
  assign N21 = mask[21] ^ data[21];
  assign N126 = ~N21;
  assign N22 = mask[22] ^ data[22];
  assign N129 = ~N22;
  assign N23 = mask[23] ^ data[23];
  assign N132 = ~N23;
  assign N24 = mask[24] ^ data[24];
  assign N135 = ~N24;
  assign N25 = mask[25] ^ data[25];
  assign N138 = ~N25;
  assign N26 = mask[26] ^ data[26];
  assign N141 = ~N26;
  assign N27 = mask[27] ^ data[27];
  assign N144 = ~N27;
  assign N28 = mask[28] ^ data[28];
  assign N147 = ~N28;
  assign N29 = mask[29] ^ data[29];
  assign N150 = ~N29;
  assign N30 = mask[30] ^ data[30];
  assign N153 = ~N30;
  assign N31 = mask[31] ^ data[31];
  assign N156 = ~N31;
  assign matchvec[1] = (N32)? 1'b1 :
                       (N65)? N66 : 1'b0;
  assign N32 = N64;
  assign matchvec[2] = (N33)? 1'b1 :
                       (N68)? N69 : 1'b0;
  assign N33 = N67;
  assign matchvec[3] = (N34)? 1'b1 :
                       (N71)? N72 : 1'b0;
  assign N34 = N70;
  assign matchvec[4] = (N35)? 1'b1 :
                       (N74)? N75 : 1'b0;
  assign N35 = N73;
  assign matchvec[5] = (N36)? 1'b1 :
                       (N77)? N78 : 1'b0;
  assign N36 = N76;
  assign matchvec[6] = (N37)? 1'b1 :
                       (N80)? N81 : 1'b0;
  assign N37 = N79;
  assign matchvec[7] = (N38)? 1'b1 :
                       (N83)? N84 : 1'b0;
  assign N38 = N82;
  assign matchvec[8] = (N39)? 1'b1 :
                       (N86)? N87 : 1'b0;
  assign N39 = N85;
  assign matchvec[9] = (N40)? 1'b1 :
                       (N89)? N90 : 1'b0;
  assign N40 = N88;
  assign matchvec[10] = (N41)? 1'b1 :
                        (N92)? N93 : 1'b0;
  assign N41 = N91;
  assign matchvec[11] = (N42)? 1'b1 :
                        (N95)? N96 : 1'b0;
  assign N42 = N94;
  assign matchvec[12] = (N43)? 1'b1 :
                        (N98)? N99 : 1'b0;
  assign N43 = N97;
  assign matchvec[13] = (N44)? 1'b1 :
                        (N101)? N102 : 1'b0;
  assign N44 = N100;
  assign matchvec[14] = (N45)? 1'b1 :
                        (N104)? N105 : 1'b0;
  assign N45 = N103;
  assign matchvec[15] = (N46)? 1'b1 :
                        (N107)? N108 : 1'b0;
  assign N46 = N106;
  assign matchvec[16] = (N47)? 1'b1 :
                        (N110)? N111 : 1'b0;
  assign N47 = N109;
  assign matchvec[17] = (N48)? 1'b1 :
                        (N113)? N114 : 1'b0;
  assign N48 = N112;
  assign matchvec[18] = (N49)? 1'b1 :
                        (N116)? N117 : 1'b0;
  assign N49 = N115;
  assign matchvec[19] = (N50)? 1'b1 :
                        (N119)? N120 : 1'b0;
  assign N50 = N118;
  assign matchvec[20] = (N51)? 1'b1 :
                        (N122)? N123 : 1'b0;
  assign N51 = N121;
  assign matchvec[21] = (N52)? 1'b1 :
                        (N125)? N126 : 1'b0;
  assign N52 = N124;
  assign matchvec[22] = (N53)? 1'b1 :
                        (N128)? N129 : 1'b0;
  assign N53 = N127;
  assign matchvec[23] = (N54)? 1'b1 :
                        (N131)? N132 : 1'b0;
  assign N54 = N130;
  assign matchvec[24] = (N55)? 1'b1 :
                        (N134)? N135 : 1'b0;
  assign N55 = N133;
  assign matchvec[25] = (N56)? 1'b1 :
                        (N137)? N138 : 1'b0;
  assign N56 = N136;
  assign matchvec[26] = (N57)? 1'b1 :
                        (N140)? N141 : 1'b0;
  assign N57 = N139;
  assign matchvec[27] = (N58)? 1'b1 :
                        (N143)? N144 : 1'b0;
  assign N58 = N142;
  assign matchvec[28] = (N59)? 1'b1 :
                        (N146)? N147 : 1'b0;
  assign N59 = N145;
  assign matchvec[29] = (N60)? 1'b1 :
                        (N149)? N150 : 1'b0;
  assign N60 = N148;
  assign matchvec[30] = (N61)? 1'b1 :
                        (N152)? N153 : 1'b0;
  assign N61 = N151;
  assign matchvec[31] = (N62)? 1'b1 :
                        (N155)? N156 : 1'b0;
  assign N62 = N154;
  assign masken_or_fullmask = masken & N188;
  assign N188 = ~N187;
  assign N187 = N186 & mask[0];
  assign N186 = N185 & mask[1];
  assign N185 = N184 & mask[2];
  assign N184 = N183 & mask[3];
  assign N183 = N182 & mask[4];
  assign N182 = N181 & mask[5];
  assign N181 = N180 & mask[6];
  assign N180 = N179 & mask[7];
  assign N179 = N178 & mask[8];
  assign N178 = N177 & mask[9];
  assign N177 = N176 & mask[10];
  assign N176 = N175 & mask[11];
  assign N175 = N174 & mask[12];
  assign N174 = N173 & mask[13];
  assign N173 = N172 & mask[14];
  assign N172 = N171 & mask[15];
  assign N171 = N170 & mask[16];
  assign N170 = N169 & mask[17];
  assign N169 = N168 & mask[18];
  assign N168 = N167 & mask[19];
  assign N167 = N166 & mask[20];
  assign N166 = N165 & mask[21];
  assign N165 = N164 & mask[22];
  assign N164 = N163 & mask[23];
  assign N163 = N162 & mask[24];
  assign N162 = N161 & mask[25];
  assign N161 = N160 & mask[26];
  assign N160 = N159 & mask[27];
  assign N159 = N158 & mask[28];
  assign N158 = N157 & mask[29];
  assign N157 = mask[31] & mask[30];
  assign matchvec[0] = masken_or_fullmask | N63;
  assign N64 = mask[0] & masken_or_fullmask;
  assign N65 = ~N64;
  assign N67 = N189 & masken_or_fullmask;
  assign N189 = mask[1] & mask[0];
  assign N68 = ~N67;
  assign N70 = N191 & masken_or_fullmask;
  assign N191 = N190 & mask[0];
  assign N190 = mask[2] & mask[1];
  assign N71 = ~N70;
  assign N73 = N194 & masken_or_fullmask;
  assign N194 = N193 & mask[0];
  assign N193 = N192 & mask[1];
  assign N192 = mask[3] & mask[2];
  assign N74 = ~N73;
  assign N76 = N198 & masken_or_fullmask;
  assign N198 = N197 & mask[0];
  assign N197 = N196 & mask[1];
  assign N196 = N195 & mask[2];
  assign N195 = mask[4] & mask[3];
  assign N77 = ~N76;
  assign N79 = N203 & masken_or_fullmask;
  assign N203 = N202 & mask[0];
  assign N202 = N201 & mask[1];
  assign N201 = N200 & mask[2];
  assign N200 = N199 & mask[3];
  assign N199 = mask[5] & mask[4];
  assign N80 = ~N79;
  assign N82 = N209 & masken_or_fullmask;
  assign N209 = N208 & mask[0];
  assign N208 = N207 & mask[1];
  assign N207 = N206 & mask[2];
  assign N206 = N205 & mask[3];
  assign N205 = N204 & mask[4];
  assign N204 = mask[6] & mask[5];
  assign N83 = ~N82;
  assign N85 = N216 & masken_or_fullmask;
  assign N216 = N215 & mask[0];
  assign N215 = N214 & mask[1];
  assign N214 = N213 & mask[2];
  assign N213 = N212 & mask[3];
  assign N212 = N211 & mask[4];
  assign N211 = N210 & mask[5];
  assign N210 = mask[7] & mask[6];
  assign N86 = ~N85;
  assign N88 = N224 & masken_or_fullmask;
  assign N224 = N223 & mask[0];
  assign N223 = N222 & mask[1];
  assign N222 = N221 & mask[2];
  assign N221 = N220 & mask[3];
  assign N220 = N219 & mask[4];
  assign N219 = N218 & mask[5];
  assign N218 = N217 & mask[6];
  assign N217 = mask[8] & mask[7];
  assign N89 = ~N88;
  assign N91 = N233 & masken_or_fullmask;
  assign N233 = N232 & mask[0];
  assign N232 = N231 & mask[1];
  assign N231 = N230 & mask[2];
  assign N230 = N229 & mask[3];
  assign N229 = N228 & mask[4];
  assign N228 = N227 & mask[5];
  assign N227 = N226 & mask[6];
  assign N226 = N225 & mask[7];
  assign N225 = mask[9] & mask[8];
  assign N92 = ~N91;
  assign N94 = N243 & masken_or_fullmask;
  assign N243 = N242 & mask[0];
  assign N242 = N241 & mask[1];
  assign N241 = N240 & mask[2];
  assign N240 = N239 & mask[3];
  assign N239 = N238 & mask[4];
  assign N238 = N237 & mask[5];
  assign N237 = N236 & mask[6];
  assign N236 = N235 & mask[7];
  assign N235 = N234 & mask[8];
  assign N234 = mask[10] & mask[9];
  assign N95 = ~N94;
  assign N97 = N254 & masken_or_fullmask;
  assign N254 = N253 & mask[0];
  assign N253 = N252 & mask[1];
  assign N252 = N251 & mask[2];
  assign N251 = N250 & mask[3];
  assign N250 = N249 & mask[4];
  assign N249 = N248 & mask[5];
  assign N248 = N247 & mask[6];
  assign N247 = N246 & mask[7];
  assign N246 = N245 & mask[8];
  assign N245 = N244 & mask[9];
  assign N244 = mask[11] & mask[10];
  assign N98 = ~N97;
  assign N100 = N266 & masken_or_fullmask;
  assign N266 = N265 & mask[0];
  assign N265 = N264 & mask[1];
  assign N264 = N263 & mask[2];
  assign N263 = N262 & mask[3];
  assign N262 = N261 & mask[4];
  assign N261 = N260 & mask[5];
  assign N260 = N259 & mask[6];
  assign N259 = N258 & mask[7];
  assign N258 = N257 & mask[8];
  assign N257 = N256 & mask[9];
  assign N256 = N255 & mask[10];
  assign N255 = mask[12] & mask[11];
  assign N101 = ~N100;
  assign N103 = N279 & masken_or_fullmask;
  assign N279 = N278 & mask[0];
  assign N278 = N277 & mask[1];
  assign N277 = N276 & mask[2];
  assign N276 = N275 & mask[3];
  assign N275 = N274 & mask[4];
  assign N274 = N273 & mask[5];
  assign N273 = N272 & mask[6];
  assign N272 = N271 & mask[7];
  assign N271 = N270 & mask[8];
  assign N270 = N269 & mask[9];
  assign N269 = N268 & mask[10];
  assign N268 = N267 & mask[11];
  assign N267 = mask[13] & mask[12];
  assign N104 = ~N103;
  assign N106 = N293 & masken_or_fullmask;
  assign N293 = N292 & mask[0];
  assign N292 = N291 & mask[1];
  assign N291 = N290 & mask[2];
  assign N290 = N289 & mask[3];
  assign N289 = N288 & mask[4];
  assign N288 = N287 & mask[5];
  assign N287 = N286 & mask[6];
  assign N286 = N285 & mask[7];
  assign N285 = N284 & mask[8];
  assign N284 = N283 & mask[9];
  assign N283 = N282 & mask[10];
  assign N282 = N281 & mask[11];
  assign N281 = N280 & mask[12];
  assign N280 = mask[14] & mask[13];
  assign N107 = ~N106;
  assign N109 = N308 & masken_or_fullmask;
  assign N308 = N307 & mask[0];
  assign N307 = N306 & mask[1];
  assign N306 = N305 & mask[2];
  assign N305 = N304 & mask[3];
  assign N304 = N303 & mask[4];
  assign N303 = N302 & mask[5];
  assign N302 = N301 & mask[6];
  assign N301 = N300 & mask[7];
  assign N300 = N299 & mask[8];
  assign N299 = N298 & mask[9];
  assign N298 = N297 & mask[10];
  assign N297 = N296 & mask[11];
  assign N296 = N295 & mask[12];
  assign N295 = N294 & mask[13];
  assign N294 = mask[15] & mask[14];
  assign N110 = ~N109;
  assign N112 = N324 & masken_or_fullmask;
  assign N324 = N323 & mask[0];
  assign N323 = N322 & mask[1];
  assign N322 = N321 & mask[2];
  assign N321 = N320 & mask[3];
  assign N320 = N319 & mask[4];
  assign N319 = N318 & mask[5];
  assign N318 = N317 & mask[6];
  assign N317 = N316 & mask[7];
  assign N316 = N315 & mask[8];
  assign N315 = N314 & mask[9];
  assign N314 = N313 & mask[10];
  assign N313 = N312 & mask[11];
  assign N312 = N311 & mask[12];
  assign N311 = N310 & mask[13];
  assign N310 = N309 & mask[14];
  assign N309 = mask[16] & mask[15];
  assign N113 = ~N112;
  assign N115 = N341 & masken_or_fullmask;
  assign N341 = N340 & mask[0];
  assign N340 = N339 & mask[1];
  assign N339 = N338 & mask[2];
  assign N338 = N337 & mask[3];
  assign N337 = N336 & mask[4];
  assign N336 = N335 & mask[5];
  assign N335 = N334 & mask[6];
  assign N334 = N333 & mask[7];
  assign N333 = N332 & mask[8];
  assign N332 = N331 & mask[9];
  assign N331 = N330 & mask[10];
  assign N330 = N329 & mask[11];
  assign N329 = N328 & mask[12];
  assign N328 = N327 & mask[13];
  assign N327 = N326 & mask[14];
  assign N326 = N325 & mask[15];
  assign N325 = mask[17] & mask[16];
  assign N116 = ~N115;
  assign N118 = N359 & masken_or_fullmask;
  assign N359 = N358 & mask[0];
  assign N358 = N357 & mask[1];
  assign N357 = N356 & mask[2];
  assign N356 = N355 & mask[3];
  assign N355 = N354 & mask[4];
  assign N354 = N353 & mask[5];
  assign N353 = N352 & mask[6];
  assign N352 = N351 & mask[7];
  assign N351 = N350 & mask[8];
  assign N350 = N349 & mask[9];
  assign N349 = N348 & mask[10];
  assign N348 = N347 & mask[11];
  assign N347 = N346 & mask[12];
  assign N346 = N345 & mask[13];
  assign N345 = N344 & mask[14];
  assign N344 = N343 & mask[15];
  assign N343 = N342 & mask[16];
  assign N342 = mask[18] & mask[17];
  assign N119 = ~N118;
  assign N121 = N378 & masken_or_fullmask;
  assign N378 = N377 & mask[0];
  assign N377 = N376 & mask[1];
  assign N376 = N375 & mask[2];
  assign N375 = N374 & mask[3];
  assign N374 = N373 & mask[4];
  assign N373 = N372 & mask[5];
  assign N372 = N371 & mask[6];
  assign N371 = N370 & mask[7];
  assign N370 = N369 & mask[8];
  assign N369 = N368 & mask[9];
  assign N368 = N367 & mask[10];
  assign N367 = N366 & mask[11];
  assign N366 = N365 & mask[12];
  assign N365 = N364 & mask[13];
  assign N364 = N363 & mask[14];
  assign N363 = N362 & mask[15];
  assign N362 = N361 & mask[16];
  assign N361 = N360 & mask[17];
  assign N360 = mask[19] & mask[18];
  assign N122 = ~N121;
  assign N124 = N398 & masken_or_fullmask;
  assign N398 = N397 & mask[0];
  assign N397 = N396 & mask[1];
  assign N396 = N395 & mask[2];
  assign N395 = N394 & mask[3];
  assign N394 = N393 & mask[4];
  assign N393 = N392 & mask[5];
  assign N392 = N391 & mask[6];
  assign N391 = N390 & mask[7];
  assign N390 = N389 & mask[8];
  assign N389 = N388 & mask[9];
  assign N388 = N387 & mask[10];
  assign N387 = N386 & mask[11];
  assign N386 = N385 & mask[12];
  assign N385 = N384 & mask[13];
  assign N384 = N383 & mask[14];
  assign N383 = N382 & mask[15];
  assign N382 = N381 & mask[16];
  assign N381 = N380 & mask[17];
  assign N380 = N379 & mask[18];
  assign N379 = mask[20] & mask[19];
  assign N125 = ~N124;
  assign N127 = N419 & masken_or_fullmask;
  assign N419 = N418 & mask[0];
  assign N418 = N417 & mask[1];
  assign N417 = N416 & mask[2];
  assign N416 = N415 & mask[3];
  assign N415 = N414 & mask[4];
  assign N414 = N413 & mask[5];
  assign N413 = N412 & mask[6];
  assign N412 = N411 & mask[7];
  assign N411 = N410 & mask[8];
  assign N410 = N409 & mask[9];
  assign N409 = N408 & mask[10];
  assign N408 = N407 & mask[11];
  assign N407 = N406 & mask[12];
  assign N406 = N405 & mask[13];
  assign N405 = N404 & mask[14];
  assign N404 = N403 & mask[15];
  assign N403 = N402 & mask[16];
  assign N402 = N401 & mask[17];
  assign N401 = N400 & mask[18];
  assign N400 = N399 & mask[19];
  assign N399 = mask[21] & mask[20];
  assign N128 = ~N127;
  assign N130 = N441 & masken_or_fullmask;
  assign N441 = N440 & mask[0];
  assign N440 = N439 & mask[1];
  assign N439 = N438 & mask[2];
  assign N438 = N437 & mask[3];
  assign N437 = N436 & mask[4];
  assign N436 = N435 & mask[5];
  assign N435 = N434 & mask[6];
  assign N434 = N433 & mask[7];
  assign N433 = N432 & mask[8];
  assign N432 = N431 & mask[9];
  assign N431 = N430 & mask[10];
  assign N430 = N429 & mask[11];
  assign N429 = N428 & mask[12];
  assign N428 = N427 & mask[13];
  assign N427 = N426 & mask[14];
  assign N426 = N425 & mask[15];
  assign N425 = N424 & mask[16];
  assign N424 = N423 & mask[17];
  assign N423 = N422 & mask[18];
  assign N422 = N421 & mask[19];
  assign N421 = N420 & mask[20];
  assign N420 = mask[22] & mask[21];
  assign N131 = ~N130;
  assign N133 = N464 & masken_or_fullmask;
  assign N464 = N463 & mask[0];
  assign N463 = N462 & mask[1];
  assign N462 = N461 & mask[2];
  assign N461 = N460 & mask[3];
  assign N460 = N459 & mask[4];
  assign N459 = N458 & mask[5];
  assign N458 = N457 & mask[6];
  assign N457 = N456 & mask[7];
  assign N456 = N455 & mask[8];
  assign N455 = N454 & mask[9];
  assign N454 = N453 & mask[10];
  assign N453 = N452 & mask[11];
  assign N452 = N451 & mask[12];
  assign N451 = N450 & mask[13];
  assign N450 = N449 & mask[14];
  assign N449 = N448 & mask[15];
  assign N448 = N447 & mask[16];
  assign N447 = N446 & mask[17];
  assign N446 = N445 & mask[18];
  assign N445 = N444 & mask[19];
  assign N444 = N443 & mask[20];
  assign N443 = N442 & mask[21];
  assign N442 = mask[23] & mask[22];
  assign N134 = ~N133;
  assign N136 = N488 & masken_or_fullmask;
  assign N488 = N487 & mask[0];
  assign N487 = N486 & mask[1];
  assign N486 = N485 & mask[2];
  assign N485 = N484 & mask[3];
  assign N484 = N483 & mask[4];
  assign N483 = N482 & mask[5];
  assign N482 = N481 & mask[6];
  assign N481 = N480 & mask[7];
  assign N480 = N479 & mask[8];
  assign N479 = N478 & mask[9];
  assign N478 = N477 & mask[10];
  assign N477 = N476 & mask[11];
  assign N476 = N475 & mask[12];
  assign N475 = N474 & mask[13];
  assign N474 = N473 & mask[14];
  assign N473 = N472 & mask[15];
  assign N472 = N471 & mask[16];
  assign N471 = N470 & mask[17];
  assign N470 = N469 & mask[18];
  assign N469 = N468 & mask[19];
  assign N468 = N467 & mask[20];
  assign N467 = N466 & mask[21];
  assign N466 = N465 & mask[22];
  assign N465 = mask[24] & mask[23];
  assign N137 = ~N136;
  assign N139 = N513 & masken_or_fullmask;
  assign N513 = N512 & mask[0];
  assign N512 = N511 & mask[1];
  assign N511 = N510 & mask[2];
  assign N510 = N509 & mask[3];
  assign N509 = N508 & mask[4];
  assign N508 = N507 & mask[5];
  assign N507 = N506 & mask[6];
  assign N506 = N505 & mask[7];
  assign N505 = N504 & mask[8];
  assign N504 = N503 & mask[9];
  assign N503 = N502 & mask[10];
  assign N502 = N501 & mask[11];
  assign N501 = N500 & mask[12];
  assign N500 = N499 & mask[13];
  assign N499 = N498 & mask[14];
  assign N498 = N497 & mask[15];
  assign N497 = N496 & mask[16];
  assign N496 = N495 & mask[17];
  assign N495 = N494 & mask[18];
  assign N494 = N493 & mask[19];
  assign N493 = N492 & mask[20];
  assign N492 = N491 & mask[21];
  assign N491 = N490 & mask[22];
  assign N490 = N489 & mask[23];
  assign N489 = mask[25] & mask[24];
  assign N140 = ~N139;
  assign N142 = N539 & masken_or_fullmask;
  assign N539 = N538 & mask[0];
  assign N538 = N537 & mask[1];
  assign N537 = N536 & mask[2];
  assign N536 = N535 & mask[3];
  assign N535 = N534 & mask[4];
  assign N534 = N533 & mask[5];
  assign N533 = N532 & mask[6];
  assign N532 = N531 & mask[7];
  assign N531 = N530 & mask[8];
  assign N530 = N529 & mask[9];
  assign N529 = N528 & mask[10];
  assign N528 = N527 & mask[11];
  assign N527 = N526 & mask[12];
  assign N526 = N525 & mask[13];
  assign N525 = N524 & mask[14];
  assign N524 = N523 & mask[15];
  assign N523 = N522 & mask[16];
  assign N522 = N521 & mask[17];
  assign N521 = N520 & mask[18];
  assign N520 = N519 & mask[19];
  assign N519 = N518 & mask[20];
  assign N518 = N517 & mask[21];
  assign N517 = N516 & mask[22];
  assign N516 = N515 & mask[23];
  assign N515 = N514 & mask[24];
  assign N514 = mask[26] & mask[25];
  assign N143 = ~N142;
  assign N145 = N566 & masken_or_fullmask;
  assign N566 = N565 & mask[0];
  assign N565 = N564 & mask[1];
  assign N564 = N563 & mask[2];
  assign N563 = N562 & mask[3];
  assign N562 = N561 & mask[4];
  assign N561 = N560 & mask[5];
  assign N560 = N559 & mask[6];
  assign N559 = N558 & mask[7];
  assign N558 = N557 & mask[8];
  assign N557 = N556 & mask[9];
  assign N556 = N555 & mask[10];
  assign N555 = N554 & mask[11];
  assign N554 = N553 & mask[12];
  assign N553 = N552 & mask[13];
  assign N552 = N551 & mask[14];
  assign N551 = N550 & mask[15];
  assign N550 = N549 & mask[16];
  assign N549 = N548 & mask[17];
  assign N548 = N547 & mask[18];
  assign N547 = N546 & mask[19];
  assign N546 = N545 & mask[20];
  assign N545 = N544 & mask[21];
  assign N544 = N543 & mask[22];
  assign N543 = N542 & mask[23];
  assign N542 = N541 & mask[24];
  assign N541 = N540 & mask[25];
  assign N540 = mask[27] & mask[26];
  assign N146 = ~N145;
  assign N148 = N594 & masken_or_fullmask;
  assign N594 = N593 & mask[0];
  assign N593 = N592 & mask[1];
  assign N592 = N591 & mask[2];
  assign N591 = N590 & mask[3];
  assign N590 = N589 & mask[4];
  assign N589 = N588 & mask[5];
  assign N588 = N587 & mask[6];
  assign N587 = N586 & mask[7];
  assign N586 = N585 & mask[8];
  assign N585 = N584 & mask[9];
  assign N584 = N583 & mask[10];
  assign N583 = N582 & mask[11];
  assign N582 = N581 & mask[12];
  assign N581 = N580 & mask[13];
  assign N580 = N579 & mask[14];
  assign N579 = N578 & mask[15];
  assign N578 = N577 & mask[16];
  assign N577 = N576 & mask[17];
  assign N576 = N575 & mask[18];
  assign N575 = N574 & mask[19];
  assign N574 = N573 & mask[20];
  assign N573 = N572 & mask[21];
  assign N572 = N571 & mask[22];
  assign N571 = N570 & mask[23];
  assign N570 = N569 & mask[24];
  assign N569 = N568 & mask[25];
  assign N568 = N567 & mask[26];
  assign N567 = mask[28] & mask[27];
  assign N149 = ~N148;
  assign N151 = N623 & masken_or_fullmask;
  assign N623 = N622 & mask[0];
  assign N622 = N621 & mask[1];
  assign N621 = N620 & mask[2];
  assign N620 = N619 & mask[3];
  assign N619 = N618 & mask[4];
  assign N618 = N617 & mask[5];
  assign N617 = N616 & mask[6];
  assign N616 = N615 & mask[7];
  assign N615 = N614 & mask[8];
  assign N614 = N613 & mask[9];
  assign N613 = N612 & mask[10];
  assign N612 = N611 & mask[11];
  assign N611 = N610 & mask[12];
  assign N610 = N609 & mask[13];
  assign N609 = N608 & mask[14];
  assign N608 = N607 & mask[15];
  assign N607 = N606 & mask[16];
  assign N606 = N605 & mask[17];
  assign N605 = N604 & mask[18];
  assign N604 = N603 & mask[19];
  assign N603 = N602 & mask[20];
  assign N602 = N601 & mask[21];
  assign N601 = N600 & mask[22];
  assign N600 = N599 & mask[23];
  assign N599 = N598 & mask[24];
  assign N598 = N597 & mask[25];
  assign N597 = N596 & mask[26];
  assign N596 = N595 & mask[27];
  assign N595 = mask[29] & mask[28];
  assign N152 = ~N151;
  assign N154 = N653 & masken_or_fullmask;
  assign N653 = N652 & mask[0];
  assign N652 = N651 & mask[1];
  assign N651 = N650 & mask[2];
  assign N650 = N649 & mask[3];
  assign N649 = N648 & mask[4];
  assign N648 = N647 & mask[5];
  assign N647 = N646 & mask[6];
  assign N646 = N645 & mask[7];
  assign N645 = N644 & mask[8];
  assign N644 = N643 & mask[9];
  assign N643 = N642 & mask[10];
  assign N642 = N641 & mask[11];
  assign N641 = N640 & mask[12];
  assign N640 = N639 & mask[13];
  assign N639 = N638 & mask[14];
  assign N638 = N637 & mask[15];
  assign N637 = N636 & mask[16];
  assign N636 = N635 & mask[17];
  assign N635 = N634 & mask[18];
  assign N634 = N633 & mask[19];
  assign N633 = N632 & mask[20];
  assign N632 = N631 & mask[21];
  assign N631 = N630 & mask[22];
  assign N630 = N629 & mask[23];
  assign N629 = N628 & mask[24];
  assign N628 = N627 & mask[25];
  assign N627 = N626 & mask[26];
  assign N626 = N625 & mask[27];
  assign N625 = N624 & mask[28];
  assign N624 = mask[30] & mask[29];
  assign N155 = ~N154;
  assign match = N683 & matchvec[0];
  assign N683 = N682 & matchvec[1];
  assign N682 = N681 & matchvec[2];
  assign N681 = N680 & matchvec[3];
  assign N680 = N679 & matchvec[4];
  assign N679 = N678 & matchvec[5];
  assign N678 = N677 & matchvec[6];
  assign N677 = N676 & matchvec[7];
  assign N676 = N675 & matchvec[8];
  assign N675 = N674 & matchvec[9];
  assign N674 = N673 & matchvec[10];
  assign N673 = N672 & matchvec[11];
  assign N672 = N671 & matchvec[12];
  assign N671 = N670 & matchvec[13];
  assign N670 = N669 & matchvec[14];
  assign N669 = N668 & matchvec[15];
  assign N668 = N667 & matchvec[16];
  assign N667 = N666 & matchvec[17];
  assign N666 = N665 & matchvec[18];
  assign N665 = N664 & matchvec[19];
  assign N664 = N663 & matchvec[20];
  assign N663 = N662 & matchvec[21];
  assign N662 = N661 & matchvec[22];
  assign N661 = N660 & matchvec[23];
  assign N660 = N659 & matchvec[24];
  assign N659 = N658 & matchvec[25];
  assign N658 = N657 & matchvec[26];
  assign N657 = N656 & matchvec[27];
  assign N656 = N655 & matchvec[28];
  assign N655 = N654 & matchvec[29];
  assign N654 = matchvec[31] & matchvec[30];

endmodule