module re_name
(
  clk_i,
  rst_ni,
  flush_i,
  flush_unissied_instr_i,
  issue_instr_i,
  issue_instr_valid_i,
  issue_ack_o,
  issue_instr_o,
  issue_instr_valid_o,
  issue_ack_i
);

  input [361:0] issue_instr_i;
  output [361:0] issue_instr_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input flush_unissied_instr_i;
  input issue_instr_valid_i;
  input issue_ack_i;
  output issue_ack_o;
  output issue_instr_valid_o;
  wire [361:0] issue_instr_o;
  wire issue_ack_o,issue_instr_valid_o,issue_ack_i,issue_instr_valid_i;
  assign issue_instr_o[271] = 1'b0;
  assign issue_instr_o[277] = 1'b0;
  assign issue_instr_o[283] = 1'b0;
  assign issue_ack_o = issue_ack_i;
  assign issue_instr_o[361] = issue_instr_i[361];
  assign issue_instr_o[360] = issue_instr_i[360];
  assign issue_instr_o[359] = issue_instr_i[359];
  assign issue_instr_o[358] = issue_instr_i[358];
  assign issue_instr_o[357] = issue_instr_i[357];
  assign issue_instr_o[356] = issue_instr_i[356];
  assign issue_instr_o[355] = issue_instr_i[355];
  assign issue_instr_o[354] = issue_instr_i[354];
  assign issue_instr_o[353] = issue_instr_i[353];
  assign issue_instr_o[352] = issue_instr_i[352];
  assign issue_instr_o[351] = issue_instr_i[351];
  assign issue_instr_o[350] = issue_instr_i[350];
  assign issue_instr_o[349] = issue_instr_i[349];
  assign issue_instr_o[348] = issue_instr_i[348];
  assign issue_instr_o[347] = issue_instr_i[347];
  assign issue_instr_o[346] = issue_instr_i[346];
  assign issue_instr_o[345] = issue_instr_i[345];
  assign issue_instr_o[344] = issue_instr_i[344];
  assign issue_instr_o[343] = issue_instr_i[343];
  assign issue_instr_o[342] = issue_instr_i[342];
  assign issue_instr_o[341] = issue_instr_i[341];
  assign issue_instr_o[340] = issue_instr_i[340];
  assign issue_instr_o[339] = issue_instr_i[339];
  assign issue_instr_o[338] = issue_instr_i[338];
  assign issue_instr_o[337] = issue_instr_i[337];
  assign issue_instr_o[336] = issue_instr_i[336];
  assign issue_instr_o[335] = issue_instr_i[335];
  assign issue_instr_o[334] = issue_instr_i[334];
  assign issue_instr_o[333] = issue_instr_i[333];
  assign issue_instr_o[332] = issue_instr_i[332];
  assign issue_instr_o[331] = issue_instr_i[331];
  assign issue_instr_o[330] = issue_instr_i[330];
  assign issue_instr_o[329] = issue_instr_i[329];
  assign issue_instr_o[328] = issue_instr_i[328];
  assign issue_instr_o[327] = issue_instr_i[327];
  assign issue_instr_o[326] = issue_instr_i[326];
  assign issue_instr_o[325] = issue_instr_i[325];
  assign issue_instr_o[324] = issue_instr_i[324];
  assign issue_instr_o[323] = issue_instr_i[323];
  assign issue_instr_o[322] = issue_instr_i[322];
  assign issue_instr_o[321] = issue_instr_i[321];
  assign issue_instr_o[320] = issue_instr_i[320];
  assign issue_instr_o[319] = issue_instr_i[319];
  assign issue_instr_o[318] = issue_instr_i[318];
  assign issue_instr_o[317] = issue_instr_i[317];
  assign issue_instr_o[316] = issue_instr_i[316];
  assign issue_instr_o[315] = issue_instr_i[315];
  assign issue_instr_o[314] = issue_instr_i[314];
  assign issue_instr_o[313] = issue_instr_i[313];
  assign issue_instr_o[312] = issue_instr_i[312];
  assign issue_instr_o[311] = issue_instr_i[311];
  assign issue_instr_o[310] = issue_instr_i[310];
  assign issue_instr_o[309] = issue_instr_i[309];
  assign issue_instr_o[308] = issue_instr_i[308];
  assign issue_instr_o[307] = issue_instr_i[307];
  assign issue_instr_o[306] = issue_instr_i[306];
  assign issue_instr_o[305] = issue_instr_i[305];
  assign issue_instr_o[304] = issue_instr_i[304];
  assign issue_instr_o[303] = issue_instr_i[303];
  assign issue_instr_o[302] = issue_instr_i[302];
  assign issue_instr_o[301] = issue_instr_i[301];
  assign issue_instr_o[300] = issue_instr_i[300];
  assign issue_instr_o[299] = issue_instr_i[299];
  assign issue_instr_o[298] = issue_instr_i[298];
  assign issue_instr_o[297] = issue_instr_i[297];
  assign issue_instr_o[296] = issue_instr_i[296];
  assign issue_instr_o[295] = issue_instr_i[295];
  assign issue_instr_o[294] = issue_instr_i[294];
  assign issue_instr_o[293] = issue_instr_i[293];
  assign issue_instr_o[292] = issue_instr_i[292];
  assign issue_instr_o[291] = issue_instr_i[291];
  assign issue_instr_o[290] = issue_instr_i[290];
  assign issue_instr_o[289] = issue_instr_i[289];
  assign issue_instr_o[288] = issue_instr_i[288];
  assign issue_instr_o[287] = issue_instr_i[287];
  assign issue_instr_o[286] = issue_instr_i[286];
  assign issue_instr_o[285] = issue_instr_i[285];
  assign issue_instr_o[284] = issue_instr_i[284];
  assign issue_instr_o[282] = issue_instr_i[282];
  assign issue_instr_o[281] = issue_instr_i[281];
  assign issue_instr_o[280] = issue_instr_i[280];
  assign issue_instr_o[279] = issue_instr_i[279];
  assign issue_instr_o[278] = issue_instr_i[278];
  assign issue_instr_o[276] = issue_instr_i[276];
  assign issue_instr_o[275] = issue_instr_i[275];
  assign issue_instr_o[274] = issue_instr_i[274];
  assign issue_instr_o[273] = issue_instr_i[273];
  assign issue_instr_o[272] = issue_instr_i[272];
  assign issue_instr_o[270] = issue_instr_i[270];
  assign issue_instr_o[269] = issue_instr_i[269];
  assign issue_instr_o[268] = issue_instr_i[268];
  assign issue_instr_o[267] = issue_instr_i[267];
  assign issue_instr_o[266] = issue_instr_i[266];
  assign issue_instr_o[265] = issue_instr_i[265];
  assign issue_instr_o[264] = issue_instr_i[264];
  assign issue_instr_o[263] = issue_instr_i[263];
  assign issue_instr_o[262] = issue_instr_i[262];
  assign issue_instr_o[261] = issue_instr_i[261];
  assign issue_instr_o[260] = issue_instr_i[260];
  assign issue_instr_o[259] = issue_instr_i[259];
  assign issue_instr_o[258] = issue_instr_i[258];
  assign issue_instr_o[257] = issue_instr_i[257];
  assign issue_instr_o[256] = issue_instr_i[256];
  assign issue_instr_o[255] = issue_instr_i[255];
  assign issue_instr_o[254] = issue_instr_i[254];
  assign issue_instr_o[253] = issue_instr_i[253];
  assign issue_instr_o[252] = issue_instr_i[252];
  assign issue_instr_o[251] = issue_instr_i[251];
  assign issue_instr_o[250] = issue_instr_i[250];
  assign issue_instr_o[249] = issue_instr_i[249];
  assign issue_instr_o[248] = issue_instr_i[248];
  assign issue_instr_o[247] = issue_instr_i[247];
  assign issue_instr_o[246] = issue_instr_i[246];
  assign issue_instr_o[245] = issue_instr_i[245];
  assign issue_instr_o[244] = issue_instr_i[244];
  assign issue_instr_o[243] = issue_instr_i[243];
  assign issue_instr_o[242] = issue_instr_i[242];
  assign issue_instr_o[241] = issue_instr_i[241];
  assign issue_instr_o[240] = issue_instr_i[240];
  assign issue_instr_o[239] = issue_instr_i[239];
  assign issue_instr_o[238] = issue_instr_i[238];
  assign issue_instr_o[237] = issue_instr_i[237];
  assign issue_instr_o[236] = issue_instr_i[236];
  assign issue_instr_o[235] = issue_instr_i[235];
  assign issue_instr_o[234] = issue_instr_i[234];
  assign issue_instr_o[233] = issue_instr_i[233];
  assign issue_instr_o[232] = issue_instr_i[232];
  assign issue_instr_o[231] = issue_instr_i[231];
  assign issue_instr_o[230] = issue_instr_i[230];
  assign issue_instr_o[229] = issue_instr_i[229];
  assign issue_instr_o[228] = issue_instr_i[228];
  assign issue_instr_o[227] = issue_instr_i[227];
  assign issue_instr_o[226] = issue_instr_i[226];
  assign issue_instr_o[225] = issue_instr_i[225];
  assign issue_instr_o[224] = issue_instr_i[224];
  assign issue_instr_o[223] = issue_instr_i[223];
  assign issue_instr_o[222] = issue_instr_i[222];
  assign issue_instr_o[221] = issue_instr_i[221];
  assign issue_instr_o[220] = issue_instr_i[220];
  assign issue_instr_o[219] = issue_instr_i[219];
  assign issue_instr_o[218] = issue_instr_i[218];
  assign issue_instr_o[217] = issue_instr_i[217];
  assign issue_instr_o[216] = issue_instr_i[216];
  assign issue_instr_o[215] = issue_instr_i[215];
  assign issue_instr_o[214] = issue_instr_i[214];
  assign issue_instr_o[213] = issue_instr_i[213];
  assign issue_instr_o[212] = issue_instr_i[212];
  assign issue_instr_o[211] = issue_instr_i[211];
  assign issue_instr_o[210] = issue_instr_i[210];
  assign issue_instr_o[209] = issue_instr_i[209];
  assign issue_instr_o[208] = issue_instr_i[208];
  assign issue_instr_o[207] = issue_instr_i[207];
  assign issue_instr_o[206] = issue_instr_i[206];
  assign issue_instr_o[205] = issue_instr_i[205];
  assign issue_instr_o[204] = issue_instr_i[204];
  assign issue_instr_o[203] = issue_instr_i[203];
  assign issue_instr_o[202] = issue_instr_i[202];
  assign issue_instr_o[201] = issue_instr_i[201];
  assign issue_instr_o[200] = issue_instr_i[200];
  assign issue_instr_o[199] = issue_instr_i[199];
  assign issue_instr_o[198] = issue_instr_i[198];
  assign issue_instr_o[197] = issue_instr_i[197];
  assign issue_instr_o[196] = issue_instr_i[196];
  assign issue_instr_o[195] = issue_instr_i[195];
  assign issue_instr_o[194] = issue_instr_i[194];
  assign issue_instr_o[193] = issue_instr_i[193];
  assign issue_instr_o[192] = issue_instr_i[192];
  assign issue_instr_o[191] = issue_instr_i[191];
  assign issue_instr_o[190] = issue_instr_i[190];
  assign issue_instr_o[189] = issue_instr_i[189];
  assign issue_instr_o[188] = issue_instr_i[188];
  assign issue_instr_o[187] = issue_instr_i[187];
  assign issue_instr_o[186] = issue_instr_i[186];
  assign issue_instr_o[185] = issue_instr_i[185];
  assign issue_instr_o[184] = issue_instr_i[184];
  assign issue_instr_o[183] = issue_instr_i[183];
  assign issue_instr_o[182] = issue_instr_i[182];
  assign issue_instr_o[181] = issue_instr_i[181];
  assign issue_instr_o[180] = issue_instr_i[180];
  assign issue_instr_o[179] = issue_instr_i[179];
  assign issue_instr_o[178] = issue_instr_i[178];
  assign issue_instr_o[177] = issue_instr_i[177];
  assign issue_instr_o[176] = issue_instr_i[176];
  assign issue_instr_o[175] = issue_instr_i[175];
  assign issue_instr_o[174] = issue_instr_i[174];
  assign issue_instr_o[173] = issue_instr_i[173];
  assign issue_instr_o[172] = issue_instr_i[172];
  assign issue_instr_o[171] = issue_instr_i[171];
  assign issue_instr_o[170] = issue_instr_i[170];
  assign issue_instr_o[169] = issue_instr_i[169];
  assign issue_instr_o[168] = issue_instr_i[168];
  assign issue_instr_o[167] = issue_instr_i[167];
  assign issue_instr_o[166] = issue_instr_i[166];
  assign issue_instr_o[165] = issue_instr_i[165];
  assign issue_instr_o[164] = issue_instr_i[164];
  assign issue_instr_o[163] = issue_instr_i[163];
  assign issue_instr_o[162] = issue_instr_i[162];
  assign issue_instr_o[161] = issue_instr_i[161];
  assign issue_instr_o[160] = issue_instr_i[160];
  assign issue_instr_o[159] = issue_instr_i[159];
  assign issue_instr_o[158] = issue_instr_i[158];
  assign issue_instr_o[157] = issue_instr_i[157];
  assign issue_instr_o[156] = issue_instr_i[156];
  assign issue_instr_o[155] = issue_instr_i[155];
  assign issue_instr_o[154] = issue_instr_i[154];
  assign issue_instr_o[153] = issue_instr_i[153];
  assign issue_instr_o[152] = issue_instr_i[152];
  assign issue_instr_o[151] = issue_instr_i[151];
  assign issue_instr_o[150] = issue_instr_i[150];
  assign issue_instr_o[149] = issue_instr_i[149];
  assign issue_instr_o[148] = issue_instr_i[148];
  assign issue_instr_o[147] = issue_instr_i[147];
  assign issue_instr_o[146] = issue_instr_i[146];
  assign issue_instr_o[145] = issue_instr_i[145];
  assign issue_instr_o[144] = issue_instr_i[144];
  assign issue_instr_o[143] = issue_instr_i[143];
  assign issue_instr_o[142] = issue_instr_i[142];
  assign issue_instr_o[141] = issue_instr_i[141];
  assign issue_instr_o[140] = issue_instr_i[140];
  assign issue_instr_o[139] = issue_instr_i[139];
  assign issue_instr_o[138] = issue_instr_i[138];
  assign issue_instr_o[137] = issue_instr_i[137];
  assign issue_instr_o[136] = issue_instr_i[136];
  assign issue_instr_o[135] = issue_instr_i[135];
  assign issue_instr_o[134] = issue_instr_i[134];
  assign issue_instr_o[133] = issue_instr_i[133];
  assign issue_instr_o[132] = issue_instr_i[132];
  assign issue_instr_o[131] = issue_instr_i[131];
  assign issue_instr_o[130] = issue_instr_i[130];
  assign issue_instr_o[129] = issue_instr_i[129];
  assign issue_instr_o[128] = issue_instr_i[128];
  assign issue_instr_o[127] = issue_instr_i[127];
  assign issue_instr_o[126] = issue_instr_i[126];
  assign issue_instr_o[125] = issue_instr_i[125];
  assign issue_instr_o[124] = issue_instr_i[124];
  assign issue_instr_o[123] = issue_instr_i[123];
  assign issue_instr_o[122] = issue_instr_i[122];
  assign issue_instr_o[121] = issue_instr_i[121];
  assign issue_instr_o[120] = issue_instr_i[120];
  assign issue_instr_o[119] = issue_instr_i[119];
  assign issue_instr_o[118] = issue_instr_i[118];
  assign issue_instr_o[117] = issue_instr_i[117];
  assign issue_instr_o[116] = issue_instr_i[116];
  assign issue_instr_o[115] = issue_instr_i[115];
  assign issue_instr_o[114] = issue_instr_i[114];
  assign issue_instr_o[113] = issue_instr_i[113];
  assign issue_instr_o[112] = issue_instr_i[112];
  assign issue_instr_o[111] = issue_instr_i[111];
  assign issue_instr_o[110] = issue_instr_i[110];
  assign issue_instr_o[109] = issue_instr_i[109];
  assign issue_instr_o[108] = issue_instr_i[108];
  assign issue_instr_o[107] = issue_instr_i[107];
  assign issue_instr_o[106] = issue_instr_i[106];
  assign issue_instr_o[105] = issue_instr_i[105];
  assign issue_instr_o[104] = issue_instr_i[104];
  assign issue_instr_o[103] = issue_instr_i[103];
  assign issue_instr_o[102] = issue_instr_i[102];
  assign issue_instr_o[101] = issue_instr_i[101];
  assign issue_instr_o[100] = issue_instr_i[100];
  assign issue_instr_o[99] = issue_instr_i[99];
  assign issue_instr_o[98] = issue_instr_i[98];
  assign issue_instr_o[97] = issue_instr_i[97];
  assign issue_instr_o[96] = issue_instr_i[96];
  assign issue_instr_o[95] = issue_instr_i[95];
  assign issue_instr_o[94] = issue_instr_i[94];
  assign issue_instr_o[93] = issue_instr_i[93];
  assign issue_instr_o[92] = issue_instr_i[92];
  assign issue_instr_o[91] = issue_instr_i[91];
  assign issue_instr_o[90] = issue_instr_i[90];
  assign issue_instr_o[89] = issue_instr_i[89];
  assign issue_instr_o[88] = issue_instr_i[88];
  assign issue_instr_o[87] = issue_instr_i[87];
  assign issue_instr_o[86] = issue_instr_i[86];
  assign issue_instr_o[85] = issue_instr_i[85];
  assign issue_instr_o[84] = issue_instr_i[84];
  assign issue_instr_o[83] = issue_instr_i[83];
  assign issue_instr_o[82] = issue_instr_i[82];
  assign issue_instr_o[81] = issue_instr_i[81];
  assign issue_instr_o[80] = issue_instr_i[80];
  assign issue_instr_o[79] = issue_instr_i[79];
  assign issue_instr_o[78] = issue_instr_i[78];
  assign issue_instr_o[77] = issue_instr_i[77];
  assign issue_instr_o[76] = issue_instr_i[76];
  assign issue_instr_o[75] = issue_instr_i[75];
  assign issue_instr_o[74] = issue_instr_i[74];
  assign issue_instr_o[73] = issue_instr_i[73];
  assign issue_instr_o[72] = issue_instr_i[72];
  assign issue_instr_o[71] = issue_instr_i[71];
  assign issue_instr_o[70] = issue_instr_i[70];
  assign issue_instr_o[69] = issue_instr_i[69];
  assign issue_instr_o[68] = issue_instr_i[68];
  assign issue_instr_o[67] = issue_instr_i[67];
  assign issue_instr_o[66] = issue_instr_i[66];
  assign issue_instr_o[65] = issue_instr_i[65];
  assign issue_instr_o[64] = issue_instr_i[64];
  assign issue_instr_o[63] = issue_instr_i[63];
  assign issue_instr_o[62] = issue_instr_i[62];
  assign issue_instr_o[61] = issue_instr_i[61];
  assign issue_instr_o[60] = issue_instr_i[60];
  assign issue_instr_o[59] = issue_instr_i[59];
  assign issue_instr_o[58] = issue_instr_i[58];
  assign issue_instr_o[57] = issue_instr_i[57];
  assign issue_instr_o[56] = issue_instr_i[56];
  assign issue_instr_o[55] = issue_instr_i[55];
  assign issue_instr_o[54] = issue_instr_i[54];
  assign issue_instr_o[53] = issue_instr_i[53];
  assign issue_instr_o[52] = issue_instr_i[52];
  assign issue_instr_o[51] = issue_instr_i[51];
  assign issue_instr_o[50] = issue_instr_i[50];
  assign issue_instr_o[49] = issue_instr_i[49];
  assign issue_instr_o[48] = issue_instr_i[48];
  assign issue_instr_o[47] = issue_instr_i[47];
  assign issue_instr_o[46] = issue_instr_i[46];
  assign issue_instr_o[45] = issue_instr_i[45];
  assign issue_instr_o[44] = issue_instr_i[44];
  assign issue_instr_o[43] = issue_instr_i[43];
  assign issue_instr_o[42] = issue_instr_i[42];
  assign issue_instr_o[41] = issue_instr_i[41];
  assign issue_instr_o[40] = issue_instr_i[40];
  assign issue_instr_o[39] = issue_instr_i[39];
  assign issue_instr_o[38] = issue_instr_i[38];
  assign issue_instr_o[37] = issue_instr_i[37];
  assign issue_instr_o[36] = issue_instr_i[36];
  assign issue_instr_o[35] = issue_instr_i[35];
  assign issue_instr_o[34] = issue_instr_i[34];
  assign issue_instr_o[33] = issue_instr_i[33];
  assign issue_instr_o[32] = issue_instr_i[32];
  assign issue_instr_o[31] = issue_instr_i[31];
  assign issue_instr_o[30] = issue_instr_i[30];
  assign issue_instr_o[29] = issue_instr_i[29];
  assign issue_instr_o[28] = issue_instr_i[28];
  assign issue_instr_o[27] = issue_instr_i[27];
  assign issue_instr_o[26] = issue_instr_i[26];
  assign issue_instr_o[25] = issue_instr_i[25];
  assign issue_instr_o[24] = issue_instr_i[24];
  assign issue_instr_o[23] = issue_instr_i[23];
  assign issue_instr_o[22] = issue_instr_i[22];
  assign issue_instr_o[21] = issue_instr_i[21];
  assign issue_instr_o[20] = issue_instr_i[20];
  assign issue_instr_o[19] = issue_instr_i[19];
  assign issue_instr_o[18] = issue_instr_i[18];
  assign issue_instr_o[17] = issue_instr_i[17];
  assign issue_instr_o[16] = issue_instr_i[16];
  assign issue_instr_o[15] = issue_instr_i[15];
  assign issue_instr_o[14] = issue_instr_i[14];
  assign issue_instr_o[13] = issue_instr_i[13];
  assign issue_instr_o[12] = issue_instr_i[12];
  assign issue_instr_o[11] = issue_instr_i[11];
  assign issue_instr_o[10] = issue_instr_i[10];
  assign issue_instr_o[9] = issue_instr_i[9];
  assign issue_instr_o[8] = issue_instr_i[8];
  assign issue_instr_o[7] = issue_instr_i[7];
  assign issue_instr_o[6] = issue_instr_i[6];
  assign issue_instr_o[5] = issue_instr_i[5];
  assign issue_instr_o[4] = issue_instr_i[4];
  assign issue_instr_o[3] = issue_instr_i[3];
  assign issue_instr_o[2] = issue_instr_i[2];
  assign issue_instr_o[1] = issue_instr_i[1];
  assign issue_instr_o[0] = issue_instr_i[0];
  assign issue_instr_valid_o = issue_instr_valid_i;

endmodule