module bp_be_dcache_lce_cmd_num_cce_p1_num_lce_p2_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_data_width_p64
(
  clk_i,
  reset_i,
  lce_id_i,
  lce_sync_done_o,
  tag_set_o,
  tag_set_wakeup_o,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_yumi_o,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_data_i,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_v_o,
  tag_mem_pkt_o,
  tag_mem_pkt_yumi_i,
  stat_mem_pkt_v_o,
  stat_mem_pkt_o,
  dirty_i,
  stat_mem_pkt_yumi_i
);

  input [0:0] lce_id_i;
  input [35:0] lce_cmd_i;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  output [538:0] lce_tr_resp_o;
  output [521:0] data_mem_pkt_o;
  input [511:0] data_mem_data_i;
  output [22:0] tag_mem_pkt_o;
  output [10:0] stat_mem_pkt_o;
  input [7:0] dirty_i;
  input clk_i;
  input reset_i;
  input lce_cmd_v_i;
  input lce_resp_yumi_i;
  input lce_data_resp_ready_i;
  input lce_tr_resp_ready_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input stat_mem_pkt_yumi_i;
  output lce_sync_done_o;
  output tag_set_o;
  output tag_set_wakeup_o;
  output lce_cmd_yumi_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_tr_resp_v_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output stat_mem_pkt_v_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o;
  wire [521:0] data_mem_pkt_o;
  wire [22:0] tag_mem_pkt_o;
  wire [10:0] stat_mem_pkt_o;
  wire lce_sync_done_o,tag_set_o,tag_set_wakeup_o,lce_cmd_yumi_o,lce_resp_v_o,
  lce_data_resp_v_o,lce_tr_resp_v_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,stat_mem_pkt_v_o,N0,
  N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,lce_tr_resp_done,lce_data_resp_done,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,
  N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,
  N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1606,
  N1607;
  wire [2:0] state_n;
  reg [511:0] data_buf_r;
  reg [2:0] state_r;
  reg [0:0] sync_ack_count_r;
  reg tr_data_buffered_r,wb_data_buffered_r,wb_data_read_r,wb_dirty_cleared_r,
  invalidated_tag_r;
  assign data_mem_pkt_o[0] = 1'b0;
  assign data_mem_pkt_o[1] = 1'b0;
  assign data_mem_pkt_o[2] = 1'b0;
  assign data_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[4] = 1'b0;
  assign data_mem_pkt_o[5] = 1'b0;
  assign data_mem_pkt_o[6] = 1'b0;
  assign data_mem_pkt_o[7] = 1'b0;
  assign data_mem_pkt_o[8] = 1'b0;
  assign data_mem_pkt_o[9] = 1'b0;
  assign data_mem_pkt_o[10] = 1'b0;
  assign data_mem_pkt_o[11] = 1'b0;
  assign data_mem_pkt_o[12] = 1'b0;
  assign data_mem_pkt_o[13] = 1'b0;
  assign data_mem_pkt_o[14] = 1'b0;
  assign data_mem_pkt_o[15] = 1'b0;
  assign data_mem_pkt_o[16] = 1'b0;
  assign data_mem_pkt_o[17] = 1'b0;
  assign data_mem_pkt_o[18] = 1'b0;
  assign data_mem_pkt_o[19] = 1'b0;
  assign data_mem_pkt_o[20] = 1'b0;
  assign data_mem_pkt_o[21] = 1'b0;
  assign data_mem_pkt_o[22] = 1'b0;
  assign data_mem_pkt_o[23] = 1'b0;
  assign data_mem_pkt_o[24] = 1'b0;
  assign data_mem_pkt_o[25] = 1'b0;
  assign data_mem_pkt_o[26] = 1'b0;
  assign data_mem_pkt_o[27] = 1'b0;
  assign data_mem_pkt_o[28] = 1'b0;
  assign data_mem_pkt_o[29] = 1'b0;
  assign data_mem_pkt_o[30] = 1'b0;
  assign data_mem_pkt_o[31] = 1'b0;
  assign data_mem_pkt_o[32] = 1'b0;
  assign data_mem_pkt_o[33] = 1'b0;
  assign data_mem_pkt_o[34] = 1'b0;
  assign data_mem_pkt_o[35] = 1'b0;
  assign data_mem_pkt_o[36] = 1'b0;
  assign data_mem_pkt_o[37] = 1'b0;
  assign data_mem_pkt_o[38] = 1'b0;
  assign data_mem_pkt_o[39] = 1'b0;
  assign data_mem_pkt_o[40] = 1'b0;
  assign data_mem_pkt_o[41] = 1'b0;
  assign data_mem_pkt_o[42] = 1'b0;
  assign data_mem_pkt_o[43] = 1'b0;
  assign data_mem_pkt_o[44] = 1'b0;
  assign data_mem_pkt_o[45] = 1'b0;
  assign data_mem_pkt_o[46] = 1'b0;
  assign data_mem_pkt_o[47] = 1'b0;
  assign data_mem_pkt_o[48] = 1'b0;
  assign data_mem_pkt_o[49] = 1'b0;
  assign data_mem_pkt_o[50] = 1'b0;
  assign data_mem_pkt_o[51] = 1'b0;
  assign data_mem_pkt_o[52] = 1'b0;
  assign data_mem_pkt_o[53] = 1'b0;
  assign data_mem_pkt_o[54] = 1'b0;
  assign data_mem_pkt_o[55] = 1'b0;
  assign data_mem_pkt_o[56] = 1'b0;
  assign data_mem_pkt_o[57] = 1'b0;
  assign data_mem_pkt_o[58] = 1'b0;
  assign data_mem_pkt_o[59] = 1'b0;
  assign data_mem_pkt_o[60] = 1'b0;
  assign data_mem_pkt_o[61] = 1'b0;
  assign data_mem_pkt_o[62] = 1'b0;
  assign data_mem_pkt_o[63] = 1'b0;
  assign data_mem_pkt_o[64] = 1'b0;
  assign data_mem_pkt_o[65] = 1'b0;
  assign data_mem_pkt_o[66] = 1'b0;
  assign data_mem_pkt_o[67] = 1'b0;
  assign data_mem_pkt_o[68] = 1'b0;
  assign data_mem_pkt_o[69] = 1'b0;
  assign data_mem_pkt_o[70] = 1'b0;
  assign data_mem_pkt_o[71] = 1'b0;
  assign data_mem_pkt_o[72] = 1'b0;
  assign data_mem_pkt_o[73] = 1'b0;
  assign data_mem_pkt_o[74] = 1'b0;
  assign data_mem_pkt_o[75] = 1'b0;
  assign data_mem_pkt_o[76] = 1'b0;
  assign data_mem_pkt_o[77] = 1'b0;
  assign data_mem_pkt_o[78] = 1'b0;
  assign data_mem_pkt_o[79] = 1'b0;
  assign data_mem_pkt_o[80] = 1'b0;
  assign data_mem_pkt_o[81] = 1'b0;
  assign data_mem_pkt_o[82] = 1'b0;
  assign data_mem_pkt_o[83] = 1'b0;
  assign data_mem_pkt_o[84] = 1'b0;
  assign data_mem_pkt_o[85] = 1'b0;
  assign data_mem_pkt_o[86] = 1'b0;
  assign data_mem_pkt_o[87] = 1'b0;
  assign data_mem_pkt_o[88] = 1'b0;
  assign data_mem_pkt_o[89] = 1'b0;
  assign data_mem_pkt_o[90] = 1'b0;
  assign data_mem_pkt_o[91] = 1'b0;
  assign data_mem_pkt_o[92] = 1'b0;
  assign data_mem_pkt_o[93] = 1'b0;
  assign data_mem_pkt_o[94] = 1'b0;
  assign data_mem_pkt_o[95] = 1'b0;
  assign data_mem_pkt_o[96] = 1'b0;
  assign data_mem_pkt_o[97] = 1'b0;
  assign data_mem_pkt_o[98] = 1'b0;
  assign data_mem_pkt_o[99] = 1'b0;
  assign data_mem_pkt_o[100] = 1'b0;
  assign data_mem_pkt_o[101] = 1'b0;
  assign data_mem_pkt_o[102] = 1'b0;
  assign data_mem_pkt_o[103] = 1'b0;
  assign data_mem_pkt_o[104] = 1'b0;
  assign data_mem_pkt_o[105] = 1'b0;
  assign data_mem_pkt_o[106] = 1'b0;
  assign data_mem_pkt_o[107] = 1'b0;
  assign data_mem_pkt_o[108] = 1'b0;
  assign data_mem_pkt_o[109] = 1'b0;
  assign data_mem_pkt_o[110] = 1'b0;
  assign data_mem_pkt_o[111] = 1'b0;
  assign data_mem_pkt_o[112] = 1'b0;
  assign data_mem_pkt_o[113] = 1'b0;
  assign data_mem_pkt_o[114] = 1'b0;
  assign data_mem_pkt_o[115] = 1'b0;
  assign data_mem_pkt_o[116] = 1'b0;
  assign data_mem_pkt_o[117] = 1'b0;
  assign data_mem_pkt_o[118] = 1'b0;
  assign data_mem_pkt_o[119] = 1'b0;
  assign data_mem_pkt_o[120] = 1'b0;
  assign data_mem_pkt_o[121] = 1'b0;
  assign data_mem_pkt_o[122] = 1'b0;
  assign data_mem_pkt_o[123] = 1'b0;
  assign data_mem_pkt_o[124] = 1'b0;
  assign data_mem_pkt_o[125] = 1'b0;
  assign data_mem_pkt_o[126] = 1'b0;
  assign data_mem_pkt_o[127] = 1'b0;
  assign data_mem_pkt_o[128] = 1'b0;
  assign data_mem_pkt_o[129] = 1'b0;
  assign data_mem_pkt_o[130] = 1'b0;
  assign data_mem_pkt_o[131] = 1'b0;
  assign data_mem_pkt_o[132] = 1'b0;
  assign data_mem_pkt_o[133] = 1'b0;
  assign data_mem_pkt_o[134] = 1'b0;
  assign data_mem_pkt_o[135] = 1'b0;
  assign data_mem_pkt_o[136] = 1'b0;
  assign data_mem_pkt_o[137] = 1'b0;
  assign data_mem_pkt_o[138] = 1'b0;
  assign data_mem_pkt_o[139] = 1'b0;
  assign data_mem_pkt_o[140] = 1'b0;
  assign data_mem_pkt_o[141] = 1'b0;
  assign data_mem_pkt_o[142] = 1'b0;
  assign data_mem_pkt_o[143] = 1'b0;
  assign data_mem_pkt_o[144] = 1'b0;
  assign data_mem_pkt_o[145] = 1'b0;
  assign data_mem_pkt_o[146] = 1'b0;
  assign data_mem_pkt_o[147] = 1'b0;
  assign data_mem_pkt_o[148] = 1'b0;
  assign data_mem_pkt_o[149] = 1'b0;
  assign data_mem_pkt_o[150] = 1'b0;
  assign data_mem_pkt_o[151] = 1'b0;
  assign data_mem_pkt_o[152] = 1'b0;
  assign data_mem_pkt_o[153] = 1'b0;
  assign data_mem_pkt_o[154] = 1'b0;
  assign data_mem_pkt_o[155] = 1'b0;
  assign data_mem_pkt_o[156] = 1'b0;
  assign data_mem_pkt_o[157] = 1'b0;
  assign data_mem_pkt_o[158] = 1'b0;
  assign data_mem_pkt_o[159] = 1'b0;
  assign data_mem_pkt_o[160] = 1'b0;
  assign data_mem_pkt_o[161] = 1'b0;
  assign data_mem_pkt_o[162] = 1'b0;
  assign data_mem_pkt_o[163] = 1'b0;
  assign data_mem_pkt_o[164] = 1'b0;
  assign data_mem_pkt_o[165] = 1'b0;
  assign data_mem_pkt_o[166] = 1'b0;
  assign data_mem_pkt_o[167] = 1'b0;
  assign data_mem_pkt_o[168] = 1'b0;
  assign data_mem_pkt_o[169] = 1'b0;
  assign data_mem_pkt_o[170] = 1'b0;
  assign data_mem_pkt_o[171] = 1'b0;
  assign data_mem_pkt_o[172] = 1'b0;
  assign data_mem_pkt_o[173] = 1'b0;
  assign data_mem_pkt_o[174] = 1'b0;
  assign data_mem_pkt_o[175] = 1'b0;
  assign data_mem_pkt_o[176] = 1'b0;
  assign data_mem_pkt_o[177] = 1'b0;
  assign data_mem_pkt_o[178] = 1'b0;
  assign data_mem_pkt_o[179] = 1'b0;
  assign data_mem_pkt_o[180] = 1'b0;
  assign data_mem_pkt_o[181] = 1'b0;
  assign data_mem_pkt_o[182] = 1'b0;
  assign data_mem_pkt_o[183] = 1'b0;
  assign data_mem_pkt_o[184] = 1'b0;
  assign data_mem_pkt_o[185] = 1'b0;
  assign data_mem_pkt_o[186] = 1'b0;
  assign data_mem_pkt_o[187] = 1'b0;
  assign data_mem_pkt_o[188] = 1'b0;
  assign data_mem_pkt_o[189] = 1'b0;
  assign data_mem_pkt_o[190] = 1'b0;
  assign data_mem_pkt_o[191] = 1'b0;
  assign data_mem_pkt_o[192] = 1'b0;
  assign data_mem_pkt_o[193] = 1'b0;
  assign data_mem_pkt_o[194] = 1'b0;
  assign data_mem_pkt_o[195] = 1'b0;
  assign data_mem_pkt_o[196] = 1'b0;
  assign data_mem_pkt_o[197] = 1'b0;
  assign data_mem_pkt_o[198] = 1'b0;
  assign data_mem_pkt_o[199] = 1'b0;
  assign data_mem_pkt_o[200] = 1'b0;
  assign data_mem_pkt_o[201] = 1'b0;
  assign data_mem_pkt_o[202] = 1'b0;
  assign data_mem_pkt_o[203] = 1'b0;
  assign data_mem_pkt_o[204] = 1'b0;
  assign data_mem_pkt_o[205] = 1'b0;
  assign data_mem_pkt_o[206] = 1'b0;
  assign data_mem_pkt_o[207] = 1'b0;
  assign data_mem_pkt_o[208] = 1'b0;
  assign data_mem_pkt_o[209] = 1'b0;
  assign data_mem_pkt_o[210] = 1'b0;
  assign data_mem_pkt_o[211] = 1'b0;
  assign data_mem_pkt_o[212] = 1'b0;
  assign data_mem_pkt_o[213] = 1'b0;
  assign data_mem_pkt_o[214] = 1'b0;
  assign data_mem_pkt_o[215] = 1'b0;
  assign data_mem_pkt_o[216] = 1'b0;
  assign data_mem_pkt_o[217] = 1'b0;
  assign data_mem_pkt_o[218] = 1'b0;
  assign data_mem_pkt_o[219] = 1'b0;
  assign data_mem_pkt_o[220] = 1'b0;
  assign data_mem_pkt_o[221] = 1'b0;
  assign data_mem_pkt_o[222] = 1'b0;
  assign data_mem_pkt_o[223] = 1'b0;
  assign data_mem_pkt_o[224] = 1'b0;
  assign data_mem_pkt_o[225] = 1'b0;
  assign data_mem_pkt_o[226] = 1'b0;
  assign data_mem_pkt_o[227] = 1'b0;
  assign data_mem_pkt_o[228] = 1'b0;
  assign data_mem_pkt_o[229] = 1'b0;
  assign data_mem_pkt_o[230] = 1'b0;
  assign data_mem_pkt_o[231] = 1'b0;
  assign data_mem_pkt_o[232] = 1'b0;
  assign data_mem_pkt_o[233] = 1'b0;
  assign data_mem_pkt_o[234] = 1'b0;
  assign data_mem_pkt_o[235] = 1'b0;
  assign data_mem_pkt_o[236] = 1'b0;
  assign data_mem_pkt_o[237] = 1'b0;
  assign data_mem_pkt_o[238] = 1'b0;
  assign data_mem_pkt_o[239] = 1'b0;
  assign data_mem_pkt_o[240] = 1'b0;
  assign data_mem_pkt_o[241] = 1'b0;
  assign data_mem_pkt_o[242] = 1'b0;
  assign data_mem_pkt_o[243] = 1'b0;
  assign data_mem_pkt_o[244] = 1'b0;
  assign data_mem_pkt_o[245] = 1'b0;
  assign data_mem_pkt_o[246] = 1'b0;
  assign data_mem_pkt_o[247] = 1'b0;
  assign data_mem_pkt_o[248] = 1'b0;
  assign data_mem_pkt_o[249] = 1'b0;
  assign data_mem_pkt_o[250] = 1'b0;
  assign data_mem_pkt_o[251] = 1'b0;
  assign data_mem_pkt_o[252] = 1'b0;
  assign data_mem_pkt_o[253] = 1'b0;
  assign data_mem_pkt_o[254] = 1'b0;
  assign data_mem_pkt_o[255] = 1'b0;
  assign data_mem_pkt_o[256] = 1'b0;
  assign data_mem_pkt_o[257] = 1'b0;
  assign data_mem_pkt_o[258] = 1'b0;
  assign data_mem_pkt_o[259] = 1'b0;
  assign data_mem_pkt_o[260] = 1'b0;
  assign data_mem_pkt_o[261] = 1'b0;
  assign data_mem_pkt_o[262] = 1'b0;
  assign data_mem_pkt_o[263] = 1'b0;
  assign data_mem_pkt_o[264] = 1'b0;
  assign data_mem_pkt_o[265] = 1'b0;
  assign data_mem_pkt_o[266] = 1'b0;
  assign data_mem_pkt_o[267] = 1'b0;
  assign data_mem_pkt_o[268] = 1'b0;
  assign data_mem_pkt_o[269] = 1'b0;
  assign data_mem_pkt_o[270] = 1'b0;
  assign data_mem_pkt_o[271] = 1'b0;
  assign data_mem_pkt_o[272] = 1'b0;
  assign data_mem_pkt_o[273] = 1'b0;
  assign data_mem_pkt_o[274] = 1'b0;
  assign data_mem_pkt_o[275] = 1'b0;
  assign data_mem_pkt_o[276] = 1'b0;
  assign data_mem_pkt_o[277] = 1'b0;
  assign data_mem_pkt_o[278] = 1'b0;
  assign data_mem_pkt_o[279] = 1'b0;
  assign data_mem_pkt_o[280] = 1'b0;
  assign data_mem_pkt_o[281] = 1'b0;
  assign data_mem_pkt_o[282] = 1'b0;
  assign data_mem_pkt_o[283] = 1'b0;
  assign data_mem_pkt_o[284] = 1'b0;
  assign data_mem_pkt_o[285] = 1'b0;
  assign data_mem_pkt_o[286] = 1'b0;
  assign data_mem_pkt_o[287] = 1'b0;
  assign data_mem_pkt_o[288] = 1'b0;
  assign data_mem_pkt_o[289] = 1'b0;
  assign data_mem_pkt_o[290] = 1'b0;
  assign data_mem_pkt_o[291] = 1'b0;
  assign data_mem_pkt_o[292] = 1'b0;
  assign data_mem_pkt_o[293] = 1'b0;
  assign data_mem_pkt_o[294] = 1'b0;
  assign data_mem_pkt_o[295] = 1'b0;
  assign data_mem_pkt_o[296] = 1'b0;
  assign data_mem_pkt_o[297] = 1'b0;
  assign data_mem_pkt_o[298] = 1'b0;
  assign data_mem_pkt_o[299] = 1'b0;
  assign data_mem_pkt_o[300] = 1'b0;
  assign data_mem_pkt_o[301] = 1'b0;
  assign data_mem_pkt_o[302] = 1'b0;
  assign data_mem_pkt_o[303] = 1'b0;
  assign data_mem_pkt_o[304] = 1'b0;
  assign data_mem_pkt_o[305] = 1'b0;
  assign data_mem_pkt_o[306] = 1'b0;
  assign data_mem_pkt_o[307] = 1'b0;
  assign data_mem_pkt_o[308] = 1'b0;
  assign data_mem_pkt_o[309] = 1'b0;
  assign data_mem_pkt_o[310] = 1'b0;
  assign data_mem_pkt_o[311] = 1'b0;
  assign data_mem_pkt_o[312] = 1'b0;
  assign data_mem_pkt_o[313] = 1'b0;
  assign data_mem_pkt_o[314] = 1'b0;
  assign data_mem_pkt_o[315] = 1'b0;
  assign data_mem_pkt_o[316] = 1'b0;
  assign data_mem_pkt_o[317] = 1'b0;
  assign data_mem_pkt_o[318] = 1'b0;
  assign data_mem_pkt_o[319] = 1'b0;
  assign data_mem_pkt_o[320] = 1'b0;
  assign data_mem_pkt_o[321] = 1'b0;
  assign data_mem_pkt_o[322] = 1'b0;
  assign data_mem_pkt_o[323] = 1'b0;
  assign data_mem_pkt_o[324] = 1'b0;
  assign data_mem_pkt_o[325] = 1'b0;
  assign data_mem_pkt_o[326] = 1'b0;
  assign data_mem_pkt_o[327] = 1'b0;
  assign data_mem_pkt_o[328] = 1'b0;
  assign data_mem_pkt_o[329] = 1'b0;
  assign data_mem_pkt_o[330] = 1'b0;
  assign data_mem_pkt_o[331] = 1'b0;
  assign data_mem_pkt_o[332] = 1'b0;
  assign data_mem_pkt_o[333] = 1'b0;
  assign data_mem_pkt_o[334] = 1'b0;
  assign data_mem_pkt_o[335] = 1'b0;
  assign data_mem_pkt_o[336] = 1'b0;
  assign data_mem_pkt_o[337] = 1'b0;
  assign data_mem_pkt_o[338] = 1'b0;
  assign data_mem_pkt_o[339] = 1'b0;
  assign data_mem_pkt_o[340] = 1'b0;
  assign data_mem_pkt_o[341] = 1'b0;
  assign data_mem_pkt_o[342] = 1'b0;
  assign data_mem_pkt_o[343] = 1'b0;
  assign data_mem_pkt_o[344] = 1'b0;
  assign data_mem_pkt_o[345] = 1'b0;
  assign data_mem_pkt_o[346] = 1'b0;
  assign data_mem_pkt_o[347] = 1'b0;
  assign data_mem_pkt_o[348] = 1'b0;
  assign data_mem_pkt_o[349] = 1'b0;
  assign data_mem_pkt_o[350] = 1'b0;
  assign data_mem_pkt_o[351] = 1'b0;
  assign data_mem_pkt_o[352] = 1'b0;
  assign data_mem_pkt_o[353] = 1'b0;
  assign data_mem_pkt_o[354] = 1'b0;
  assign data_mem_pkt_o[355] = 1'b0;
  assign data_mem_pkt_o[356] = 1'b0;
  assign data_mem_pkt_o[357] = 1'b0;
  assign data_mem_pkt_o[358] = 1'b0;
  assign data_mem_pkt_o[359] = 1'b0;
  assign data_mem_pkt_o[360] = 1'b0;
  assign data_mem_pkt_o[361] = 1'b0;
  assign data_mem_pkt_o[362] = 1'b0;
  assign data_mem_pkt_o[363] = 1'b0;
  assign data_mem_pkt_o[364] = 1'b0;
  assign data_mem_pkt_o[365] = 1'b0;
  assign data_mem_pkt_o[366] = 1'b0;
  assign data_mem_pkt_o[367] = 1'b0;
  assign data_mem_pkt_o[368] = 1'b0;
  assign data_mem_pkt_o[369] = 1'b0;
  assign data_mem_pkt_o[370] = 1'b0;
  assign data_mem_pkt_o[371] = 1'b0;
  assign data_mem_pkt_o[372] = 1'b0;
  assign data_mem_pkt_o[373] = 1'b0;
  assign data_mem_pkt_o[374] = 1'b0;
  assign data_mem_pkt_o[375] = 1'b0;
  assign data_mem_pkt_o[376] = 1'b0;
  assign data_mem_pkt_o[377] = 1'b0;
  assign data_mem_pkt_o[378] = 1'b0;
  assign data_mem_pkt_o[379] = 1'b0;
  assign data_mem_pkt_o[380] = 1'b0;
  assign data_mem_pkt_o[381] = 1'b0;
  assign data_mem_pkt_o[382] = 1'b0;
  assign data_mem_pkt_o[383] = 1'b0;
  assign data_mem_pkt_o[384] = 1'b0;
  assign data_mem_pkt_o[385] = 1'b0;
  assign data_mem_pkt_o[386] = 1'b0;
  assign data_mem_pkt_o[387] = 1'b0;
  assign data_mem_pkt_o[388] = 1'b0;
  assign data_mem_pkt_o[389] = 1'b0;
  assign data_mem_pkt_o[390] = 1'b0;
  assign data_mem_pkt_o[391] = 1'b0;
  assign data_mem_pkt_o[392] = 1'b0;
  assign data_mem_pkt_o[393] = 1'b0;
  assign data_mem_pkt_o[394] = 1'b0;
  assign data_mem_pkt_o[395] = 1'b0;
  assign data_mem_pkt_o[396] = 1'b0;
  assign data_mem_pkt_o[397] = 1'b0;
  assign data_mem_pkt_o[398] = 1'b0;
  assign data_mem_pkt_o[399] = 1'b0;
  assign data_mem_pkt_o[400] = 1'b0;
  assign data_mem_pkt_o[401] = 1'b0;
  assign data_mem_pkt_o[402] = 1'b0;
  assign data_mem_pkt_o[403] = 1'b0;
  assign data_mem_pkt_o[404] = 1'b0;
  assign data_mem_pkt_o[405] = 1'b0;
  assign data_mem_pkt_o[406] = 1'b0;
  assign data_mem_pkt_o[407] = 1'b0;
  assign data_mem_pkt_o[408] = 1'b0;
  assign data_mem_pkt_o[409] = 1'b0;
  assign data_mem_pkt_o[410] = 1'b0;
  assign data_mem_pkt_o[411] = 1'b0;
  assign data_mem_pkt_o[412] = 1'b0;
  assign data_mem_pkt_o[413] = 1'b0;
  assign data_mem_pkt_o[414] = 1'b0;
  assign data_mem_pkt_o[415] = 1'b0;
  assign data_mem_pkt_o[416] = 1'b0;
  assign data_mem_pkt_o[417] = 1'b0;
  assign data_mem_pkt_o[418] = 1'b0;
  assign data_mem_pkt_o[419] = 1'b0;
  assign data_mem_pkt_o[420] = 1'b0;
  assign data_mem_pkt_o[421] = 1'b0;
  assign data_mem_pkt_o[422] = 1'b0;
  assign data_mem_pkt_o[423] = 1'b0;
  assign data_mem_pkt_o[424] = 1'b0;
  assign data_mem_pkt_o[425] = 1'b0;
  assign data_mem_pkt_o[426] = 1'b0;
  assign data_mem_pkt_o[427] = 1'b0;
  assign data_mem_pkt_o[428] = 1'b0;
  assign data_mem_pkt_o[429] = 1'b0;
  assign data_mem_pkt_o[430] = 1'b0;
  assign data_mem_pkt_o[431] = 1'b0;
  assign data_mem_pkt_o[432] = 1'b0;
  assign data_mem_pkt_o[433] = 1'b0;
  assign data_mem_pkt_o[434] = 1'b0;
  assign data_mem_pkt_o[435] = 1'b0;
  assign data_mem_pkt_o[436] = 1'b0;
  assign data_mem_pkt_o[437] = 1'b0;
  assign data_mem_pkt_o[438] = 1'b0;
  assign data_mem_pkt_o[439] = 1'b0;
  assign data_mem_pkt_o[440] = 1'b0;
  assign data_mem_pkt_o[441] = 1'b0;
  assign data_mem_pkt_o[442] = 1'b0;
  assign data_mem_pkt_o[443] = 1'b0;
  assign data_mem_pkt_o[444] = 1'b0;
  assign data_mem_pkt_o[445] = 1'b0;
  assign data_mem_pkt_o[446] = 1'b0;
  assign data_mem_pkt_o[447] = 1'b0;
  assign data_mem_pkt_o[448] = 1'b0;
  assign data_mem_pkt_o[449] = 1'b0;
  assign data_mem_pkt_o[450] = 1'b0;
  assign data_mem_pkt_o[451] = 1'b0;
  assign data_mem_pkt_o[452] = 1'b0;
  assign data_mem_pkt_o[453] = 1'b0;
  assign data_mem_pkt_o[454] = 1'b0;
  assign data_mem_pkt_o[455] = 1'b0;
  assign data_mem_pkt_o[456] = 1'b0;
  assign data_mem_pkt_o[457] = 1'b0;
  assign data_mem_pkt_o[458] = 1'b0;
  assign data_mem_pkt_o[459] = 1'b0;
  assign data_mem_pkt_o[460] = 1'b0;
  assign data_mem_pkt_o[461] = 1'b0;
  assign data_mem_pkt_o[462] = 1'b0;
  assign data_mem_pkt_o[463] = 1'b0;
  assign data_mem_pkt_o[464] = 1'b0;
  assign data_mem_pkt_o[465] = 1'b0;
  assign data_mem_pkt_o[466] = 1'b0;
  assign data_mem_pkt_o[467] = 1'b0;
  assign data_mem_pkt_o[468] = 1'b0;
  assign data_mem_pkt_o[469] = 1'b0;
  assign data_mem_pkt_o[470] = 1'b0;
  assign data_mem_pkt_o[471] = 1'b0;
  assign data_mem_pkt_o[472] = 1'b0;
  assign data_mem_pkt_o[473] = 1'b0;
  assign data_mem_pkt_o[474] = 1'b0;
  assign data_mem_pkt_o[475] = 1'b0;
  assign data_mem_pkt_o[476] = 1'b0;
  assign data_mem_pkt_o[477] = 1'b0;
  assign data_mem_pkt_o[478] = 1'b0;
  assign data_mem_pkt_o[479] = 1'b0;
  assign data_mem_pkt_o[480] = 1'b0;
  assign data_mem_pkt_o[481] = 1'b0;
  assign data_mem_pkt_o[482] = 1'b0;
  assign data_mem_pkt_o[483] = 1'b0;
  assign data_mem_pkt_o[484] = 1'b0;
  assign data_mem_pkt_o[485] = 1'b0;
  assign data_mem_pkt_o[486] = 1'b0;
  assign data_mem_pkt_o[487] = 1'b0;
  assign data_mem_pkt_o[488] = 1'b0;
  assign data_mem_pkt_o[489] = 1'b0;
  assign data_mem_pkt_o[490] = 1'b0;
  assign data_mem_pkt_o[491] = 1'b0;
  assign data_mem_pkt_o[492] = 1'b0;
  assign data_mem_pkt_o[493] = 1'b0;
  assign data_mem_pkt_o[494] = 1'b0;
  assign data_mem_pkt_o[495] = 1'b0;
  assign data_mem_pkt_o[496] = 1'b0;
  assign data_mem_pkt_o[497] = 1'b0;
  assign data_mem_pkt_o[498] = 1'b0;
  assign data_mem_pkt_o[499] = 1'b0;
  assign data_mem_pkt_o[500] = 1'b0;
  assign data_mem_pkt_o[501] = 1'b0;
  assign data_mem_pkt_o[502] = 1'b0;
  assign data_mem_pkt_o[503] = 1'b0;
  assign data_mem_pkt_o[504] = 1'b0;
  assign data_mem_pkt_o[505] = 1'b0;
  assign data_mem_pkt_o[506] = 1'b0;
  assign data_mem_pkt_o[507] = 1'b0;
  assign data_mem_pkt_o[508] = 1'b0;
  assign data_mem_pkt_o[509] = 1'b0;
  assign data_mem_pkt_o[510] = 1'b0;
  assign data_mem_pkt_o[511] = 1'b0;
  assign data_mem_pkt_o[512] = 1'b0;
  assign lce_resp_o[23] = 1'b0;
  assign lce_tr_resp_o[537] = lce_id_i[0];
  assign lce_data_resp_o[535] = lce_id_i[0];
  assign lce_resp_o[24] = lce_id_i[0];
  assign N31 = N28 & N29;
  assign N32 = N31 & N30;
  assign N33 = state_r[2] | state_r[1];
  assign N34 = N33 | N30;
  assign N36 = state_r[2] | N29;
  assign N37 = N36 | state_r[0];
  assign N39 = state_r[2] | N29;
  assign N40 = N39 | N30;
  assign N42 = N28 | state_r[1];
  assign N43 = N42 | state_r[0];
  assign N45 = N28 | state_r[1];
  assign N46 = N45 | N30;
  assign N48 = state_r[2] & state_r[1];
  assign N49 = N86 & N75;
  assign N50 = lce_cmd_i[33] | lce_cmd_i[32];
  assign N51 = N50 | N75;
  assign N68 = N70 | lce_cmd_i[31];
  assign N70 = lce_cmd_i[33] | N80;
  assign N71 = N70 | N75;
  assign N73 = N76 | lce_cmd_i[31];
  assign N76 = N79 | lce_cmd_i[32];
  assign N77 = N76 | N75;
  assign N81 = N79 | N80;
  assign N82 = N81 | lce_cmd_i[31];
  assign N84 = lce_cmd_i[33] & lce_cmd_i[32];
  assign N85 = N84 & lce_cmd_i[31];
  assign N86 = N79 & N80;
  assign N698 = (N690)? dirty_i[0] : 
                (N692)? dirty_i[1] : 
                (N694)? dirty_i[2] : 
                (N696)? dirty_i[3] : 
                (N691)? dirty_i[4] : 
                (N693)? dirty_i[5] : 
                (N695)? dirty_i[6] : 
                (N697)? dirty_i[7] : 1'b0;
  assign N1604 = state_r[1] | state_r[2];
  assign lce_sync_done_o = state_r[0] | N1604;
  assign N1606 = ~sync_ack_count_r[0];
  assign N55 = sync_ack_count_r[0] ^ 1'b1;
  assign N58 = (N0)? lce_cmd_i[34] : 
               (N1)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N0 = N49;
  assign N1 = N52;
  assign N2 = N53;
  assign N59 = (N0)? lce_cmd_v_i : 
               (N1)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N60 = (N0)? lce_resp_yumi_i : 
               (N1)? N57 : 
               (N2)? 1'b0 : 1'b0;
  assign { N66, N65, N64, N63, N62, N61 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N1)? lce_cmd_i[20:15] : 
                                            (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = (N0)? 1'b0 : 
               (N1)? lce_cmd_v_i : 
               (N2)? 1'b0 : 1'b0;
  assign N90 = (N3)? 1'b0 : 
               (N4)? lce_cmd_v_i : 1'b0;
  assign N3 = invalidated_tag_r;
  assign N4 = N89;
  assign N93 = (N5)? 1'b0 : 
               (N1237)? 1'b1 : 
               (N92)? tag_mem_pkt_yumi_i : 1'b0;
  assign N5 = lce_resp_yumi_i;
  assign { N103, N102, N101, N100, N99, N98, N97, N96, N95 } = (N6)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                                               (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N69;
  assign N7 = N72;
  assign N8 = N74;
  assign N9 = N78;
  assign N10 = N83;
  assign N11 = N87;
  assign N104 = (N6)? lce_cmd_v_i : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign { N106, N105 } = (N6)? { data_mem_pkt_yumi_i, N88 } : 
                          (N7)? { stat_mem_pkt_yumi_i, 1'b1 } : 1'b0;
  assign { N116, N115, N114, N113, N112, N111, N110, N109, N108, N107 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N7)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b1 } : 
                                                                          (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N117 = (N6)? 1'b0 : 
                (N7)? lce_cmd_v_i : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign { N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                  (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                  (N8)? { lce_cmd_i[20:15], lce_cmd_i[8:4], lce_cmd_i[30:21], 1'b1 } : 
                                                                                                                                                  (N9)? { lce_cmd_i[20:15], lce_cmd_i[8:4], lce_cmd_i[30:21], 1'b1 } : 
                                                                                                                                                  (N10)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                  (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N140 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? lce_cmd_v_i : 
                (N9)? lce_cmd_v_i : 
                (N10)? N90 : 
                (N11)? 1'b0 : 1'b0;
  assign N141 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? tag_mem_pkt_yumi_i : 
                (N9)? tag_mem_pkt_yumi_i : 
                (N10)? lce_resp_yumi_i : 
                (N11)? 1'b0 : 1'b0;
  assign N142 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? tag_mem_pkt_yumi_i : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign N143 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? tag_mem_pkt_yumi_i : 
                (N10)? 1'b0 : 
                (N11)? 1'b0 : 1'b0;
  assign { N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N10)? { lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9] } : 
                                                                                                                                                              (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N168 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? N94 : 
                (N11)? 1'b0 : 1'b0;
  assign { N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171 } = (N12)? data_buf_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? data_mem_data_i : 1'b0;
  assign N12 = tr_data_buffered_r;
  assign N13 = N170;
  assign N699 = ~N698;
  assign N710 = (N14)? 1'b0 : 
                (N1241)? 1'b1 : 
                (N709)? wb_data_read_r : 1'b0;
  assign N14 = lce_data_resp_done;
  assign N713 = (N14)? 1'b0 : 
                (N1242)? 1'b1 : 
                (N712)? data_mem_pkt_yumi_i : 1'b0;
  assign N716 = (N15)? 1'b0 : 
                (N16)? N715 : 1'b0;
  assign N15 = wb_dirty_cleared_r;
  assign N16 = N714;
  assign N719 = (N14)? 1'b0 : 
                (N1243)? 1'b1 : 
                (N718)? stat_mem_pkt_yumi_i : 1'b0;
  assign { N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721 } = (N17)? data_buf_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N18)? data_mem_data_i : 1'b0;
  assign N17 = wb_data_buffered_r;
  assign N18 = N720;
  assign stat_mem_pkt_o[0] = (N19)? N107 : 
                             (N1235)? 1'b0 : 1'b0;
  assign N19 = N35;
  assign stat_mem_pkt_o[10:2] = (N20)? { N66, N65, N64, N63, N62, N61, 1'b0, 1'b0, 1'b0 } : 
                                (N19)? { N116, N115, N114, N113, N112, N111, N110, N109, N108 } : 
                                (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N23)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = N32;
  assign N21 = N38;
  assign N22 = N41;
  assign N23 = stat_mem_pkt_o[1];
  assign N24 = N47;
  assign N25 = N48;
  assign stat_mem_pkt_v_o = (N20)? N67 : 
                            (N19)? N117 : 
                            (N21)? 1'b0 : 
                            (N22)? 1'b0 : 
                            (N23)? N716 : 
                            (N24)? 1'b0 : 
                            (N25)? 1'b0 : 1'b0;
  assign { lce_resp_o[25:25], lce_resp_o[22:0] } = (N20)? { N58, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N19)? { N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144 } : 
                                                   (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_resp_v_o = (N20)? N59 : 
                        (N19)? N168 : 
                        (N21)? 1'b0 : 
                        (N22)? 1'b0 : 
                        (N23)? 1'b0 : 
                        (N24)? 1'b0 : 
                        (N25)? 1'b0 : 1'b0;
  assign lce_cmd_yumi_o = (N20)? N60 : 
                          (N19)? N141 : 
                          (N21)? lce_tr_resp_done : 
                          (N22)? 1'b0 : 
                          (N23)? lce_data_resp_done : 
                          (N24)? lce_data_resp_done : 
                          (N25)? 1'b0 : 1'b0;
  assign state_n = (N20)? { 1'b0, 1'b0, N56 } : 
                   (N19)? { 1'b0, N106, N105 } : 
                   (N21)? { 1'b0, N169, lce_tr_resp_done } : 
                   (N22)? { 1'b1, 1'b0, N699 } : 
                   (N23)? { N1234, 1'b0, lce_data_resp_done } : 
                   (N24)? { N1234, 1'b0, 1'b1 } : 
                   (N25)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_o = (N20)? { N66, N65, N64, N63, N62, N61, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N19)? { N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N83 } : 
                         (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_v_o = (N20)? N67 : 
                           (N19)? N140 : 
                           (N21)? 1'b0 : 
                           (N22)? 1'b0 : 
                           (N23)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N25)? 1'b0 : 1'b0;
  assign data_mem_pkt_o[521:513] = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N19)? { N103, N102, N101, N100, N99, N98, N97, N96, N95 } : 
                                   (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N23)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                   (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                   (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_mem_pkt_v_o = (N20)? 1'b0 : 
                            (N19)? N104 : 
                            (N21)? 1'b0 : 
                            (N22)? 1'b0 : 
                            (N23)? N700 : 
                            (N24)? 1'b0 : 
                            (N25)? 1'b0 : 1'b0;
  assign tag_set_o = (N20)? 1'b0 : 
                     (N19)? N142 : 
                     (N21)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N25)? 1'b0 : 1'b0;
  assign tag_set_wakeup_o = (N20)? 1'b0 : 
                            (N19)? N143 : 
                            (N21)? 1'b0 : 
                            (N22)? 1'b0 : 
                            (N23)? 1'b0 : 
                            (N24)? 1'b0 : 
                            (N25)? 1'b0 : 1'b0;
  assign { lce_tr_resp_o[538:538], lce_tr_resp_o[536:0] } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N21)? { lce_cmd_i[3:0], lce_cmd_i[30:9], N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171 } : 
                                                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                            (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_tr_resp_v_o = (N20)? 1'b0 : 
                           (N19)? 1'b0 : 
                           (N21)? 1'b1 : 
                           (N22)? 1'b0 : 
                           (N23)? 1'b0 : 
                           (N24)? 1'b0 : 
                           (N25)? 1'b0 : 1'b0;
  assign { lce_data_resp_o[536:536], lce_data_resp_o[534:0] } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N23)? { lce_cmd_i[34:34], 1'b0, lce_cmd_i[30:9], N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721 } : 
                                                                (N24)? { lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_resp_v_o = (N20)? 1'b0 : 
                             (N19)? 1'b0 : 
                             (N21)? 1'b0 : 
                             (N22)? 1'b0 : 
                             (N23)? N1233 : 
                             (N24)? 1'b1 : 
                             (N25)? 1'b0 : 1'b0;
  assign { N1247, N1246, N1245 } = (N26)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N27)? state_n : 1'b0;
  assign N26 = reset_i;
  assign N27 = N1244;
  assign N1248 = (N26)? 1'b0 : 
                 (N27)? N55 : 1'b0;
  assign N1249 = (N26)? 1'b0 : 
                 (N27)? N169 : 1'b0;
  assign N1250 = (N26)? 1'b0 : 
                 (N27)? N710 : 1'b0;
  assign N1251 = (N26)? 1'b0 : 
                 (N27)? N713 : 1'b0;
  assign N1252 = (N26)? 1'b0 : 
                 (N27)? N719 : 1'b0;
  assign N1253 = (N26)? 1'b0 : 
                 (N27)? N93 : 1'b0;
  assign lce_tr_resp_done = lce_tr_resp_v_o & lce_tr_resp_ready_i;
  assign lce_data_resp_done = lce_data_resp_ready_i & lce_data_resp_v_o;
  assign N28 = ~state_r[2];
  assign N29 = ~state_r[1];
  assign N30 = ~state_r[0];
  assign N35 = ~N34;
  assign N38 = ~N37;
  assign N41 = ~N40;
  assign N44 = ~N43;
  assign N47 = ~N46;
  assign stat_mem_pkt_o[1] = N44;
  assign N52 = ~N51;
  assign N53 = lce_cmd_i[33] | lce_cmd_i[32];
  assign N54 = ~lce_resp_yumi_i;
  assign N56 = N1606 & lce_resp_yumi_i;
  assign N57 = tag_mem_pkt_yumi_i & stat_mem_pkt_yumi_i;
  assign N69 = ~N68;
  assign N72 = ~N71;
  assign N74 = ~N73;
  assign N75 = ~lce_cmd_i[31];
  assign N78 = ~N77;
  assign N79 = ~lce_cmd_i[33];
  assign N80 = ~lce_cmd_i[32];
  assign N83 = ~N82;
  assign N87 = N85 | N86;
  assign N88 = ~data_mem_pkt_yumi_i;
  assign N89 = ~invalidated_tag_r;
  assign N91 = invalidated_tag_r | lce_resp_yumi_i;
  assign N92 = ~N91;
  assign N94 = invalidated_tag_r | tag_mem_pkt_yumi_i;
  assign N169 = ~lce_tr_resp_done;
  assign N170 = ~tr_data_buffered_r;
  assign N683 = ~lce_cmd_i[6];
  assign N684 = ~lce_cmd_i[7];
  assign N685 = N683 & N684;
  assign N686 = N683 & lce_cmd_i[7];
  assign N687 = lce_cmd_i[6] & N684;
  assign N688 = lce_cmd_i[6] & lce_cmd_i[7];
  assign N689 = ~lce_cmd_i[8];
  assign N690 = N685 & N689;
  assign N691 = N685 & lce_cmd_i[8];
  assign N692 = N687 & N689;
  assign N693 = N687 & lce_cmd_i[8];
  assign N694 = N686 & N689;
  assign N695 = N686 & lce_cmd_i[8];
  assign N696 = N688 & N689;
  assign N697 = N688 & lce_cmd_i[8];
  assign N700 = ~wb_data_read_r;
  assign N701 = ~N1239;
  assign N702 = N701;
  assign N703 = N701;
  assign N704 = N701;
  assign N705 = N701;
  assign N706 = N701;
  assign N707 = N701;
  assign N708 = wb_data_buffered_r | lce_data_resp_done;
  assign N709 = ~N708;
  assign N711 = wb_data_read_r | lce_data_resp_done;
  assign N712 = ~N711;
  assign N714 = ~wb_dirty_cleared_r;
  assign N715 = wb_data_read_r | data_mem_pkt_yumi_i;
  assign N717 = wb_dirty_cleared_r | lce_data_resp_done;
  assign N718 = ~N717;
  assign N720 = ~wb_data_buffered_r;
  assign N1233 = wb_data_read_r & N1607;
  assign N1607 = wb_dirty_cleared_r | stat_mem_pkt_yumi_i;
  assign N1234 = ~lce_data_resp_done;
  assign N1235 = N34;
  assign N1236 = ~lce_resp_yumi_i;
  assign N1237 = invalidated_tag_r & N1236;
  assign N1238 = ~wb_data_buffered_r;
  assign N1239 = wb_data_read_r & N1238;
  assign N1240 = ~lce_data_resp_done;
  assign N1241 = wb_data_buffered_r & N1240;
  assign N1242 = wb_data_read_r & N1240;
  assign N1243 = wb_dirty_cleared_r & N1240;
  assign N1244 = ~reset_i;
  assign N1254 = N32 & N1244;
  assign N1255 = N35 & N1244;
  assign N1256 = N1254 | N1255;
  assign N1257 = N38 & N1244;
  assign N1258 = tr_data_buffered_r & N1257;
  assign N1259 = N1256 | N1258;
  assign N1260 = N41 & N1244;
  assign N1261 = N1259 | N1260;
  assign N1262 = stat_mem_pkt_o[1] & N1244;
  assign N1263 = N702 & N1262;
  assign N1264 = N1261 | N1263;
  assign N1265 = N47 & N1244;
  assign N1266 = N1264 | N1265;
  assign N1267 = N48 & N1244;
  assign N1268 = N1266 | N1267;
  assign N1269 = ~N1268;
  assign N1270 = N1244 & N1269;
  assign N1271 = N32 & N1244;
  assign N1272 = N35 & N1244;
  assign N1273 = N1271 | N1272;
  assign N1274 = N38 & N1244;
  assign N1275 = tr_data_buffered_r & N1274;
  assign N1276 = N1273 | N1275;
  assign N1277 = N41 & N1244;
  assign N1278 = N1276 | N1277;
  assign N1279 = stat_mem_pkt_o[1] & N1244;
  assign N1280 = N702 & N1279;
  assign N1281 = N1278 | N1280;
  assign N1282 = N47 & N1244;
  assign N1283 = N1281 | N1282;
  assign N1284 = N48 & N1244;
  assign N1285 = N1283 | N1284;
  assign N1286 = ~N1285;
  assign N1287 = N1244 & N1286;
  assign N1288 = N32 & N1244;
  assign N1289 = N35 & N1244;
  assign N1290 = N1288 | N1289;
  assign N1291 = N38 & N1244;
  assign N1292 = tr_data_buffered_r & N1291;
  assign N1293 = N1290 | N1292;
  assign N1294 = N41 & N1244;
  assign N1295 = N1293 | N1294;
  assign N1296 = stat_mem_pkt_o[1] & N1244;
  assign N1297 = N702 & N1296;
  assign N1298 = N1295 | N1297;
  assign N1299 = N47 & N1244;
  assign N1300 = N1298 | N1299;
  assign N1301 = N48 & N1244;
  assign N1302 = N1300 | N1301;
  assign N1303 = ~N1302;
  assign N1304 = N1244 & N1303;
  assign N1305 = N32 & N1244;
  assign N1306 = N35 & N1244;
  assign N1307 = N1305 | N1306;
  assign N1308 = N38 & N1244;
  assign N1309 = tr_data_buffered_r & N1308;
  assign N1310 = N1307 | N1309;
  assign N1311 = N41 & N1244;
  assign N1312 = N1310 | N1311;
  assign N1313 = stat_mem_pkt_o[1] & N1244;
  assign N1314 = N702 & N1313;
  assign N1315 = N1312 | N1314;
  assign N1316 = N47 & N1244;
  assign N1317 = N1315 | N1316;
  assign N1318 = N48 & N1244;
  assign N1319 = N1317 | N1318;
  assign N1320 = ~N1319;
  assign N1321 = N1244 & N1320;
  assign N1322 = N32 & N1244;
  assign N1323 = N35 & N1244;
  assign N1324 = N1322 | N1323;
  assign N1325 = N38 & N1244;
  assign N1326 = tr_data_buffered_r & N1325;
  assign N1327 = N1324 | N1326;
  assign N1328 = N41 & N1244;
  assign N1329 = N1327 | N1328;
  assign N1330 = stat_mem_pkt_o[1] & N1244;
  assign N1331 = N702 & N1330;
  assign N1332 = N1329 | N1331;
  assign N1333 = N47 & N1244;
  assign N1334 = N1332 | N1333;
  assign N1335 = N48 & N1244;
  assign N1336 = N1334 | N1335;
  assign N1337 = ~N1336;
  assign N1338 = N1244 & N1337;
  assign N1339 = N32 & N1244;
  assign N1340 = N35 & N1244;
  assign N1341 = N1339 | N1340;
  assign N1342 = N38 & N1244;
  assign N1343 = tr_data_buffered_r & N1342;
  assign N1344 = N1341 | N1343;
  assign N1345 = N41 & N1244;
  assign N1346 = N1344 | N1345;
  assign N1347 = stat_mem_pkt_o[1] & N1244;
  assign N1348 = N702 & N1347;
  assign N1349 = N1346 | N1348;
  assign N1350 = N47 & N1244;
  assign N1351 = N1349 | N1350;
  assign N1352 = N48 & N1244;
  assign N1353 = N1351 | N1352;
  assign N1354 = ~N1353;
  assign N1355 = N1244 & N1354;
  assign N1356 = N1346 | N1331;
  assign N1357 = N1356 | N1350;
  assign N1358 = N1357 | N1352;
  assign N1359 = ~N1358;
  assign N1360 = N1244 & N1359;
  assign N1361 = N1341 | N1326;
  assign N1362 = N1361 | N1345;
  assign N1363 = N1362 | N1331;
  assign N1364 = N1363 | N1350;
  assign N1365 = N1364 | N1352;
  assign N1366 = ~N1365;
  assign N1367 = N1244 & N1366;
  assign N1368 = N1361 | N1328;
  assign N1369 = N1368 | N1331;
  assign N1370 = N1369 | N1333;
  assign N1371 = N1370 | N1335;
  assign N1372 = ~N1371;
  assign N1373 = N1244 & N1372;
  assign N1374 = N1322 | N1340;
  assign N1375 = N1374 | N1326;
  assign N1376 = N1375 | N1328;
  assign N1377 = N1376 | N1331;
  assign N1378 = N1377 | N1333;
  assign N1379 = N1378 | N1335;
  assign N1380 = ~N1379;
  assign N1381 = N1244 & N1380;
  assign N1382 = N703 & N1330;
  assign N1383 = N1329 | N1382;
  assign N1384 = N1383 | N1333;
  assign N1385 = N1384 | N1335;
  assign N1386 = ~N1385;
  assign N1387 = N1244 & N1386;
  assign N1388 = N703 & N1313;
  assign N1389 = N1329 | N1388;
  assign N1390 = N1389 | N1333;
  assign N1391 = N1390 | N1335;
  assign N1392 = ~N1391;
  assign N1393 = N1244 & N1392;
  assign N1394 = N1324 | N1309;
  assign N1395 = N1394 | N1328;
  assign N1396 = N1395 | N1388;
  assign N1397 = N1396 | N1333;
  assign N1398 = N1397 | N1335;
  assign N1399 = ~N1398;
  assign N1400 = N1244 & N1399;
  assign N1401 = N1394 | N1311;
  assign N1402 = N1401 | N1388;
  assign N1403 = N1402 | N1316;
  assign N1404 = N1403 | N1318;
  assign N1405 = ~N1404;
  assign N1406 = N1244 & N1405;
  assign N1407 = N1305 | N1323;
  assign N1408 = N1407 | N1309;
  assign N1409 = N1408 | N1311;
  assign N1410 = N1409 | N1388;
  assign N1411 = N1410 | N1316;
  assign N1412 = N1411 | N1318;
  assign N1413 = ~N1412;
  assign N1414 = N1244 & N1413;
  assign N1415 = N1312 | N1388;
  assign N1416 = N1415 | N1316;
  assign N1417 = N1416 | N1318;
  assign N1418 = ~N1417;
  assign N1419 = N1244 & N1418;
  assign N1420 = N704 & N1313;
  assign N1421 = N1312 | N1420;
  assign N1422 = N1421 | N1316;
  assign N1423 = N1422 | N1318;
  assign N1424 = ~N1423;
  assign N1425 = N1244 & N1424;
  assign N1426 = N704 & N1296;
  assign N1427 = N1312 | N1426;
  assign N1428 = N1427 | N1316;
  assign N1429 = N1428 | N1318;
  assign N1430 = ~N1429;
  assign N1431 = N1244 & N1430;
  assign N1432 = N1307 | N1292;
  assign N1433 = N1432 | N1311;
  assign N1434 = N1433 | N1426;
  assign N1435 = N1434 | N1316;
  assign N1436 = N1435 | N1318;
  assign N1437 = ~N1436;
  assign N1438 = N1244 & N1437;
  assign N1439 = N1432 | N1294;
  assign N1440 = N1439 | N1426;
  assign N1441 = N1440 | N1299;
  assign N1442 = N1441 | N1301;
  assign N1443 = ~N1442;
  assign N1444 = N1244 & N1443;
  assign N1445 = N1288 | N1306;
  assign N1446 = N1445 | N1292;
  assign N1447 = N1446 | N1294;
  assign N1448 = N1447 | N1426;
  assign N1449 = N1448 | N1299;
  assign N1450 = N1449 | N1301;
  assign N1451 = ~N1450;
  assign N1452 = N1244 & N1451;
  assign N1453 = N1295 | N1426;
  assign N1454 = N1453 | N1299;
  assign N1455 = N1454 | N1301;
  assign N1456 = ~N1455;
  assign N1457 = N1244 & N1456;
  assign N1458 = N705 & N1296;
  assign N1459 = N1295 | N1458;
  assign N1460 = N1459 | N1299;
  assign N1461 = N1460 | N1301;
  assign N1462 = ~N1461;
  assign N1463 = N1244 & N1462;
  assign N1464 = N705 & N1279;
  assign N1465 = N1295 | N1464;
  assign N1466 = N1465 | N1299;
  assign N1467 = N1466 | N1301;
  assign N1468 = ~N1467;
  assign N1469 = N1244 & N1468;
  assign N1470 = N1290 | N1275;
  assign N1471 = N1470 | N1294;
  assign N1472 = N1471 | N1464;
  assign N1473 = N1472 | N1299;
  assign N1474 = N1473 | N1301;
  assign N1475 = ~N1474;
  assign N1476 = N1244 & N1475;
  assign N1477 = N1470 | N1277;
  assign N1478 = N1477 | N1464;
  assign N1479 = N1478 | N1282;
  assign N1480 = N1479 | N1284;
  assign N1481 = ~N1480;
  assign N1482 = N1244 & N1481;
  assign N1483 = N1271 | N1289;
  assign N1484 = N1483 | N1275;
  assign N1485 = N1484 | N1277;
  assign N1486 = N1485 | N1464;
  assign N1487 = N1486 | N1282;
  assign N1488 = N1487 | N1284;
  assign N1489 = ~N1488;
  assign N1490 = N1244 & N1489;
  assign N1491 = N1278 | N1464;
  assign N1492 = N1491 | N1282;
  assign N1493 = N1492 | N1284;
  assign N1494 = ~N1493;
  assign N1495 = N1244 & N1494;
  assign N1496 = N706 & N1279;
  assign N1497 = N1278 | N1496;
  assign N1498 = N1497 | N1282;
  assign N1499 = N1498 | N1284;
  assign N1500 = ~N1499;
  assign N1501 = N1244 & N1500;
  assign N1502 = N706 & N1262;
  assign N1503 = N1278 | N1502;
  assign N1504 = N1503 | N1282;
  assign N1505 = N1504 | N1284;
  assign N1506 = ~N1505;
  assign N1507 = N1244 & N1506;
  assign N1508 = N1273 | N1258;
  assign N1509 = N1508 | N1277;
  assign N1510 = N1509 | N1502;
  assign N1511 = N1510 | N1282;
  assign N1512 = N1511 | N1284;
  assign N1513 = ~N1512;
  assign N1514 = N1244 & N1513;
  assign N1515 = N1508 | N1260;
  assign N1516 = N1515 | N1502;
  assign N1517 = N1516 | N1265;
  assign N1518 = N1517 | N1267;
  assign N1519 = ~N1518;
  assign N1520 = N1244 & N1519;
  assign N1521 = N1254 | N1272;
  assign N1522 = N1521 | N1258;
  assign N1523 = N1522 | N1260;
  assign N1524 = N1523 | N1502;
  assign N1525 = N1524 | N1265;
  assign N1526 = N1525 | N1267;
  assign N1527 = ~N1526;
  assign N1528 = N1244 & N1527;
  assign N1529 = N1261 | N1502;
  assign N1530 = N1529 | N1265;
  assign N1531 = N1530 | N1267;
  assign N1532 = ~N1531;
  assign N1533 = N1244 & N1532;
  assign N1534 = N707 & N1262;
  assign N1535 = N1261 | N1534;
  assign N1536 = N1535 | N1265;
  assign N1537 = N1536 | N1267;
  assign N1538 = ~N1537;
  assign N1539 = N1244 & N1538;
  assign N1540 = N705 & N1262;
  assign N1541 = N1261 | N1540;
  assign N1542 = N1541 | N1265;
  assign N1543 = N1542 | N1267;
  assign N1544 = ~N1543;
  assign N1545 = N1244 & N1544;
  assign N1546 = N704 & N1262;
  assign N1547 = N1261 | N1546;
  assign N1548 = N1547 | N1265;
  assign N1549 = N1548 | N1267;
  assign N1550 = ~N1549;
  assign N1551 = N1244 & N1550;
  assign N1552 = N703 & N1262;
  assign N1553 = N1261 | N1552;
  assign N1554 = N1553 | N1265;
  assign N1555 = N1554 | N1267;
  assign N1556 = ~N1555;
  assign N1557 = N1244 & N1556;
  assign N1558 = N52 & N1254;
  assign N1559 = N53 & N1254;
  assign N1560 = N1558 | N1559;
  assign N1561 = N74 & N1255;
  assign N1562 = N1560 | N1561;
  assign N1563 = N78 & N1255;
  assign N1564 = N1562 | N1563;
  assign N1565 = N83 & N1255;
  assign N1566 = N1564 | N1565;
  assign N1567 = N87 & N1255;
  assign N1568 = N1566 | N1567;
  assign N1569 = ~N1568;
  assign N1570 = N49 & N1254;
  assign N1571 = N54 & N1570;
  assign N1572 = N1571 | N1558;
  assign N1573 = N1572 | N1559;
  assign N1574 = N1573 | N1255;
  assign N1575 = N1574 | N1257;
  assign N1576 = N1575 | N1260;
  assign N1577 = N1576 | N1262;
  assign N1578 = N1577 | N1265;
  assign N1579 = N1578 | N1267;
  assign N1580 = ~N1579;
  assign N1581 = N1256 | N1260;
  assign N1582 = N1581 | N1262;
  assign N1583 = N1582 | N1265;
  assign N1584 = N1583 | N1267;
  assign N1585 = ~N1584;
  assign N1586 = N1256 | N1257;
  assign N1587 = N1586 | N1260;
  assign N1588 = N1587 | N1265;
  assign N1589 = N1588 | N1267;
  assign N1590 = ~N1589;
  assign N1591 = N69 & N1255;
  assign N1592 = N1254 | N1591;
  assign N1593 = N72 & N1255;
  assign N1594 = N1592 | N1593;
  assign N1595 = N1594 | N1561;
  assign N1596 = N1595 | N1563;
  assign N1597 = N1596 | N1567;
  assign N1598 = N1597 | N1257;
  assign N1599 = N1598 | N1260;
  assign N1600 = N1599 | N1262;
  assign N1601 = N1600 | N1265;
  assign N1602 = N1601 | N1267;
  assign N1603 = ~N1602;

  always @(posedge clk_i) begin
    if(N1270) begin
      { data_buf_r[511:511], data_buf_r[0:0] } <= { data_mem_data_i[511:511], data_mem_data_i[0:0] };
    end 
    if(N1287) begin
      { data_buf_r[510:510] } <= { data_mem_data_i[510:510] };
    end 
    if(N1304) begin
      { data_buf_r[509:509] } <= { data_mem_data_i[509:509] };
    end 
    if(N1321) begin
      { data_buf_r[508:508] } <= { data_mem_data_i[508:508] };
    end 
    if(N1338) begin
      { data_buf_r[507:507], data_buf_r[472:413] } <= { data_mem_data_i[507:507], data_mem_data_i[472:413] };
    end 
    if(N1355) begin
      { data_buf_r[506:492] } <= { data_mem_data_i[506:492] };
    end 
    if(N1360) begin
      { data_buf_r[491:490] } <= { data_mem_data_i[491:490] };
    end 
    if(N1367) begin
      { data_buf_r[489:489] } <= { data_mem_data_i[489:489] };
    end 
    if(N1373) begin
      { data_buf_r[488:481] } <= { data_mem_data_i[488:481] };
    end 
    if(N1381) begin
      { data_buf_r[480:473] } <= { data_mem_data_i[480:473] };
    end 
    if(N1387) begin
      { data_buf_r[412:393] } <= { data_mem_data_i[412:393] };
    end 
    if(N1393) begin
      { data_buf_r[392:391] } <= { data_mem_data_i[392:391] };
    end 
    if(N1400) begin
      { data_buf_r[390:390] } <= { data_mem_data_i[390:390] };
    end 
    if(N1406) begin
      { data_buf_r[389:382] } <= { data_mem_data_i[389:382] };
    end 
    if(N1414) begin
      { data_buf_r[381:374] } <= { data_mem_data_i[381:374] };
    end 
    if(N1419) begin
      { data_buf_r[373:314] } <= { data_mem_data_i[373:314] };
    end 
    if(N1425) begin
      { data_buf_r[313:294] } <= { data_mem_data_i[313:294] };
    end 
    if(N1431) begin
      { data_buf_r[293:292] } <= { data_mem_data_i[293:292] };
    end 
    if(N1438) begin
      { data_buf_r[291:291] } <= { data_mem_data_i[291:291] };
    end 
    if(N1444) begin
      { data_buf_r[290:283] } <= { data_mem_data_i[290:283] };
    end 
    if(N1452) begin
      { data_buf_r[282:275] } <= { data_mem_data_i[282:275] };
    end 
    if(N1457) begin
      { data_buf_r[274:215] } <= { data_mem_data_i[274:215] };
    end 
    if(N1463) begin
      { data_buf_r[214:195] } <= { data_mem_data_i[214:195] };
    end 
    if(N1469) begin
      { data_buf_r[194:193] } <= { data_mem_data_i[194:193] };
    end 
    if(N1476) begin
      { data_buf_r[192:192] } <= { data_mem_data_i[192:192] };
    end 
    if(N1482) begin
      { data_buf_r[191:184] } <= { data_mem_data_i[191:184] };
    end 
    if(N1490) begin
      { data_buf_r[183:176] } <= { data_mem_data_i[183:176] };
    end 
    if(N1495) begin
      { data_buf_r[175:116] } <= { data_mem_data_i[175:116] };
    end 
    if(N1501) begin
      { data_buf_r[115:96] } <= { data_mem_data_i[115:96] };
    end 
    if(N1507) begin
      { data_buf_r[95:94] } <= { data_mem_data_i[95:94] };
    end 
    if(N1514) begin
      { data_buf_r[93:93] } <= { data_mem_data_i[93:93] };
    end 
    if(N1520) begin
      { data_buf_r[92:85] } <= { data_mem_data_i[92:85] };
    end 
    if(N1528) begin
      { data_buf_r[84:77] } <= { data_mem_data_i[84:77] };
    end 
    if(N1533) begin
      { data_buf_r[76:17], data_buf_r[4:4] } <= { data_mem_data_i[76:17], data_mem_data_i[4:4] };
    end 
    if(N1539) begin
      { data_buf_r[16:5] } <= { data_mem_data_i[16:5] };
    end 
    if(N1545) begin
      { data_buf_r[3:3] } <= { data_mem_data_i[3:3] };
    end 
    if(N1551) begin
      { data_buf_r[2:2] } <= { data_mem_data_i[2:2] };
    end 
    if(N1557) begin
      { data_buf_r[1:1] } <= { data_mem_data_i[1:1] };
    end 
    if(N1569) begin
      { state_r[2:0] } <= { N1247, N1246, N1245 };
    end 
    if(N1580) begin
      { sync_ack_count_r[0:0] } <= { N1248 };
    end 
    if(N1585) begin
      tr_data_buffered_r <= N1249;
    end 
    if(N1590) begin
      wb_data_buffered_r <= N1250;
      wb_data_read_r <= N1251;
      wb_dirty_cleared_r <= N1252;
    end 
    if(N1603) begin
      invalidated_tag_r <= N1253;
    end 
  end


endmodule