module Queue_4
(
  clk,
  reset,
  io_enq_ready,
  io_enq_valid,
  io_enq_bits_resp,
  io_enq_bits_data,
  io_enq_bits_last,
  io_enq_bits_id,
  io_enq_bits_user,
  io_deq_ready,
  io_deq_valid,
  io_deq_bits_resp,
  io_deq_bits_data,
  io_deq_bits_last,
  io_deq_bits_id,
  io_deq_bits_user,
  io_count
);

  input [1:0] io_enq_bits_resp;
  input [63:0] io_enq_bits_data;
  input [5:0] io_enq_bits_id;
  output [1:0] io_deq_bits_resp;
  output [63:0] io_deq_bits_data;
  output [5:0] io_deq_bits_id;
  output [3:0] io_count;
  input clk;
  input reset;
  input io_enq_valid;
  input io_enq_bits_last;
  input io_enq_bits_user;
  input io_deq_ready;
  output io_enq_ready;
  output io_deq_valid;
  output io_deq_bits_last;
  output io_deq_bits_user;
  wire [1:0] io_deq_bits_resp;
  wire [63:0] io_deq_bits_data;
  wire [5:0] io_deq_bits_id;
  wire [3:0] io_count;
  wire io_enq_ready,io_deq_valid,io_deq_bits_last,io_deq_bits_user,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,do_deq,do_enq,ptr_match,T9,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,empty,T23,full,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74;
  wire [2:0] T3,T6;
  reg [2:0] R1,R4;
  reg maybe_full;
  reg [591:0] ram;
  assign ptr_match = R4 == R1;
  assign T9 = do_enq ^ do_deq;
  assign io_deq_bits_resp[1] = (N22)? ram[73] : 
                               (N24)? ram[147] : 
                               (N26)? ram[221] : 
                               (N28)? ram[295] : 
                               (N23)? ram[369] : 
                               (N25)? ram[443] : 
                               (N27)? ram[517] : 
                               (N29)? ram[591] : 1'b0;
  assign io_deq_bits_resp[0] = (N22)? ram[72] : 
                               (N24)? ram[146] : 
                               (N26)? ram[220] : 
                               (N28)? ram[294] : 
                               (N23)? ram[368] : 
                               (N25)? ram[442] : 
                               (N27)? ram[516] : 
                               (N29)? ram[590] : 1'b0;
  assign io_deq_bits_data[63] = (N22)? ram[71] : 
                                (N24)? ram[145] : 
                                (N26)? ram[219] : 
                                (N28)? ram[293] : 
                                (N23)? ram[367] : 
                                (N25)? ram[441] : 
                                (N27)? ram[515] : 
                                (N29)? ram[589] : 1'b0;
  assign io_deq_bits_data[62] = (N22)? ram[70] : 
                                (N24)? ram[144] : 
                                (N26)? ram[218] : 
                                (N28)? ram[292] : 
                                (N23)? ram[366] : 
                                (N25)? ram[440] : 
                                (N27)? ram[514] : 
                                (N29)? ram[588] : 1'b0;
  assign io_deq_bits_data[61] = (N22)? ram[69] : 
                                (N24)? ram[143] : 
                                (N26)? ram[217] : 
                                (N28)? ram[291] : 
                                (N23)? ram[365] : 
                                (N25)? ram[439] : 
                                (N27)? ram[513] : 
                                (N29)? ram[587] : 1'b0;
  assign io_deq_bits_data[60] = (N22)? ram[68] : 
                                (N24)? ram[142] : 
                                (N26)? ram[216] : 
                                (N28)? ram[290] : 
                                (N23)? ram[364] : 
                                (N25)? ram[438] : 
                                (N27)? ram[512] : 
                                (N29)? ram[586] : 1'b0;
  assign io_deq_bits_data[59] = (N22)? ram[67] : 
                                (N24)? ram[141] : 
                                (N26)? ram[215] : 
                                (N28)? ram[289] : 
                                (N23)? ram[363] : 
                                (N25)? ram[437] : 
                                (N27)? ram[511] : 
                                (N29)? ram[585] : 1'b0;
  assign io_deq_bits_data[58] = (N22)? ram[66] : 
                                (N24)? ram[140] : 
                                (N26)? ram[214] : 
                                (N28)? ram[288] : 
                                (N23)? ram[362] : 
                                (N25)? ram[436] : 
                                (N27)? ram[510] : 
                                (N29)? ram[584] : 1'b0;
  assign io_deq_bits_data[57] = (N22)? ram[65] : 
                                (N24)? ram[139] : 
                                (N26)? ram[213] : 
                                (N28)? ram[287] : 
                                (N23)? ram[361] : 
                                (N25)? ram[435] : 
                                (N27)? ram[509] : 
                                (N29)? ram[583] : 1'b0;
  assign io_deq_bits_data[56] = (N22)? ram[64] : 
                                (N24)? ram[138] : 
                                (N26)? ram[212] : 
                                (N28)? ram[286] : 
                                (N23)? ram[360] : 
                                (N25)? ram[434] : 
                                (N27)? ram[508] : 
                                (N29)? ram[582] : 1'b0;
  assign io_deq_bits_data[55] = (N22)? ram[63] : 
                                (N24)? ram[137] : 
                                (N26)? ram[211] : 
                                (N28)? ram[285] : 
                                (N23)? ram[359] : 
                                (N25)? ram[433] : 
                                (N27)? ram[507] : 
                                (N29)? ram[581] : 1'b0;
  assign io_deq_bits_data[54] = (N22)? ram[62] : 
                                (N24)? ram[136] : 
                                (N26)? ram[210] : 
                                (N28)? ram[284] : 
                                (N23)? ram[358] : 
                                (N25)? ram[432] : 
                                (N27)? ram[506] : 
                                (N29)? ram[580] : 1'b0;
  assign io_deq_bits_data[53] = (N22)? ram[61] : 
                                (N24)? ram[135] : 
                                (N26)? ram[209] : 
                                (N28)? ram[283] : 
                                (N23)? ram[357] : 
                                (N25)? ram[431] : 
                                (N27)? ram[505] : 
                                (N29)? ram[579] : 1'b0;
  assign io_deq_bits_data[52] = (N22)? ram[60] : 
                                (N24)? ram[134] : 
                                (N26)? ram[208] : 
                                (N28)? ram[282] : 
                                (N23)? ram[356] : 
                                (N25)? ram[430] : 
                                (N27)? ram[504] : 
                                (N29)? ram[578] : 1'b0;
  assign io_deq_bits_data[51] = (N22)? ram[59] : 
                                (N24)? ram[133] : 
                                (N26)? ram[207] : 
                                (N28)? ram[281] : 
                                (N23)? ram[355] : 
                                (N25)? ram[429] : 
                                (N27)? ram[503] : 
                                (N29)? ram[577] : 1'b0;
  assign io_deq_bits_data[50] = (N22)? ram[58] : 
                                (N24)? ram[132] : 
                                (N26)? ram[206] : 
                                (N28)? ram[280] : 
                                (N23)? ram[354] : 
                                (N25)? ram[428] : 
                                (N27)? ram[502] : 
                                (N29)? ram[576] : 1'b0;
  assign io_deq_bits_data[49] = (N22)? ram[57] : 
                                (N24)? ram[131] : 
                                (N26)? ram[205] : 
                                (N28)? ram[279] : 
                                (N23)? ram[353] : 
                                (N25)? ram[427] : 
                                (N27)? ram[501] : 
                                (N29)? ram[575] : 1'b0;
  assign io_deq_bits_data[48] = (N22)? ram[56] : 
                                (N24)? ram[130] : 
                                (N26)? ram[204] : 
                                (N28)? ram[278] : 
                                (N23)? ram[352] : 
                                (N25)? ram[426] : 
                                (N27)? ram[500] : 
                                (N29)? ram[574] : 1'b0;
  assign io_deq_bits_data[47] = (N22)? ram[55] : 
                                (N24)? ram[129] : 
                                (N26)? ram[203] : 
                                (N28)? ram[277] : 
                                (N23)? ram[351] : 
                                (N25)? ram[425] : 
                                (N27)? ram[499] : 
                                (N29)? ram[573] : 1'b0;
  assign io_deq_bits_data[46] = (N22)? ram[54] : 
                                (N24)? ram[128] : 
                                (N26)? ram[202] : 
                                (N28)? ram[276] : 
                                (N23)? ram[350] : 
                                (N25)? ram[424] : 
                                (N27)? ram[498] : 
                                (N29)? ram[572] : 1'b0;
  assign io_deq_bits_data[45] = (N22)? ram[53] : 
                                (N24)? ram[127] : 
                                (N26)? ram[201] : 
                                (N28)? ram[275] : 
                                (N23)? ram[349] : 
                                (N25)? ram[423] : 
                                (N27)? ram[497] : 
                                (N29)? ram[571] : 1'b0;
  assign io_deq_bits_data[44] = (N22)? ram[52] : 
                                (N24)? ram[126] : 
                                (N26)? ram[200] : 
                                (N28)? ram[274] : 
                                (N23)? ram[348] : 
                                (N25)? ram[422] : 
                                (N27)? ram[496] : 
                                (N29)? ram[570] : 1'b0;
  assign io_deq_bits_data[43] = (N22)? ram[51] : 
                                (N24)? ram[125] : 
                                (N26)? ram[199] : 
                                (N28)? ram[273] : 
                                (N23)? ram[347] : 
                                (N25)? ram[421] : 
                                (N27)? ram[495] : 
                                (N29)? ram[569] : 1'b0;
  assign io_deq_bits_data[42] = (N22)? ram[50] : 
                                (N24)? ram[124] : 
                                (N26)? ram[198] : 
                                (N28)? ram[272] : 
                                (N23)? ram[346] : 
                                (N25)? ram[420] : 
                                (N27)? ram[494] : 
                                (N29)? ram[568] : 1'b0;
  assign io_deq_bits_data[41] = (N22)? ram[49] : 
                                (N24)? ram[123] : 
                                (N26)? ram[197] : 
                                (N28)? ram[271] : 
                                (N23)? ram[345] : 
                                (N25)? ram[419] : 
                                (N27)? ram[493] : 
                                (N29)? ram[567] : 1'b0;
  assign io_deq_bits_data[40] = (N22)? ram[48] : 
                                (N24)? ram[122] : 
                                (N26)? ram[196] : 
                                (N28)? ram[270] : 
                                (N23)? ram[344] : 
                                (N25)? ram[418] : 
                                (N27)? ram[492] : 
                                (N29)? ram[566] : 1'b0;
  assign io_deq_bits_data[39] = (N22)? ram[47] : 
                                (N24)? ram[121] : 
                                (N26)? ram[195] : 
                                (N28)? ram[269] : 
                                (N23)? ram[343] : 
                                (N25)? ram[417] : 
                                (N27)? ram[491] : 
                                (N29)? ram[565] : 1'b0;
  assign io_deq_bits_data[38] = (N22)? ram[46] : 
                                (N24)? ram[120] : 
                                (N26)? ram[194] : 
                                (N28)? ram[268] : 
                                (N23)? ram[342] : 
                                (N25)? ram[416] : 
                                (N27)? ram[490] : 
                                (N29)? ram[564] : 1'b0;
  assign io_deq_bits_data[37] = (N22)? ram[45] : 
                                (N24)? ram[119] : 
                                (N26)? ram[193] : 
                                (N28)? ram[267] : 
                                (N23)? ram[341] : 
                                (N25)? ram[415] : 
                                (N27)? ram[489] : 
                                (N29)? ram[563] : 1'b0;
  assign io_deq_bits_data[36] = (N22)? ram[44] : 
                                (N24)? ram[118] : 
                                (N26)? ram[192] : 
                                (N28)? ram[266] : 
                                (N23)? ram[340] : 
                                (N25)? ram[414] : 
                                (N27)? ram[488] : 
                                (N29)? ram[562] : 1'b0;
  assign io_deq_bits_data[35] = (N22)? ram[43] : 
                                (N24)? ram[117] : 
                                (N26)? ram[191] : 
                                (N28)? ram[265] : 
                                (N23)? ram[339] : 
                                (N25)? ram[413] : 
                                (N27)? ram[487] : 
                                (N29)? ram[561] : 1'b0;
  assign io_deq_bits_data[34] = (N22)? ram[42] : 
                                (N24)? ram[116] : 
                                (N26)? ram[190] : 
                                (N28)? ram[264] : 
                                (N23)? ram[338] : 
                                (N25)? ram[412] : 
                                (N27)? ram[486] : 
                                (N29)? ram[560] : 1'b0;
  assign io_deq_bits_data[33] = (N22)? ram[41] : 
                                (N24)? ram[115] : 
                                (N26)? ram[189] : 
                                (N28)? ram[263] : 
                                (N23)? ram[337] : 
                                (N25)? ram[411] : 
                                (N27)? ram[485] : 
                                (N29)? ram[559] : 1'b0;
  assign io_deq_bits_data[32] = (N22)? ram[40] : 
                                (N24)? ram[114] : 
                                (N26)? ram[188] : 
                                (N28)? ram[262] : 
                                (N23)? ram[336] : 
                                (N25)? ram[410] : 
                                (N27)? ram[484] : 
                                (N29)? ram[558] : 1'b0;
  assign io_deq_bits_data[31] = (N22)? ram[39] : 
                                (N24)? ram[113] : 
                                (N26)? ram[187] : 
                                (N28)? ram[261] : 
                                (N23)? ram[335] : 
                                (N25)? ram[409] : 
                                (N27)? ram[483] : 
                                (N29)? ram[557] : 1'b0;
  assign io_deq_bits_data[30] = (N22)? ram[38] : 
                                (N24)? ram[112] : 
                                (N26)? ram[186] : 
                                (N28)? ram[260] : 
                                (N23)? ram[334] : 
                                (N25)? ram[408] : 
                                (N27)? ram[482] : 
                                (N29)? ram[556] : 1'b0;
  assign io_deq_bits_data[29] = (N22)? ram[37] : 
                                (N24)? ram[111] : 
                                (N26)? ram[185] : 
                                (N28)? ram[259] : 
                                (N23)? ram[333] : 
                                (N25)? ram[407] : 
                                (N27)? ram[481] : 
                                (N29)? ram[555] : 1'b0;
  assign io_deq_bits_data[28] = (N22)? ram[36] : 
                                (N24)? ram[110] : 
                                (N26)? ram[184] : 
                                (N28)? ram[258] : 
                                (N23)? ram[332] : 
                                (N25)? ram[406] : 
                                (N27)? ram[480] : 
                                (N29)? ram[554] : 1'b0;
  assign io_deq_bits_data[27] = (N22)? ram[35] : 
                                (N24)? ram[109] : 
                                (N26)? ram[183] : 
                                (N28)? ram[257] : 
                                (N23)? ram[331] : 
                                (N25)? ram[405] : 
                                (N27)? ram[479] : 
                                (N29)? ram[553] : 1'b0;
  assign io_deq_bits_data[26] = (N22)? ram[34] : 
                                (N24)? ram[108] : 
                                (N26)? ram[182] : 
                                (N28)? ram[256] : 
                                (N23)? ram[330] : 
                                (N25)? ram[404] : 
                                (N27)? ram[478] : 
                                (N29)? ram[552] : 1'b0;
  assign io_deq_bits_data[25] = (N22)? ram[33] : 
                                (N24)? ram[107] : 
                                (N26)? ram[181] : 
                                (N28)? ram[255] : 
                                (N23)? ram[329] : 
                                (N25)? ram[403] : 
                                (N27)? ram[477] : 
                                (N29)? ram[551] : 1'b0;
  assign io_deq_bits_data[24] = (N22)? ram[32] : 
                                (N24)? ram[106] : 
                                (N26)? ram[180] : 
                                (N28)? ram[254] : 
                                (N23)? ram[328] : 
                                (N25)? ram[402] : 
                                (N27)? ram[476] : 
                                (N29)? ram[550] : 1'b0;
  assign io_deq_bits_data[23] = (N22)? ram[31] : 
                                (N24)? ram[105] : 
                                (N26)? ram[179] : 
                                (N28)? ram[253] : 
                                (N23)? ram[327] : 
                                (N25)? ram[401] : 
                                (N27)? ram[475] : 
                                (N29)? ram[549] : 1'b0;
  assign io_deq_bits_data[22] = (N22)? ram[30] : 
                                (N24)? ram[104] : 
                                (N26)? ram[178] : 
                                (N28)? ram[252] : 
                                (N23)? ram[326] : 
                                (N25)? ram[400] : 
                                (N27)? ram[474] : 
                                (N29)? ram[548] : 1'b0;
  assign io_deq_bits_data[21] = (N22)? ram[29] : 
                                (N24)? ram[103] : 
                                (N26)? ram[177] : 
                                (N28)? ram[251] : 
                                (N23)? ram[325] : 
                                (N25)? ram[399] : 
                                (N27)? ram[473] : 
                                (N29)? ram[547] : 1'b0;
  assign io_deq_bits_data[20] = (N22)? ram[28] : 
                                (N24)? ram[102] : 
                                (N26)? ram[176] : 
                                (N28)? ram[250] : 
                                (N23)? ram[324] : 
                                (N25)? ram[398] : 
                                (N27)? ram[472] : 
                                (N29)? ram[546] : 1'b0;
  assign io_deq_bits_data[19] = (N22)? ram[27] : 
                                (N24)? ram[101] : 
                                (N26)? ram[175] : 
                                (N28)? ram[249] : 
                                (N23)? ram[323] : 
                                (N25)? ram[397] : 
                                (N27)? ram[471] : 
                                (N29)? ram[545] : 1'b0;
  assign io_deq_bits_data[18] = (N22)? ram[26] : 
                                (N24)? ram[100] : 
                                (N26)? ram[174] : 
                                (N28)? ram[248] : 
                                (N23)? ram[322] : 
                                (N25)? ram[396] : 
                                (N27)? ram[470] : 
                                (N29)? ram[544] : 1'b0;
  assign io_deq_bits_data[17] = (N22)? ram[25] : 
                                (N24)? ram[99] : 
                                (N26)? ram[173] : 
                                (N28)? ram[247] : 
                                (N23)? ram[321] : 
                                (N25)? ram[395] : 
                                (N27)? ram[469] : 
                                (N29)? ram[543] : 1'b0;
  assign io_deq_bits_data[16] = (N22)? ram[24] : 
                                (N24)? ram[98] : 
                                (N26)? ram[172] : 
                                (N28)? ram[246] : 
                                (N23)? ram[320] : 
                                (N25)? ram[394] : 
                                (N27)? ram[468] : 
                                (N29)? ram[542] : 1'b0;
  assign io_deq_bits_data[15] = (N22)? ram[23] : 
                                (N24)? ram[97] : 
                                (N26)? ram[171] : 
                                (N28)? ram[245] : 
                                (N23)? ram[319] : 
                                (N25)? ram[393] : 
                                (N27)? ram[467] : 
                                (N29)? ram[541] : 1'b0;
  assign io_deq_bits_data[14] = (N22)? ram[22] : 
                                (N24)? ram[96] : 
                                (N26)? ram[170] : 
                                (N28)? ram[244] : 
                                (N23)? ram[318] : 
                                (N25)? ram[392] : 
                                (N27)? ram[466] : 
                                (N29)? ram[540] : 1'b0;
  assign io_deq_bits_data[13] = (N22)? ram[21] : 
                                (N24)? ram[95] : 
                                (N26)? ram[169] : 
                                (N28)? ram[243] : 
                                (N23)? ram[317] : 
                                (N25)? ram[391] : 
                                (N27)? ram[465] : 
                                (N29)? ram[539] : 1'b0;
  assign io_deq_bits_data[12] = (N22)? ram[20] : 
                                (N24)? ram[94] : 
                                (N26)? ram[168] : 
                                (N28)? ram[242] : 
                                (N23)? ram[316] : 
                                (N25)? ram[390] : 
                                (N27)? ram[464] : 
                                (N29)? ram[538] : 1'b0;
  assign io_deq_bits_data[11] = (N22)? ram[19] : 
                                (N24)? ram[93] : 
                                (N26)? ram[167] : 
                                (N28)? ram[241] : 
                                (N23)? ram[315] : 
                                (N25)? ram[389] : 
                                (N27)? ram[463] : 
                                (N29)? ram[537] : 1'b0;
  assign io_deq_bits_data[10] = (N22)? ram[18] : 
                                (N24)? ram[92] : 
                                (N26)? ram[166] : 
                                (N28)? ram[240] : 
                                (N23)? ram[314] : 
                                (N25)? ram[388] : 
                                (N27)? ram[462] : 
                                (N29)? ram[536] : 1'b0;
  assign io_deq_bits_data[9] = (N22)? ram[17] : 
                               (N24)? ram[91] : 
                               (N26)? ram[165] : 
                               (N28)? ram[239] : 
                               (N23)? ram[313] : 
                               (N25)? ram[387] : 
                               (N27)? ram[461] : 
                               (N29)? ram[535] : 1'b0;
  assign io_deq_bits_data[8] = (N22)? ram[16] : 
                               (N24)? ram[90] : 
                               (N26)? ram[164] : 
                               (N28)? ram[238] : 
                               (N23)? ram[312] : 
                               (N25)? ram[386] : 
                               (N27)? ram[460] : 
                               (N29)? ram[534] : 1'b0;
  assign io_deq_bits_data[7] = (N22)? ram[15] : 
                               (N24)? ram[89] : 
                               (N26)? ram[163] : 
                               (N28)? ram[237] : 
                               (N23)? ram[311] : 
                               (N25)? ram[385] : 
                               (N27)? ram[459] : 
                               (N29)? ram[533] : 1'b0;
  assign io_deq_bits_data[6] = (N22)? ram[14] : 
                               (N24)? ram[88] : 
                               (N26)? ram[162] : 
                               (N28)? ram[236] : 
                               (N23)? ram[310] : 
                               (N25)? ram[384] : 
                               (N27)? ram[458] : 
                               (N29)? ram[532] : 1'b0;
  assign io_deq_bits_data[5] = (N22)? ram[13] : 
                               (N24)? ram[87] : 
                               (N26)? ram[161] : 
                               (N28)? ram[235] : 
                               (N23)? ram[309] : 
                               (N25)? ram[383] : 
                               (N27)? ram[457] : 
                               (N29)? ram[531] : 1'b0;
  assign io_deq_bits_data[4] = (N22)? ram[12] : 
                               (N24)? ram[86] : 
                               (N26)? ram[160] : 
                               (N28)? ram[234] : 
                               (N23)? ram[308] : 
                               (N25)? ram[382] : 
                               (N27)? ram[456] : 
                               (N29)? ram[530] : 1'b0;
  assign io_deq_bits_data[3] = (N22)? ram[11] : 
                               (N24)? ram[85] : 
                               (N26)? ram[159] : 
                               (N28)? ram[233] : 
                               (N23)? ram[307] : 
                               (N25)? ram[381] : 
                               (N27)? ram[455] : 
                               (N29)? ram[529] : 1'b0;
  assign io_deq_bits_data[2] = (N22)? ram[10] : 
                               (N24)? ram[84] : 
                               (N26)? ram[158] : 
                               (N28)? ram[232] : 
                               (N23)? ram[306] : 
                               (N25)? ram[380] : 
                               (N27)? ram[454] : 
                               (N29)? ram[528] : 1'b0;
  assign io_deq_bits_data[1] = (N22)? ram[9] : 
                               (N24)? ram[83] : 
                               (N26)? ram[157] : 
                               (N28)? ram[231] : 
                               (N23)? ram[305] : 
                               (N25)? ram[379] : 
                               (N27)? ram[453] : 
                               (N29)? ram[527] : 1'b0;
  assign io_deq_bits_data[0] = (N22)? ram[8] : 
                               (N24)? ram[82] : 
                               (N26)? ram[156] : 
                               (N28)? ram[230] : 
                               (N23)? ram[304] : 
                               (N25)? ram[378] : 
                               (N27)? ram[452] : 
                               (N29)? ram[526] : 1'b0;
  assign io_deq_bits_last = (N22)? ram[7] : 
                            (N24)? ram[81] : 
                            (N26)? ram[155] : 
                            (N28)? ram[229] : 
                            (N23)? ram[303] : 
                            (N25)? ram[377] : 
                            (N27)? ram[451] : 
                            (N29)? ram[525] : 1'b0;
  assign io_deq_bits_id[5] = (N22)? ram[6] : 
                             (N24)? ram[80] : 
                             (N26)? ram[154] : 
                             (N28)? ram[228] : 
                             (N23)? ram[302] : 
                             (N25)? ram[376] : 
                             (N27)? ram[450] : 
                             (N29)? ram[524] : 1'b0;
  assign io_deq_bits_id[4] = (N22)? ram[5] : 
                             (N24)? ram[79] : 
                             (N26)? ram[153] : 
                             (N28)? ram[227] : 
                             (N23)? ram[301] : 
                             (N25)? ram[375] : 
                             (N27)? ram[449] : 
                             (N29)? ram[523] : 1'b0;
  assign io_deq_bits_id[3] = (N22)? ram[4] : 
                             (N24)? ram[78] : 
                             (N26)? ram[152] : 
                             (N28)? ram[226] : 
                             (N23)? ram[300] : 
                             (N25)? ram[374] : 
                             (N27)? ram[448] : 
                             (N29)? ram[522] : 1'b0;
  assign io_deq_bits_id[2] = (N22)? ram[3] : 
                             (N24)? ram[77] : 
                             (N26)? ram[151] : 
                             (N28)? ram[225] : 
                             (N23)? ram[299] : 
                             (N25)? ram[373] : 
                             (N27)? ram[447] : 
                             (N29)? ram[521] : 1'b0;
  assign io_deq_bits_id[1] = (N22)? ram[2] : 
                             (N24)? ram[76] : 
                             (N26)? ram[150] : 
                             (N28)? ram[224] : 
                             (N23)? ram[298] : 
                             (N25)? ram[372] : 
                             (N27)? ram[446] : 
                             (N29)? ram[520] : 1'b0;
  assign io_deq_bits_id[0] = (N22)? ram[1] : 
                             (N24)? ram[75] : 
                             (N26)? ram[149] : 
                             (N28)? ram[223] : 
                             (N23)? ram[297] : 
                             (N25)? ram[371] : 
                             (N27)? ram[445] : 
                             (N29)? ram[519] : 1'b0;
  assign io_deq_bits_user = (N22)? ram[0] : 
                            (N24)? ram[74] : 
                            (N26)? ram[148] : 
                            (N28)? ram[222] : 
                            (N23)? ram[296] : 
                            (N25)? ram[370] : 
                            (N27)? ram[444] : 
                            (N29)? ram[518] : 1'b0;

  always @(posedge clk) begin
    if(N32) begin
      R1[2] <= N35;
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      R1[1] <= N34;
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      R1[0] <= N33;
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      R4[2] <= N41;
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      R4[1] <= N40;
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      R4[0] <= N39;
    end 
  end


  always @(posedge clk) begin
    if(N44) begin
      maybe_full <= N45;
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[591] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[590] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[589] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[588] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[587] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[586] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[585] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[584] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[583] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[582] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[581] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[580] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[579] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[578] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[577] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[576] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[575] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[574] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[573] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[572] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[571] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[570] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[569] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[568] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[567] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[566] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[565] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[564] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[563] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[562] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[561] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[560] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[559] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[558] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[557] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[556] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[555] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[554] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[553] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[552] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[551] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[550] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[549] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[548] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[547] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[546] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[545] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[544] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[543] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[542] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[541] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[540] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[539] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[538] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[537] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[536] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[535] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[534] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[533] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[532] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[531] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[530] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[529] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[528] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[527] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[526] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[525] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[524] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[523] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[522] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[521] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[520] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[519] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N62) begin
      ram[518] <= io_enq_bits_user;
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[517] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[516] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[515] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[514] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[513] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[512] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[511] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[510] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[509] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[508] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[507] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[506] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[505] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[504] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[503] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[502] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[501] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[500] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[499] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[498] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[497] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[496] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[495] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[494] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[493] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[492] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[491] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[490] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[489] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[488] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[487] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[486] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[485] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[484] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[483] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[482] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[481] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[480] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[479] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[478] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[477] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[476] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[475] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[474] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[473] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[472] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[471] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[470] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[469] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[468] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[467] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[466] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[465] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[464] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[463] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[462] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[461] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[460] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[459] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[458] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[457] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[456] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[455] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[454] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[453] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[452] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[451] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[450] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[449] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[448] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[447] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[446] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[445] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N61) begin
      ram[444] <= io_enq_bits_user;
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[443] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[442] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[441] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[440] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[439] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[438] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[437] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[436] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[435] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[434] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[433] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[432] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[431] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[430] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[429] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[428] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[427] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[426] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[425] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[424] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[423] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[422] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[421] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[420] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[419] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[418] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[417] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[416] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[415] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[414] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[413] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[412] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[411] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[410] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[409] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[408] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[407] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[406] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[405] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[404] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[403] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[402] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[401] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[400] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[399] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[398] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[397] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[396] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[395] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[394] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[393] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[392] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[391] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[390] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[389] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[388] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[387] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[386] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[385] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[384] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[383] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[382] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[381] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[380] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[379] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[378] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[377] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[376] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[375] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[374] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[373] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[372] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[371] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N60) begin
      ram[370] <= io_enq_bits_user;
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[369] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[368] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[367] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[366] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[365] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[364] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[363] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[362] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[361] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[360] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[359] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[358] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[357] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[356] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[355] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[354] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[353] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[352] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[351] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[350] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[349] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[348] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[347] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[346] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[345] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[344] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[343] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[342] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[341] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[340] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[339] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[338] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[337] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[336] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[335] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[334] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[333] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[332] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[331] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[330] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[329] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[328] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[327] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[326] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[325] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[324] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[323] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[322] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[321] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[320] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[319] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[318] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[317] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[316] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[315] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[314] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[313] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[312] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[311] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[310] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[309] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[308] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[307] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[306] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[305] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[304] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[303] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[302] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[301] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[300] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[299] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[298] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[297] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      ram[296] <= io_enq_bits_user;
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[295] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[294] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[293] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[292] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[291] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[290] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[289] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[288] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[287] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[286] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[285] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[284] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[283] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[282] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[281] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[280] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[279] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[278] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[277] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[276] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[275] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[274] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[273] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[272] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[271] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[270] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[269] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[268] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[267] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[266] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[265] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[264] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[263] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[262] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[261] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[260] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[259] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[258] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[257] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[256] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[255] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[254] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[253] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[252] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[251] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[250] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[249] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[248] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[247] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[246] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[245] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[244] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[243] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[242] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[241] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[240] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[239] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[238] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[237] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[236] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[235] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[234] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[233] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[232] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[231] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[230] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[229] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[228] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[227] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[226] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[225] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[224] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[223] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N58) begin
      ram[222] <= io_enq_bits_user;
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[221] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[220] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[219] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[218] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[217] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[216] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[215] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[214] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[213] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[212] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[211] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[210] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[209] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[208] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[207] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[206] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[205] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[204] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[203] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[202] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[201] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[200] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[199] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[198] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[197] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[196] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[195] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[194] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[193] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[192] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[191] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[190] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[189] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[188] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[187] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[186] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[185] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[184] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[183] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[182] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[181] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[180] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[179] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[178] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[177] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[176] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[175] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[174] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[173] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[172] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[171] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[170] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[169] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[168] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[167] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[166] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[165] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[164] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[163] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[162] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[161] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[160] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[159] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[158] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[157] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[156] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[155] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[154] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[153] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[152] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[151] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[150] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[149] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N57) begin
      ram[148] <= io_enq_bits_user;
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[147] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[146] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[145] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[144] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[143] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[142] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[141] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[140] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[139] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[138] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[137] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[136] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[135] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[134] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[133] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[132] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[131] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[130] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[129] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[128] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[127] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[126] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[125] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[124] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[123] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[122] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[121] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[120] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[119] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[118] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[117] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[116] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[115] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[114] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[113] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[112] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[111] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[110] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[109] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[108] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[107] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[106] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[105] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[104] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[103] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[102] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[101] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[100] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[99] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[98] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[97] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[96] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[95] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[94] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[93] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[92] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[91] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[90] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[89] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[88] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[87] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[86] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[85] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[84] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[83] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[82] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[81] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[80] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[79] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[78] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[77] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[76] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[75] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N56) begin
      ram[74] <= io_enq_bits_user;
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[73] <= io_enq_bits_resp[1];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[72] <= io_enq_bits_resp[0];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[71] <= io_enq_bits_data[63];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[70] <= io_enq_bits_data[62];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[69] <= io_enq_bits_data[61];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[68] <= io_enq_bits_data[60];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[67] <= io_enq_bits_data[59];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[66] <= io_enq_bits_data[58];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[65] <= io_enq_bits_data[57];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[64] <= io_enq_bits_data[56];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[63] <= io_enq_bits_data[55];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[62] <= io_enq_bits_data[54];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[61] <= io_enq_bits_data[53];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[60] <= io_enq_bits_data[52];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[59] <= io_enq_bits_data[51];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[58] <= io_enq_bits_data[50];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[57] <= io_enq_bits_data[49];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[56] <= io_enq_bits_data[48];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[55] <= io_enq_bits_data[47];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[54] <= io_enq_bits_data[46];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[53] <= io_enq_bits_data[45];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[52] <= io_enq_bits_data[44];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[51] <= io_enq_bits_data[43];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[50] <= io_enq_bits_data[42];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[49] <= io_enq_bits_data[41];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[48] <= io_enq_bits_data[40];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[47] <= io_enq_bits_data[39];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[46] <= io_enq_bits_data[38];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[45] <= io_enq_bits_data[37];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[44] <= io_enq_bits_data[36];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[43] <= io_enq_bits_data[35];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[42] <= io_enq_bits_data[34];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[41] <= io_enq_bits_data[33];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[40] <= io_enq_bits_data[32];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[39] <= io_enq_bits_data[31];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[38] <= io_enq_bits_data[30];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[37] <= io_enq_bits_data[29];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[36] <= io_enq_bits_data[28];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[35] <= io_enq_bits_data[27];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[34] <= io_enq_bits_data[26];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[33] <= io_enq_bits_data[25];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[32] <= io_enq_bits_data[24];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[31] <= io_enq_bits_data[23];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[30] <= io_enq_bits_data[22];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[29] <= io_enq_bits_data[21];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[28] <= io_enq_bits_data[20];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[27] <= io_enq_bits_data[19];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[26] <= io_enq_bits_data[18];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[25] <= io_enq_bits_data[17];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[24] <= io_enq_bits_data[16];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[23] <= io_enq_bits_data[15];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[22] <= io_enq_bits_data[14];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[21] <= io_enq_bits_data[13];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[20] <= io_enq_bits_data[12];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[19] <= io_enq_bits_data[11];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[18] <= io_enq_bits_data[10];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[17] <= io_enq_bits_data[9];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[16] <= io_enq_bits_data[8];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[15] <= io_enq_bits_data[7];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[14] <= io_enq_bits_data[6];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[13] <= io_enq_bits_data[5];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[12] <= io_enq_bits_data[4];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[11] <= io_enq_bits_data[3];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[10] <= io_enq_bits_data[2];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[9] <= io_enq_bits_data[1];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[8] <= io_enq_bits_data[0];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[7] <= io_enq_bits_last;
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[6] <= io_enq_bits_id[5];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[5] <= io_enq_bits_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[4] <= io_enq_bits_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[3] <= io_enq_bits_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[2] <= io_enq_bits_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[1] <= io_enq_bits_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N55) begin
      ram[0] <= io_enq_bits_user;
    end 
  end

  assign io_count[2:0] = R4 - R1;
  assign T3 = R1 + 1'b1;
  assign T6 = R4 + 1'b1;
  assign N67 = R4[0] & R4[1];
  assign N54 = N67 & R4[2];
  assign N68 = N0 & R4[1];
  assign N0 = ~R4[0];
  assign N53 = N68 & R4[2];
  assign N69 = R4[0] & N1;
  assign N1 = ~R4[1];
  assign N52 = N69 & R4[2];
  assign N70 = N2 & N3;
  assign N2 = ~R4[0];
  assign N3 = ~R4[1];
  assign N51 = N70 & R4[2];
  assign N71 = R4[0] & R4[1];
  assign N50 = N71 & N4;
  assign N4 = ~R4[2];
  assign N72 = N5 & R4[1];
  assign N5 = ~R4[0];
  assign N49 = N72 & N6;
  assign N6 = ~R4[2];
  assign N73 = R4[0] & N7;
  assign N7 = ~R4[1];
  assign N48 = N73 & N8;
  assign N8 = ~R4[2];
  assign N74 = N9 & N10;
  assign N9 = ~R4[0];
  assign N10 = ~R4[1];
  assign N47 = N74 & N11;
  assign N11 = ~R4[2];
  assign N32 = (N12)? 1'b1 : 
               (N64)? 1'b1 : 
               (N31)? 1'b0 : 1'b0;
  assign N12 = reset;
  assign { N35, N34, N33 } = (N12)? { 1'b0, 1'b0, 1'b0 } : 
                             (N64)? T3 : 1'b0;
  assign N38 = (N12)? 1'b1 : 
               (N65)? 1'b1 : 
               (N37)? 1'b0 : 1'b0;
  assign { N41, N40, N39 } = (N12)? { 1'b0, 1'b0, 1'b0 } : 
                             (N65)? T6 : 1'b0;
  assign N44 = (N12)? 1'b1 : 
               (N66)? 1'b1 : 
               (N43)? 1'b0 : 1'b0;
  assign N45 = (N12)? 1'b0 : 
               (N66)? do_enq : 1'b0;
  assign { N62, N61, N60, N59, N58, N57, N56, N55 } = (N13)? { N54, N53, N52, N51, N50, N49, N48, N47 } : 
                                                      (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = do_enq;
  assign N14 = N46;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_count[3] = maybe_full & ptr_match;
  assign N15 = ~R1[0];
  assign N16 = ~R1[1];
  assign N17 = N15 & N16;
  assign N18 = N15 & R1[1];
  assign N19 = R1[0] & N16;
  assign N20 = R1[0] & R1[1];
  assign N21 = ~R1[2];
  assign N22 = N17 & N21;
  assign N23 = N17 & R1[2];
  assign N24 = N19 & N21;
  assign N25 = N19 & R1[2];
  assign N26 = N18 & N21;
  assign N27 = N18 & R1[2];
  assign N28 = N20 & N21;
  assign N29 = N20 & R1[2];
  assign io_deq_valid = ~empty;
  assign empty = ptr_match & T23;
  assign T23 = ~maybe_full;
  assign io_enq_ready = ~full;
  assign full = ptr_match & maybe_full;
  assign N30 = do_deq | reset;
  assign N31 = ~N30;
  assign N36 = do_enq | reset;
  assign N37 = ~N36;
  assign N42 = T9 | reset;
  assign N43 = ~N42;
  assign N46 = ~do_enq;
  assign N63 = ~reset;
  assign N64 = do_deq & N63;
  assign N65 = do_enq & N63;
  assign N66 = T9 & N63;

endmodule