module bsg_mem_1r1w_synth_width_p572_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [571:0] w_data_i;
  input [0:0] r_addr_i;
  output [571:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [571:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  wire [1143:0] mem;
  reg mem_1143_sv2v_reg,mem_1142_sv2v_reg,mem_1141_sv2v_reg,mem_1140_sv2v_reg,
  mem_1139_sv2v_reg,mem_1138_sv2v_reg,mem_1137_sv2v_reg,mem_1136_sv2v_reg,
  mem_1135_sv2v_reg,mem_1134_sv2v_reg,mem_1133_sv2v_reg,mem_1132_sv2v_reg,mem_1131_sv2v_reg,
  mem_1130_sv2v_reg,mem_1129_sv2v_reg,mem_1128_sv2v_reg,mem_1127_sv2v_reg,
  mem_1126_sv2v_reg,mem_1125_sv2v_reg,mem_1124_sv2v_reg,mem_1123_sv2v_reg,mem_1122_sv2v_reg,
  mem_1121_sv2v_reg,mem_1120_sv2v_reg,mem_1119_sv2v_reg,mem_1118_sv2v_reg,
  mem_1117_sv2v_reg,mem_1116_sv2v_reg,mem_1115_sv2v_reg,mem_1114_sv2v_reg,mem_1113_sv2v_reg,
  mem_1112_sv2v_reg,mem_1111_sv2v_reg,mem_1110_sv2v_reg,mem_1109_sv2v_reg,
  mem_1108_sv2v_reg,mem_1107_sv2v_reg,mem_1106_sv2v_reg,mem_1105_sv2v_reg,mem_1104_sv2v_reg,
  mem_1103_sv2v_reg,mem_1102_sv2v_reg,mem_1101_sv2v_reg,mem_1100_sv2v_reg,
  mem_1099_sv2v_reg,mem_1098_sv2v_reg,mem_1097_sv2v_reg,mem_1096_sv2v_reg,
  mem_1095_sv2v_reg,mem_1094_sv2v_reg,mem_1093_sv2v_reg,mem_1092_sv2v_reg,mem_1091_sv2v_reg,
  mem_1090_sv2v_reg,mem_1089_sv2v_reg,mem_1088_sv2v_reg,mem_1087_sv2v_reg,
  mem_1086_sv2v_reg,mem_1085_sv2v_reg,mem_1084_sv2v_reg,mem_1083_sv2v_reg,mem_1082_sv2v_reg,
  mem_1081_sv2v_reg,mem_1080_sv2v_reg,mem_1079_sv2v_reg,mem_1078_sv2v_reg,
  mem_1077_sv2v_reg,mem_1076_sv2v_reg,mem_1075_sv2v_reg,mem_1074_sv2v_reg,mem_1073_sv2v_reg,
  mem_1072_sv2v_reg,mem_1071_sv2v_reg,mem_1070_sv2v_reg,mem_1069_sv2v_reg,
  mem_1068_sv2v_reg,mem_1067_sv2v_reg,mem_1066_sv2v_reg,mem_1065_sv2v_reg,mem_1064_sv2v_reg,
  mem_1063_sv2v_reg,mem_1062_sv2v_reg,mem_1061_sv2v_reg,mem_1060_sv2v_reg,
  mem_1059_sv2v_reg,mem_1058_sv2v_reg,mem_1057_sv2v_reg,mem_1056_sv2v_reg,
  mem_1055_sv2v_reg,mem_1054_sv2v_reg,mem_1053_sv2v_reg,mem_1052_sv2v_reg,mem_1051_sv2v_reg,
  mem_1050_sv2v_reg,mem_1049_sv2v_reg,mem_1048_sv2v_reg,mem_1047_sv2v_reg,
  mem_1046_sv2v_reg,mem_1045_sv2v_reg,mem_1044_sv2v_reg,mem_1043_sv2v_reg,mem_1042_sv2v_reg,
  mem_1041_sv2v_reg,mem_1040_sv2v_reg,mem_1039_sv2v_reg,mem_1038_sv2v_reg,
  mem_1037_sv2v_reg,mem_1036_sv2v_reg,mem_1035_sv2v_reg,mem_1034_sv2v_reg,mem_1033_sv2v_reg,
  mem_1032_sv2v_reg,mem_1031_sv2v_reg,mem_1030_sv2v_reg,mem_1029_sv2v_reg,
  mem_1028_sv2v_reg,mem_1027_sv2v_reg,mem_1026_sv2v_reg,mem_1025_sv2v_reg,mem_1024_sv2v_reg,
  mem_1023_sv2v_reg,mem_1022_sv2v_reg,mem_1021_sv2v_reg,mem_1020_sv2v_reg,
  mem_1019_sv2v_reg,mem_1018_sv2v_reg,mem_1017_sv2v_reg,mem_1016_sv2v_reg,
  mem_1015_sv2v_reg,mem_1014_sv2v_reg,mem_1013_sv2v_reg,mem_1012_sv2v_reg,mem_1011_sv2v_reg,
  mem_1010_sv2v_reg,mem_1009_sv2v_reg,mem_1008_sv2v_reg,mem_1007_sv2v_reg,
  mem_1006_sv2v_reg,mem_1005_sv2v_reg,mem_1004_sv2v_reg,mem_1003_sv2v_reg,mem_1002_sv2v_reg,
  mem_1001_sv2v_reg,mem_1000_sv2v_reg,mem_999_sv2v_reg,mem_998_sv2v_reg,
  mem_997_sv2v_reg,mem_996_sv2v_reg,mem_995_sv2v_reg,mem_994_sv2v_reg,mem_993_sv2v_reg,
  mem_992_sv2v_reg,mem_991_sv2v_reg,mem_990_sv2v_reg,mem_989_sv2v_reg,mem_988_sv2v_reg,
  mem_987_sv2v_reg,mem_986_sv2v_reg,mem_985_sv2v_reg,mem_984_sv2v_reg,
  mem_983_sv2v_reg,mem_982_sv2v_reg,mem_981_sv2v_reg,mem_980_sv2v_reg,mem_979_sv2v_reg,
  mem_978_sv2v_reg,mem_977_sv2v_reg,mem_976_sv2v_reg,mem_975_sv2v_reg,mem_974_sv2v_reg,
  mem_973_sv2v_reg,mem_972_sv2v_reg,mem_971_sv2v_reg,mem_970_sv2v_reg,mem_969_sv2v_reg,
  mem_968_sv2v_reg,mem_967_sv2v_reg,mem_966_sv2v_reg,mem_965_sv2v_reg,
  mem_964_sv2v_reg,mem_963_sv2v_reg,mem_962_sv2v_reg,mem_961_sv2v_reg,mem_960_sv2v_reg,
  mem_959_sv2v_reg,mem_958_sv2v_reg,mem_957_sv2v_reg,mem_956_sv2v_reg,mem_955_sv2v_reg,
  mem_954_sv2v_reg,mem_953_sv2v_reg,mem_952_sv2v_reg,mem_951_sv2v_reg,
  mem_950_sv2v_reg,mem_949_sv2v_reg,mem_948_sv2v_reg,mem_947_sv2v_reg,mem_946_sv2v_reg,
  mem_945_sv2v_reg,mem_944_sv2v_reg,mem_943_sv2v_reg,mem_942_sv2v_reg,mem_941_sv2v_reg,
  mem_940_sv2v_reg,mem_939_sv2v_reg,mem_938_sv2v_reg,mem_937_sv2v_reg,mem_936_sv2v_reg,
  mem_935_sv2v_reg,mem_934_sv2v_reg,mem_933_sv2v_reg,mem_932_sv2v_reg,
  mem_931_sv2v_reg,mem_930_sv2v_reg,mem_929_sv2v_reg,mem_928_sv2v_reg,mem_927_sv2v_reg,
  mem_926_sv2v_reg,mem_925_sv2v_reg,mem_924_sv2v_reg,mem_923_sv2v_reg,mem_922_sv2v_reg,
  mem_921_sv2v_reg,mem_920_sv2v_reg,mem_919_sv2v_reg,mem_918_sv2v_reg,
  mem_917_sv2v_reg,mem_916_sv2v_reg,mem_915_sv2v_reg,mem_914_sv2v_reg,mem_913_sv2v_reg,
  mem_912_sv2v_reg,mem_911_sv2v_reg,mem_910_sv2v_reg,mem_909_sv2v_reg,mem_908_sv2v_reg,
  mem_907_sv2v_reg,mem_906_sv2v_reg,mem_905_sv2v_reg,mem_904_sv2v_reg,
  mem_903_sv2v_reg,mem_902_sv2v_reg,mem_901_sv2v_reg,mem_900_sv2v_reg,mem_899_sv2v_reg,
  mem_898_sv2v_reg,mem_897_sv2v_reg,mem_896_sv2v_reg,mem_895_sv2v_reg,mem_894_sv2v_reg,
  mem_893_sv2v_reg,mem_892_sv2v_reg,mem_891_sv2v_reg,mem_890_sv2v_reg,mem_889_sv2v_reg,
  mem_888_sv2v_reg,mem_887_sv2v_reg,mem_886_sv2v_reg,mem_885_sv2v_reg,
  mem_884_sv2v_reg,mem_883_sv2v_reg,mem_882_sv2v_reg,mem_881_sv2v_reg,mem_880_sv2v_reg,
  mem_879_sv2v_reg,mem_878_sv2v_reg,mem_877_sv2v_reg,mem_876_sv2v_reg,mem_875_sv2v_reg,
  mem_874_sv2v_reg,mem_873_sv2v_reg,mem_872_sv2v_reg,mem_871_sv2v_reg,
  mem_870_sv2v_reg,mem_869_sv2v_reg,mem_868_sv2v_reg,mem_867_sv2v_reg,mem_866_sv2v_reg,
  mem_865_sv2v_reg,mem_864_sv2v_reg,mem_863_sv2v_reg,mem_862_sv2v_reg,mem_861_sv2v_reg,
  mem_860_sv2v_reg,mem_859_sv2v_reg,mem_858_sv2v_reg,mem_857_sv2v_reg,mem_856_sv2v_reg,
  mem_855_sv2v_reg,mem_854_sv2v_reg,mem_853_sv2v_reg,mem_852_sv2v_reg,
  mem_851_sv2v_reg,mem_850_sv2v_reg,mem_849_sv2v_reg,mem_848_sv2v_reg,mem_847_sv2v_reg,
  mem_846_sv2v_reg,mem_845_sv2v_reg,mem_844_sv2v_reg,mem_843_sv2v_reg,mem_842_sv2v_reg,
  mem_841_sv2v_reg,mem_840_sv2v_reg,mem_839_sv2v_reg,mem_838_sv2v_reg,
  mem_837_sv2v_reg,mem_836_sv2v_reg,mem_835_sv2v_reg,mem_834_sv2v_reg,mem_833_sv2v_reg,
  mem_832_sv2v_reg,mem_831_sv2v_reg,mem_830_sv2v_reg,mem_829_sv2v_reg,mem_828_sv2v_reg,
  mem_827_sv2v_reg,mem_826_sv2v_reg,mem_825_sv2v_reg,mem_824_sv2v_reg,
  mem_823_sv2v_reg,mem_822_sv2v_reg,mem_821_sv2v_reg,mem_820_sv2v_reg,mem_819_sv2v_reg,
  mem_818_sv2v_reg,mem_817_sv2v_reg,mem_816_sv2v_reg,mem_815_sv2v_reg,mem_814_sv2v_reg,
  mem_813_sv2v_reg,mem_812_sv2v_reg,mem_811_sv2v_reg,mem_810_sv2v_reg,mem_809_sv2v_reg,
  mem_808_sv2v_reg,mem_807_sv2v_reg,mem_806_sv2v_reg,mem_805_sv2v_reg,
  mem_804_sv2v_reg,mem_803_sv2v_reg,mem_802_sv2v_reg,mem_801_sv2v_reg,mem_800_sv2v_reg,
  mem_799_sv2v_reg,mem_798_sv2v_reg,mem_797_sv2v_reg,mem_796_sv2v_reg,mem_795_sv2v_reg,
  mem_794_sv2v_reg,mem_793_sv2v_reg,mem_792_sv2v_reg,mem_791_sv2v_reg,
  mem_790_sv2v_reg,mem_789_sv2v_reg,mem_788_sv2v_reg,mem_787_sv2v_reg,mem_786_sv2v_reg,
  mem_785_sv2v_reg,mem_784_sv2v_reg,mem_783_sv2v_reg,mem_782_sv2v_reg,mem_781_sv2v_reg,
  mem_780_sv2v_reg,mem_779_sv2v_reg,mem_778_sv2v_reg,mem_777_sv2v_reg,mem_776_sv2v_reg,
  mem_775_sv2v_reg,mem_774_sv2v_reg,mem_773_sv2v_reg,mem_772_sv2v_reg,
  mem_771_sv2v_reg,mem_770_sv2v_reg,mem_769_sv2v_reg,mem_768_sv2v_reg,mem_767_sv2v_reg,
  mem_766_sv2v_reg,mem_765_sv2v_reg,mem_764_sv2v_reg,mem_763_sv2v_reg,mem_762_sv2v_reg,
  mem_761_sv2v_reg,mem_760_sv2v_reg,mem_759_sv2v_reg,mem_758_sv2v_reg,
  mem_757_sv2v_reg,mem_756_sv2v_reg,mem_755_sv2v_reg,mem_754_sv2v_reg,mem_753_sv2v_reg,
  mem_752_sv2v_reg,mem_751_sv2v_reg,mem_750_sv2v_reg,mem_749_sv2v_reg,mem_748_sv2v_reg,
  mem_747_sv2v_reg,mem_746_sv2v_reg,mem_745_sv2v_reg,mem_744_sv2v_reg,
  mem_743_sv2v_reg,mem_742_sv2v_reg,mem_741_sv2v_reg,mem_740_sv2v_reg,mem_739_sv2v_reg,
  mem_738_sv2v_reg,mem_737_sv2v_reg,mem_736_sv2v_reg,mem_735_sv2v_reg,mem_734_sv2v_reg,
  mem_733_sv2v_reg,mem_732_sv2v_reg,mem_731_sv2v_reg,mem_730_sv2v_reg,mem_729_sv2v_reg,
  mem_728_sv2v_reg,mem_727_sv2v_reg,mem_726_sv2v_reg,mem_725_sv2v_reg,
  mem_724_sv2v_reg,mem_723_sv2v_reg,mem_722_sv2v_reg,mem_721_sv2v_reg,mem_720_sv2v_reg,
  mem_719_sv2v_reg,mem_718_sv2v_reg,mem_717_sv2v_reg,mem_716_sv2v_reg,mem_715_sv2v_reg,
  mem_714_sv2v_reg,mem_713_sv2v_reg,mem_712_sv2v_reg,mem_711_sv2v_reg,
  mem_710_sv2v_reg,mem_709_sv2v_reg,mem_708_sv2v_reg,mem_707_sv2v_reg,mem_706_sv2v_reg,
  mem_705_sv2v_reg,mem_704_sv2v_reg,mem_703_sv2v_reg,mem_702_sv2v_reg,mem_701_sv2v_reg,
  mem_700_sv2v_reg,mem_699_sv2v_reg,mem_698_sv2v_reg,mem_697_sv2v_reg,mem_696_sv2v_reg,
  mem_695_sv2v_reg,mem_694_sv2v_reg,mem_693_sv2v_reg,mem_692_sv2v_reg,
  mem_691_sv2v_reg,mem_690_sv2v_reg,mem_689_sv2v_reg,mem_688_sv2v_reg,mem_687_sv2v_reg,
  mem_686_sv2v_reg,mem_685_sv2v_reg,mem_684_sv2v_reg,mem_683_sv2v_reg,mem_682_sv2v_reg,
  mem_681_sv2v_reg,mem_680_sv2v_reg,mem_679_sv2v_reg,mem_678_sv2v_reg,
  mem_677_sv2v_reg,mem_676_sv2v_reg,mem_675_sv2v_reg,mem_674_sv2v_reg,mem_673_sv2v_reg,
  mem_672_sv2v_reg,mem_671_sv2v_reg,mem_670_sv2v_reg,mem_669_sv2v_reg,mem_668_sv2v_reg,
  mem_667_sv2v_reg,mem_666_sv2v_reg,mem_665_sv2v_reg,mem_664_sv2v_reg,
  mem_663_sv2v_reg,mem_662_sv2v_reg,mem_661_sv2v_reg,mem_660_sv2v_reg,mem_659_sv2v_reg,
  mem_658_sv2v_reg,mem_657_sv2v_reg,mem_656_sv2v_reg,mem_655_sv2v_reg,mem_654_sv2v_reg,
  mem_653_sv2v_reg,mem_652_sv2v_reg,mem_651_sv2v_reg,mem_650_sv2v_reg,mem_649_sv2v_reg,
  mem_648_sv2v_reg,mem_647_sv2v_reg,mem_646_sv2v_reg,mem_645_sv2v_reg,
  mem_644_sv2v_reg,mem_643_sv2v_reg,mem_642_sv2v_reg,mem_641_sv2v_reg,mem_640_sv2v_reg,
  mem_639_sv2v_reg,mem_638_sv2v_reg,mem_637_sv2v_reg,mem_636_sv2v_reg,mem_635_sv2v_reg,
  mem_634_sv2v_reg,mem_633_sv2v_reg,mem_632_sv2v_reg,mem_631_sv2v_reg,
  mem_630_sv2v_reg,mem_629_sv2v_reg,mem_628_sv2v_reg,mem_627_sv2v_reg,mem_626_sv2v_reg,
  mem_625_sv2v_reg,mem_624_sv2v_reg,mem_623_sv2v_reg,mem_622_sv2v_reg,mem_621_sv2v_reg,
  mem_620_sv2v_reg,mem_619_sv2v_reg,mem_618_sv2v_reg,mem_617_sv2v_reg,mem_616_sv2v_reg,
  mem_615_sv2v_reg,mem_614_sv2v_reg,mem_613_sv2v_reg,mem_612_sv2v_reg,
  mem_611_sv2v_reg,mem_610_sv2v_reg,mem_609_sv2v_reg,mem_608_sv2v_reg,mem_607_sv2v_reg,
  mem_606_sv2v_reg,mem_605_sv2v_reg,mem_604_sv2v_reg,mem_603_sv2v_reg,mem_602_sv2v_reg,
  mem_601_sv2v_reg,mem_600_sv2v_reg,mem_599_sv2v_reg,mem_598_sv2v_reg,
  mem_597_sv2v_reg,mem_596_sv2v_reg,mem_595_sv2v_reg,mem_594_sv2v_reg,mem_593_sv2v_reg,
  mem_592_sv2v_reg,mem_591_sv2v_reg,mem_590_sv2v_reg,mem_589_sv2v_reg,mem_588_sv2v_reg,
  mem_587_sv2v_reg,mem_586_sv2v_reg,mem_585_sv2v_reg,mem_584_sv2v_reg,
  mem_583_sv2v_reg,mem_582_sv2v_reg,mem_581_sv2v_reg,mem_580_sv2v_reg,mem_579_sv2v_reg,
  mem_578_sv2v_reg,mem_577_sv2v_reg,mem_576_sv2v_reg,mem_575_sv2v_reg,mem_574_sv2v_reg,
  mem_573_sv2v_reg,mem_572_sv2v_reg,mem_571_sv2v_reg,mem_570_sv2v_reg,mem_569_sv2v_reg,
  mem_568_sv2v_reg,mem_567_sv2v_reg,mem_566_sv2v_reg,mem_565_sv2v_reg,
  mem_564_sv2v_reg,mem_563_sv2v_reg,mem_562_sv2v_reg,mem_561_sv2v_reg,mem_560_sv2v_reg,
  mem_559_sv2v_reg,mem_558_sv2v_reg,mem_557_sv2v_reg,mem_556_sv2v_reg,mem_555_sv2v_reg,
  mem_554_sv2v_reg,mem_553_sv2v_reg,mem_552_sv2v_reg,mem_551_sv2v_reg,
  mem_550_sv2v_reg,mem_549_sv2v_reg,mem_548_sv2v_reg,mem_547_sv2v_reg,mem_546_sv2v_reg,
  mem_545_sv2v_reg,mem_544_sv2v_reg,mem_543_sv2v_reg,mem_542_sv2v_reg,mem_541_sv2v_reg,
  mem_540_sv2v_reg,mem_539_sv2v_reg,mem_538_sv2v_reg,mem_537_sv2v_reg,mem_536_sv2v_reg,
  mem_535_sv2v_reg,mem_534_sv2v_reg,mem_533_sv2v_reg,mem_532_sv2v_reg,
  mem_531_sv2v_reg,mem_530_sv2v_reg,mem_529_sv2v_reg,mem_528_sv2v_reg,mem_527_sv2v_reg,
  mem_526_sv2v_reg,mem_525_sv2v_reg,mem_524_sv2v_reg,mem_523_sv2v_reg,mem_522_sv2v_reg,
  mem_521_sv2v_reg,mem_520_sv2v_reg,mem_519_sv2v_reg,mem_518_sv2v_reg,
  mem_517_sv2v_reg,mem_516_sv2v_reg,mem_515_sv2v_reg,mem_514_sv2v_reg,mem_513_sv2v_reg,
  mem_512_sv2v_reg,mem_511_sv2v_reg,mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,
  mem_507_sv2v_reg,mem_506_sv2v_reg,mem_505_sv2v_reg,mem_504_sv2v_reg,
  mem_503_sv2v_reg,mem_502_sv2v_reg,mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,
  mem_498_sv2v_reg,mem_497_sv2v_reg,mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,
  mem_493_sv2v_reg,mem_492_sv2v_reg,mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,
  mem_488_sv2v_reg,mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,
  mem_484_sv2v_reg,mem_483_sv2v_reg,mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,
  mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,
  mem_474_sv2v_reg,mem_473_sv2v_reg,mem_472_sv2v_reg,mem_471_sv2v_reg,
  mem_470_sv2v_reg,mem_469_sv2v_reg,mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,
  mem_465_sv2v_reg,mem_464_sv2v_reg,mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,
  mem_460_sv2v_reg,mem_459_sv2v_reg,mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,
  mem_455_sv2v_reg,mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,
  mem_451_sv2v_reg,mem_450_sv2v_reg,mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,
  mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,
  mem_441_sv2v_reg,mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,
  mem_437_sv2v_reg,mem_436_sv2v_reg,mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,
  mem_432_sv2v_reg,mem_431_sv2v_reg,mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,
  mem_427_sv2v_reg,mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,
  mem_423_sv2v_reg,mem_422_sv2v_reg,mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,
  mem_418_sv2v_reg,mem_417_sv2v_reg,mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,
  mem_413_sv2v_reg,mem_412_sv2v_reg,mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,
  mem_408_sv2v_reg,mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,
  mem_404_sv2v_reg,mem_403_sv2v_reg,mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,
  mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,
  mem_394_sv2v_reg,mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,
  mem_390_sv2v_reg,mem_389_sv2v_reg,mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,
  mem_385_sv2v_reg,mem_384_sv2v_reg,mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,
  mem_380_sv2v_reg,mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,
  mem_375_sv2v_reg,mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,
  mem_371_sv2v_reg,mem_370_sv2v_reg,mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,
  mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,
  mem_361_sv2v_reg,mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,
  mem_357_sv2v_reg,mem_356_sv2v_reg,mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,
  mem_352_sv2v_reg,mem_351_sv2v_reg,mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,
  mem_347_sv2v_reg,mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,
  mem_343_sv2v_reg,mem_342_sv2v_reg,mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,
  mem_338_sv2v_reg,mem_337_sv2v_reg,mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,
  mem_333_sv2v_reg,mem_332_sv2v_reg,mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,
  mem_328_sv2v_reg,mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,
  mem_324_sv2v_reg,mem_323_sv2v_reg,mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,
  mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,
  mem_314_sv2v_reg,mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,
  mem_310_sv2v_reg,mem_309_sv2v_reg,mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,
  mem_305_sv2v_reg,mem_304_sv2v_reg,mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,
  mem_300_sv2v_reg,mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,
  mem_295_sv2v_reg,mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,
  mem_291_sv2v_reg,mem_290_sv2v_reg,mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,
  mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,
  mem_281_sv2v_reg,mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,
  mem_277_sv2v_reg,mem_276_sv2v_reg,mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,
  mem_272_sv2v_reg,mem_271_sv2v_reg,mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,
  mem_267_sv2v_reg,mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,
  mem_263_sv2v_reg,mem_262_sv2v_reg,mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,
  mem_258_sv2v_reg,mem_257_sv2v_reg,mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,
  mem_253_sv2v_reg,mem_252_sv2v_reg,mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,
  mem_248_sv2v_reg,mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,
  mem_244_sv2v_reg,mem_243_sv2v_reg,mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,
  mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,
  mem_234_sv2v_reg,mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,
  mem_230_sv2v_reg,mem_229_sv2v_reg,mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,
  mem_225_sv2v_reg,mem_224_sv2v_reg,mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,
  mem_220_sv2v_reg,mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,
  mem_215_sv2v_reg,mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,
  mem_211_sv2v_reg,mem_210_sv2v_reg,mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,
  mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,
  mem_201_sv2v_reg,mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,
  mem_197_sv2v_reg,mem_196_sv2v_reg,mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,
  mem_192_sv2v_reg,mem_191_sv2v_reg,mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,
  mem_187_sv2v_reg,mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,
  mem_183_sv2v_reg,mem_182_sv2v_reg,mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,
  mem_178_sv2v_reg,mem_177_sv2v_reg,mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,
  mem_173_sv2v_reg,mem_172_sv2v_reg,mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,
  mem_168_sv2v_reg,mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,
  mem_164_sv2v_reg,mem_163_sv2v_reg,mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,
  mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,
  mem_154_sv2v_reg,mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,
  mem_150_sv2v_reg,mem_149_sv2v_reg,mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,
  mem_145_sv2v_reg,mem_144_sv2v_reg,mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,
  mem_140_sv2v_reg,mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,
  mem_135_sv2v_reg,mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,
  mem_131_sv2v_reg,mem_130_sv2v_reg,mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,
  mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,
  mem_121_sv2v_reg,mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,
  mem_117_sv2v_reg,mem_116_sv2v_reg,mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,
  mem_112_sv2v_reg,mem_111_sv2v_reg,mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,
  mem_107_sv2v_reg,mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,
  mem_103_sv2v_reg,mem_102_sv2v_reg,mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,
  mem_98_sv2v_reg,mem_97_sv2v_reg,mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,
  mem_93_sv2v_reg,mem_92_sv2v_reg,mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,
  mem_88_sv2v_reg,mem_87_sv2v_reg,mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,
  mem_83_sv2v_reg,mem_82_sv2v_reg,mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,
  mem_78_sv2v_reg,mem_77_sv2v_reg,mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,
  mem_73_sv2v_reg,mem_72_sv2v_reg,mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,
  mem_68_sv2v_reg,mem_67_sv2v_reg,mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,
  mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,
  mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,
  mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,
  mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,
  mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,
  mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,
  mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,
  mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,
  mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,
  mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,
  mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,
  mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,
  mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[1143] = mem_1143_sv2v_reg;
  assign mem[1142] = mem_1142_sv2v_reg;
  assign mem[1141] = mem_1141_sv2v_reg;
  assign mem[1140] = mem_1140_sv2v_reg;
  assign mem[1139] = mem_1139_sv2v_reg;
  assign mem[1138] = mem_1138_sv2v_reg;
  assign mem[1137] = mem_1137_sv2v_reg;
  assign mem[1136] = mem_1136_sv2v_reg;
  assign mem[1135] = mem_1135_sv2v_reg;
  assign mem[1134] = mem_1134_sv2v_reg;
  assign mem[1133] = mem_1133_sv2v_reg;
  assign mem[1132] = mem_1132_sv2v_reg;
  assign mem[1131] = mem_1131_sv2v_reg;
  assign mem[1130] = mem_1130_sv2v_reg;
  assign mem[1129] = mem_1129_sv2v_reg;
  assign mem[1128] = mem_1128_sv2v_reg;
  assign mem[1127] = mem_1127_sv2v_reg;
  assign mem[1126] = mem_1126_sv2v_reg;
  assign mem[1125] = mem_1125_sv2v_reg;
  assign mem[1124] = mem_1124_sv2v_reg;
  assign mem[1123] = mem_1123_sv2v_reg;
  assign mem[1122] = mem_1122_sv2v_reg;
  assign mem[1121] = mem_1121_sv2v_reg;
  assign mem[1120] = mem_1120_sv2v_reg;
  assign mem[1119] = mem_1119_sv2v_reg;
  assign mem[1118] = mem_1118_sv2v_reg;
  assign mem[1117] = mem_1117_sv2v_reg;
  assign mem[1116] = mem_1116_sv2v_reg;
  assign mem[1115] = mem_1115_sv2v_reg;
  assign mem[1114] = mem_1114_sv2v_reg;
  assign mem[1113] = mem_1113_sv2v_reg;
  assign mem[1112] = mem_1112_sv2v_reg;
  assign mem[1111] = mem_1111_sv2v_reg;
  assign mem[1110] = mem_1110_sv2v_reg;
  assign mem[1109] = mem_1109_sv2v_reg;
  assign mem[1108] = mem_1108_sv2v_reg;
  assign mem[1107] = mem_1107_sv2v_reg;
  assign mem[1106] = mem_1106_sv2v_reg;
  assign mem[1105] = mem_1105_sv2v_reg;
  assign mem[1104] = mem_1104_sv2v_reg;
  assign mem[1103] = mem_1103_sv2v_reg;
  assign mem[1102] = mem_1102_sv2v_reg;
  assign mem[1101] = mem_1101_sv2v_reg;
  assign mem[1100] = mem_1100_sv2v_reg;
  assign mem[1099] = mem_1099_sv2v_reg;
  assign mem[1098] = mem_1098_sv2v_reg;
  assign mem[1097] = mem_1097_sv2v_reg;
  assign mem[1096] = mem_1096_sv2v_reg;
  assign mem[1095] = mem_1095_sv2v_reg;
  assign mem[1094] = mem_1094_sv2v_reg;
  assign mem[1093] = mem_1093_sv2v_reg;
  assign mem[1092] = mem_1092_sv2v_reg;
  assign mem[1091] = mem_1091_sv2v_reg;
  assign mem[1090] = mem_1090_sv2v_reg;
  assign mem[1089] = mem_1089_sv2v_reg;
  assign mem[1088] = mem_1088_sv2v_reg;
  assign mem[1087] = mem_1087_sv2v_reg;
  assign mem[1086] = mem_1086_sv2v_reg;
  assign mem[1085] = mem_1085_sv2v_reg;
  assign mem[1084] = mem_1084_sv2v_reg;
  assign mem[1083] = mem_1083_sv2v_reg;
  assign mem[1082] = mem_1082_sv2v_reg;
  assign mem[1081] = mem_1081_sv2v_reg;
  assign mem[1080] = mem_1080_sv2v_reg;
  assign mem[1079] = mem_1079_sv2v_reg;
  assign mem[1078] = mem_1078_sv2v_reg;
  assign mem[1077] = mem_1077_sv2v_reg;
  assign mem[1076] = mem_1076_sv2v_reg;
  assign mem[1075] = mem_1075_sv2v_reg;
  assign mem[1074] = mem_1074_sv2v_reg;
  assign mem[1073] = mem_1073_sv2v_reg;
  assign mem[1072] = mem_1072_sv2v_reg;
  assign mem[1071] = mem_1071_sv2v_reg;
  assign mem[1070] = mem_1070_sv2v_reg;
  assign mem[1069] = mem_1069_sv2v_reg;
  assign mem[1068] = mem_1068_sv2v_reg;
  assign mem[1067] = mem_1067_sv2v_reg;
  assign mem[1066] = mem_1066_sv2v_reg;
  assign mem[1065] = mem_1065_sv2v_reg;
  assign mem[1064] = mem_1064_sv2v_reg;
  assign mem[1063] = mem_1063_sv2v_reg;
  assign mem[1062] = mem_1062_sv2v_reg;
  assign mem[1061] = mem_1061_sv2v_reg;
  assign mem[1060] = mem_1060_sv2v_reg;
  assign mem[1059] = mem_1059_sv2v_reg;
  assign mem[1058] = mem_1058_sv2v_reg;
  assign mem[1057] = mem_1057_sv2v_reg;
  assign mem[1056] = mem_1056_sv2v_reg;
  assign mem[1055] = mem_1055_sv2v_reg;
  assign mem[1054] = mem_1054_sv2v_reg;
  assign mem[1053] = mem_1053_sv2v_reg;
  assign mem[1052] = mem_1052_sv2v_reg;
  assign mem[1051] = mem_1051_sv2v_reg;
  assign mem[1050] = mem_1050_sv2v_reg;
  assign mem[1049] = mem_1049_sv2v_reg;
  assign mem[1048] = mem_1048_sv2v_reg;
  assign mem[1047] = mem_1047_sv2v_reg;
  assign mem[1046] = mem_1046_sv2v_reg;
  assign mem[1045] = mem_1045_sv2v_reg;
  assign mem[1044] = mem_1044_sv2v_reg;
  assign mem[1043] = mem_1043_sv2v_reg;
  assign mem[1042] = mem_1042_sv2v_reg;
  assign mem[1041] = mem_1041_sv2v_reg;
  assign mem[1040] = mem_1040_sv2v_reg;
  assign mem[1039] = mem_1039_sv2v_reg;
  assign mem[1038] = mem_1038_sv2v_reg;
  assign mem[1037] = mem_1037_sv2v_reg;
  assign mem[1036] = mem_1036_sv2v_reg;
  assign mem[1035] = mem_1035_sv2v_reg;
  assign mem[1034] = mem_1034_sv2v_reg;
  assign mem[1033] = mem_1033_sv2v_reg;
  assign mem[1032] = mem_1032_sv2v_reg;
  assign mem[1031] = mem_1031_sv2v_reg;
  assign mem[1030] = mem_1030_sv2v_reg;
  assign mem[1029] = mem_1029_sv2v_reg;
  assign mem[1028] = mem_1028_sv2v_reg;
  assign mem[1027] = mem_1027_sv2v_reg;
  assign mem[1026] = mem_1026_sv2v_reg;
  assign mem[1025] = mem_1025_sv2v_reg;
  assign mem[1024] = mem_1024_sv2v_reg;
  assign mem[1023] = mem_1023_sv2v_reg;
  assign mem[1022] = mem_1022_sv2v_reg;
  assign mem[1021] = mem_1021_sv2v_reg;
  assign mem[1020] = mem_1020_sv2v_reg;
  assign mem[1019] = mem_1019_sv2v_reg;
  assign mem[1018] = mem_1018_sv2v_reg;
  assign mem[1017] = mem_1017_sv2v_reg;
  assign mem[1016] = mem_1016_sv2v_reg;
  assign mem[1015] = mem_1015_sv2v_reg;
  assign mem[1014] = mem_1014_sv2v_reg;
  assign mem[1013] = mem_1013_sv2v_reg;
  assign mem[1012] = mem_1012_sv2v_reg;
  assign mem[1011] = mem_1011_sv2v_reg;
  assign mem[1010] = mem_1010_sv2v_reg;
  assign mem[1009] = mem_1009_sv2v_reg;
  assign mem[1008] = mem_1008_sv2v_reg;
  assign mem[1007] = mem_1007_sv2v_reg;
  assign mem[1006] = mem_1006_sv2v_reg;
  assign mem[1005] = mem_1005_sv2v_reg;
  assign mem[1004] = mem_1004_sv2v_reg;
  assign mem[1003] = mem_1003_sv2v_reg;
  assign mem[1002] = mem_1002_sv2v_reg;
  assign mem[1001] = mem_1001_sv2v_reg;
  assign mem[1000] = mem_1000_sv2v_reg;
  assign mem[999] = mem_999_sv2v_reg;
  assign mem[998] = mem_998_sv2v_reg;
  assign mem[997] = mem_997_sv2v_reg;
  assign mem[996] = mem_996_sv2v_reg;
  assign mem[995] = mem_995_sv2v_reg;
  assign mem[994] = mem_994_sv2v_reg;
  assign mem[993] = mem_993_sv2v_reg;
  assign mem[992] = mem_992_sv2v_reg;
  assign mem[991] = mem_991_sv2v_reg;
  assign mem[990] = mem_990_sv2v_reg;
  assign mem[989] = mem_989_sv2v_reg;
  assign mem[988] = mem_988_sv2v_reg;
  assign mem[987] = mem_987_sv2v_reg;
  assign mem[986] = mem_986_sv2v_reg;
  assign mem[985] = mem_985_sv2v_reg;
  assign mem[984] = mem_984_sv2v_reg;
  assign mem[983] = mem_983_sv2v_reg;
  assign mem[982] = mem_982_sv2v_reg;
  assign mem[981] = mem_981_sv2v_reg;
  assign mem[980] = mem_980_sv2v_reg;
  assign mem[979] = mem_979_sv2v_reg;
  assign mem[978] = mem_978_sv2v_reg;
  assign mem[977] = mem_977_sv2v_reg;
  assign mem[976] = mem_976_sv2v_reg;
  assign mem[975] = mem_975_sv2v_reg;
  assign mem[974] = mem_974_sv2v_reg;
  assign mem[973] = mem_973_sv2v_reg;
  assign mem[972] = mem_972_sv2v_reg;
  assign mem[971] = mem_971_sv2v_reg;
  assign mem[970] = mem_970_sv2v_reg;
  assign mem[969] = mem_969_sv2v_reg;
  assign mem[968] = mem_968_sv2v_reg;
  assign mem[967] = mem_967_sv2v_reg;
  assign mem[966] = mem_966_sv2v_reg;
  assign mem[965] = mem_965_sv2v_reg;
  assign mem[964] = mem_964_sv2v_reg;
  assign mem[963] = mem_963_sv2v_reg;
  assign mem[962] = mem_962_sv2v_reg;
  assign mem[961] = mem_961_sv2v_reg;
  assign mem[960] = mem_960_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[571] = (N3)? mem[571] : 
                         (N0)? mem[1143] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[570] = (N3)? mem[570] : 
                         (N0)? mem[1142] : 1'b0;
  assign r_data_o[569] = (N3)? mem[569] : 
                         (N0)? mem[1141] : 1'b0;
  assign r_data_o[568] = (N3)? mem[568] : 
                         (N0)? mem[1140] : 1'b0;
  assign r_data_o[567] = (N3)? mem[567] : 
                         (N0)? mem[1139] : 1'b0;
  assign r_data_o[566] = (N3)? mem[566] : 
                         (N0)? mem[1138] : 1'b0;
  assign r_data_o[565] = (N3)? mem[565] : 
                         (N0)? mem[1137] : 1'b0;
  assign r_data_o[564] = (N3)? mem[564] : 
                         (N0)? mem[1136] : 1'b0;
  assign r_data_o[563] = (N3)? mem[563] : 
                         (N0)? mem[1135] : 1'b0;
  assign r_data_o[562] = (N3)? mem[562] : 
                         (N0)? mem[1134] : 1'b0;
  assign r_data_o[561] = (N3)? mem[561] : 
                         (N0)? mem[1133] : 1'b0;
  assign r_data_o[560] = (N3)? mem[560] : 
                         (N0)? mem[1132] : 1'b0;
  assign r_data_o[559] = (N3)? mem[559] : 
                         (N0)? mem[1131] : 1'b0;
  assign r_data_o[558] = (N3)? mem[558] : 
                         (N0)? mem[1130] : 1'b0;
  assign r_data_o[557] = (N3)? mem[557] : 
                         (N0)? mem[1129] : 1'b0;
  assign r_data_o[556] = (N3)? mem[556] : 
                         (N0)? mem[1128] : 1'b0;
  assign r_data_o[555] = (N3)? mem[555] : 
                         (N0)? mem[1127] : 1'b0;
  assign r_data_o[554] = (N3)? mem[554] : 
                         (N0)? mem[1126] : 1'b0;
  assign r_data_o[553] = (N3)? mem[553] : 
                         (N0)? mem[1125] : 1'b0;
  assign r_data_o[552] = (N3)? mem[552] : 
                         (N0)? mem[1124] : 1'b0;
  assign r_data_o[551] = (N3)? mem[551] : 
                         (N0)? mem[1123] : 1'b0;
  assign r_data_o[550] = (N3)? mem[550] : 
                         (N0)? mem[1122] : 1'b0;
  assign r_data_o[549] = (N3)? mem[549] : 
                         (N0)? mem[1121] : 1'b0;
  assign r_data_o[548] = (N3)? mem[548] : 
                         (N0)? mem[1120] : 1'b0;
  assign r_data_o[547] = (N3)? mem[547] : 
                         (N0)? mem[1119] : 1'b0;
  assign r_data_o[546] = (N3)? mem[546] : 
                         (N0)? mem[1118] : 1'b0;
  assign r_data_o[545] = (N3)? mem[545] : 
                         (N0)? mem[1117] : 1'b0;
  assign r_data_o[544] = (N3)? mem[544] : 
                         (N0)? mem[1116] : 1'b0;
  assign r_data_o[543] = (N3)? mem[543] : 
                         (N0)? mem[1115] : 1'b0;
  assign r_data_o[542] = (N3)? mem[542] : 
                         (N0)? mem[1114] : 1'b0;
  assign r_data_o[541] = (N3)? mem[541] : 
                         (N0)? mem[1113] : 1'b0;
  assign r_data_o[540] = (N3)? mem[540] : 
                         (N0)? mem[1112] : 1'b0;
  assign r_data_o[539] = (N3)? mem[539] : 
                         (N0)? mem[1111] : 1'b0;
  assign r_data_o[538] = (N3)? mem[538] : 
                         (N0)? mem[1110] : 1'b0;
  assign r_data_o[537] = (N3)? mem[537] : 
                         (N0)? mem[1109] : 1'b0;
  assign r_data_o[536] = (N3)? mem[536] : 
                         (N0)? mem[1108] : 1'b0;
  assign r_data_o[535] = (N3)? mem[535] : 
                         (N0)? mem[1107] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] : 
                         (N0)? mem[1106] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] : 
                         (N0)? mem[1105] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] : 
                         (N0)? mem[1104] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] : 
                         (N0)? mem[1103] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] : 
                         (N0)? mem[1102] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] : 
                         (N0)? mem[1101] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] : 
                         (N0)? mem[1100] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] : 
                         (N0)? mem[1099] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] : 
                         (N0)? mem[1098] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] : 
                         (N0)? mem[1097] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] : 
                         (N0)? mem[1096] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] : 
                         (N0)? mem[1095] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] : 
                         (N0)? mem[1094] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] : 
                         (N0)? mem[1093] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] : 
                         (N0)? mem[1092] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] : 
                         (N0)? mem[1091] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] : 
                         (N0)? mem[1090] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] : 
                         (N0)? mem[1089] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] : 
                         (N0)? mem[1088] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] : 
                         (N0)? mem[1087] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] : 
                         (N0)? mem[1086] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] : 
                         (N0)? mem[1085] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] : 
                         (N0)? mem[1084] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] : 
                         (N0)? mem[1083] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] : 
                         (N0)? mem[1082] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] : 
                         (N0)? mem[1081] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] : 
                         (N0)? mem[1080] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] : 
                         (N0)? mem[1079] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] : 
                         (N0)? mem[1078] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] : 
                         (N0)? mem[1077] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] : 
                         (N0)? mem[1076] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] : 
                         (N0)? mem[1075] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] : 
                         (N0)? mem[1074] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] : 
                         (N0)? mem[1073] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] : 
                         (N0)? mem[1072] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] : 
                         (N0)? mem[1071] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] : 
                         (N0)? mem[1070] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] : 
                         (N0)? mem[1069] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] : 
                         (N0)? mem[1068] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] : 
                         (N0)? mem[1067] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] : 
                         (N0)? mem[1066] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] : 
                         (N0)? mem[1065] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] : 
                         (N0)? mem[1064] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] : 
                         (N0)? mem[1063] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] : 
                         (N0)? mem[1062] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] : 
                         (N0)? mem[1061] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] : 
                         (N0)? mem[1060] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] : 
                         (N0)? mem[1059] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] : 
                         (N0)? mem[1058] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] : 
                         (N0)? mem[1057] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] : 
                         (N0)? mem[1056] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] : 
                         (N0)? mem[1055] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] : 
                         (N0)? mem[1054] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] : 
                         (N0)? mem[1053] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] : 
                         (N0)? mem[1052] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] : 
                         (N0)? mem[1051] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] : 
                         (N0)? mem[1050] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] : 
                         (N0)? mem[1049] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] : 
                         (N0)? mem[1048] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] : 
                         (N0)? mem[1047] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] : 
                         (N0)? mem[1046] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] : 
                         (N0)? mem[1045] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] : 
                         (N0)? mem[1044] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] : 
                         (N0)? mem[1043] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] : 
                         (N0)? mem[1042] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] : 
                         (N0)? mem[1041] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] : 
                         (N0)? mem[1040] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] : 
                         (N0)? mem[1039] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] : 
                         (N0)? mem[1038] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] : 
                         (N0)? mem[1037] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] : 
                         (N0)? mem[1036] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] : 
                         (N0)? mem[1035] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] : 
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] : 
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] : 
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] : 
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] : 
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] : 
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] : 
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] : 
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] : 
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] : 
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] : 
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] : 
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] : 
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] : 
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] : 
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] : 
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] : 
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] : 
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] : 
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] : 
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] : 
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] : 
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] : 
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] : 
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] : 
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] : 
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] : 
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] : 
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] : 
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] : 
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] : 
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] : 
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] : 
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] : 
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] : 
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] : 
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] : 
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] : 
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] : 
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] : 
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] : 
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] : 
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] : 
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] : 
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] : 
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] : 
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] : 
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] : 
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] : 
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] : 
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] : 
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] : 
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] : 
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] : 
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] : 
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] : 
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] : 
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] : 
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] : 
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] : 
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] : 
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] : 
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] : 
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] : 
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] : 
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] : 
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] : 
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] : 
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] : 
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] : 
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] : 
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] : 
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] : 
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] : 
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] : 
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] : 
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] : 
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] : 
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] : 
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] : 
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] : 
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] : 
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] : 
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] : 
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] : 
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] : 
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] : 
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] : 
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] : 
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] : 
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] : 
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] : 
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] : 
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] : 
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] : 
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] : 
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] : 
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] : 
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] : 
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] : 
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] : 
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] : 
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] : 
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] : 
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] : 
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] : 
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] : 
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] : 
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] : 
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] : 
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] : 
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] : 
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] : 
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] : 
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] : 
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] : 
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] : 
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] : 
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] : 
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] : 
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] : 
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] : 
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] : 
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] : 
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] : 
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] : 
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] : 
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] : 
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] : 
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] : 
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] : 
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] : 
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] : 
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] : 
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] : 
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] : 
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] : 
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] : 
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] : 
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] : 
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] : 
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] : 
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] : 
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] : 
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] : 
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] : 
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] : 
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] : 
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] : 
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] : 
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] : 
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] : 
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] : 
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] : 
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] : 
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] : 
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] : 
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] : 
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] : 
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] : 
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] : 
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] : 
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] : 
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] : 
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] : 
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] : 
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] : 
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] : 
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] : 
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] : 
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] : 
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] : 
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] : 
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] : 
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] : 
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] : 
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] : 
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] : 
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] : 
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] : 
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] : 
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] : 
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] : 
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] : 
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] : 
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] : 
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] : 
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] : 
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] : 
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] : 
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] : 
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] : 
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] : 
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] : 
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] : 
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] : 
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] : 
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] : 
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] : 
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] : 
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] : 
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] : 
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] : 
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] : 
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] : 
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] : 
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] : 
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] : 
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] : 
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] : 
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] : 
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] : 
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] : 
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] : 
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] : 
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] : 
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] : 
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] : 
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] : 
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] : 
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] : 
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] : 
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] : 
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] : 
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] : 
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] : 
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] : 
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] : 
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] : 
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] : 
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] : 
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] : 
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] : 
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] : 
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] : 
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] : 
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] : 
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] : 
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] : 
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] : 
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] : 
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] : 
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] : 
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] : 
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] : 
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] : 
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] : 
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] : 
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] : 
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] : 
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] : 
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] : 
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] : 
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] : 
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] : 
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] : 
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] : 
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] : 
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] : 
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] : 
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] : 
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] : 
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] : 
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] : 
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] : 
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] : 
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] : 
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] : 
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] : 
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] : 
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] : 
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] : 
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] : 
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] : 
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] : 
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] : 
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] : 
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] : 
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] : 
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] : 
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] : 
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] : 
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] : 
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] : 
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] : 
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] : 
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] : 
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] : 
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] : 
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] : 
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] : 
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] : 
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] : 
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] : 
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] : 
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] : 
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] : 
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] : 
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] : 
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] : 
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] : 
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] : 
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] : 
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] : 
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] : 
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] : 
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] : 
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] : 
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] : 
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] : 
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] : 
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] : 
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] : 
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] : 
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] : 
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] : 
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] : 
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] : 
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] : 
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] : 
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] : 
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] : 
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] : 
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] : 
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] : 
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] : 
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] : 
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] : 
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] : 
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] : 
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] : 
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] : 
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] : 
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] : 
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] : 
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[671] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[670] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[669] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[668] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[667] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[666] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[665] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[664] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[663] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[662] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[661] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[660] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[659] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[658] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[657] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[656] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[655] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[654] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[653] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[652] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[651] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[650] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[649] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[648] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[647] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[646] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[645] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[644] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[643] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[642] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[641] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[640] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[639] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[638] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[637] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[636] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[635] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[634] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[633] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[632] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[631] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[630] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[629] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[628] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[627] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[626] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[625] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[624] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[623] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[622] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[621] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[620] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[619] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[618] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[581] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[580] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[579] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[578] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[577] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[576] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[575] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[574] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[573] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[572] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1143_sv2v_reg <= w_data_i[571];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1142_sv2v_reg <= w_data_i[570];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1141_sv2v_reg <= w_data_i[569];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1140_sv2v_reg <= w_data_i[568];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1139_sv2v_reg <= w_data_i[567];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1138_sv2v_reg <= w_data_i[566];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1137_sv2v_reg <= w_data_i[565];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1136_sv2v_reg <= w_data_i[564];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1135_sv2v_reg <= w_data_i[563];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1134_sv2v_reg <= w_data_i[562];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1133_sv2v_reg <= w_data_i[561];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1132_sv2v_reg <= w_data_i[560];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1131_sv2v_reg <= w_data_i[559];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1130_sv2v_reg <= w_data_i[558];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1129_sv2v_reg <= w_data_i[557];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1128_sv2v_reg <= w_data_i[556];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1127_sv2v_reg <= w_data_i[555];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1126_sv2v_reg <= w_data_i[554];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1125_sv2v_reg <= w_data_i[553];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1124_sv2v_reg <= w_data_i[552];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1123_sv2v_reg <= w_data_i[551];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1122_sv2v_reg <= w_data_i[550];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1121_sv2v_reg <= w_data_i[549];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1120_sv2v_reg <= w_data_i[548];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1119_sv2v_reg <= w_data_i[547];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1118_sv2v_reg <= w_data_i[546];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1117_sv2v_reg <= w_data_i[545];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1116_sv2v_reg <= w_data_i[544];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1115_sv2v_reg <= w_data_i[543];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1114_sv2v_reg <= w_data_i[542];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1113_sv2v_reg <= w_data_i[541];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1112_sv2v_reg <= w_data_i[540];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1111_sv2v_reg <= w_data_i[539];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1110_sv2v_reg <= w_data_i[538];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1109_sv2v_reg <= w_data_i[537];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1108_sv2v_reg <= w_data_i[536];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1107_sv2v_reg <= w_data_i[535];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1106_sv2v_reg <= w_data_i[534];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1105_sv2v_reg <= w_data_i[533];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1104_sv2v_reg <= w_data_i[532];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1103_sv2v_reg <= w_data_i[531];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1102_sv2v_reg <= w_data_i[530];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1101_sv2v_reg <= w_data_i[529];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1100_sv2v_reg <= w_data_i[528];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1099_sv2v_reg <= w_data_i[527];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1098_sv2v_reg <= w_data_i[526];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1097_sv2v_reg <= w_data_i[525];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1096_sv2v_reg <= w_data_i[524];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1095_sv2v_reg <= w_data_i[523];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1094_sv2v_reg <= w_data_i[522];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1093_sv2v_reg <= w_data_i[521];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1092_sv2v_reg <= w_data_i[520];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1091_sv2v_reg <= w_data_i[519];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1090_sv2v_reg <= w_data_i[518];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1089_sv2v_reg <= w_data_i[517];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1088_sv2v_reg <= w_data_i[516];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1087_sv2v_reg <= w_data_i[515];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1086_sv2v_reg <= w_data_i[514];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1085_sv2v_reg <= w_data_i[513];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1084_sv2v_reg <= w_data_i[512];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1083_sv2v_reg <= w_data_i[511];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1082_sv2v_reg <= w_data_i[510];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1081_sv2v_reg <= w_data_i[509];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1080_sv2v_reg <= w_data_i[508];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1079_sv2v_reg <= w_data_i[507];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1078_sv2v_reg <= w_data_i[506];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1077_sv2v_reg <= w_data_i[505];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1076_sv2v_reg <= w_data_i[504];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1075_sv2v_reg <= w_data_i[503];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1074_sv2v_reg <= w_data_i[502];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1073_sv2v_reg <= w_data_i[501];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1072_sv2v_reg <= w_data_i[500];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1071_sv2v_reg <= w_data_i[499];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1070_sv2v_reg <= w_data_i[498];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1069_sv2v_reg <= w_data_i[497];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1068_sv2v_reg <= w_data_i[496];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1067_sv2v_reg <= w_data_i[495];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1066_sv2v_reg <= w_data_i[494];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1065_sv2v_reg <= w_data_i[493];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1064_sv2v_reg <= w_data_i[492];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1063_sv2v_reg <= w_data_i[491];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1062_sv2v_reg <= w_data_i[490];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1061_sv2v_reg <= w_data_i[489];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1060_sv2v_reg <= w_data_i[488];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1059_sv2v_reg <= w_data_i[487];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1058_sv2v_reg <= w_data_i[486];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1057_sv2v_reg <= w_data_i[485];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1056_sv2v_reg <= w_data_i[484];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1055_sv2v_reg <= w_data_i[483];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1054_sv2v_reg <= w_data_i[482];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1053_sv2v_reg <= w_data_i[481];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1052_sv2v_reg <= w_data_i[480];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1051_sv2v_reg <= w_data_i[479];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1050_sv2v_reg <= w_data_i[478];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1049_sv2v_reg <= w_data_i[477];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1048_sv2v_reg <= w_data_i[476];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1047_sv2v_reg <= w_data_i[475];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1046_sv2v_reg <= w_data_i[474];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_1045_sv2v_reg <= w_data_i[473];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1044_sv2v_reg <= w_data_i[472];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1043_sv2v_reg <= w_data_i[471];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1042_sv2v_reg <= w_data_i[470];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1041_sv2v_reg <= w_data_i[469];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1040_sv2v_reg <= w_data_i[468];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1039_sv2v_reg <= w_data_i[467];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1038_sv2v_reg <= w_data_i[466];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1037_sv2v_reg <= w_data_i[465];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1036_sv2v_reg <= w_data_i[464];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1035_sv2v_reg <= w_data_i[463];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1034_sv2v_reg <= w_data_i[462];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1033_sv2v_reg <= w_data_i[461];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1032_sv2v_reg <= w_data_i[460];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1031_sv2v_reg <= w_data_i[459];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1030_sv2v_reg <= w_data_i[458];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1029_sv2v_reg <= w_data_i[457];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1028_sv2v_reg <= w_data_i[456];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1027_sv2v_reg <= w_data_i[455];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1026_sv2v_reg <= w_data_i[454];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1025_sv2v_reg <= w_data_i[453];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1024_sv2v_reg <= w_data_i[452];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1023_sv2v_reg <= w_data_i[451];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1022_sv2v_reg <= w_data_i[450];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1021_sv2v_reg <= w_data_i[449];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1020_sv2v_reg <= w_data_i[448];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1019_sv2v_reg <= w_data_i[447];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1018_sv2v_reg <= w_data_i[446];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1017_sv2v_reg <= w_data_i[445];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1016_sv2v_reg <= w_data_i[444];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1015_sv2v_reg <= w_data_i[443];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1014_sv2v_reg <= w_data_i[442];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1013_sv2v_reg <= w_data_i[441];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1012_sv2v_reg <= w_data_i[440];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1011_sv2v_reg <= w_data_i[439];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1010_sv2v_reg <= w_data_i[438];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1009_sv2v_reg <= w_data_i[437];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1008_sv2v_reg <= w_data_i[436];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1007_sv2v_reg <= w_data_i[435];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1006_sv2v_reg <= w_data_i[434];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1005_sv2v_reg <= w_data_i[433];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1004_sv2v_reg <= w_data_i[432];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1003_sv2v_reg <= w_data_i[431];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1002_sv2v_reg <= w_data_i[430];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1001_sv2v_reg <= w_data_i[429];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_1000_sv2v_reg <= w_data_i[428];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_999_sv2v_reg <= w_data_i[427];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_998_sv2v_reg <= w_data_i[426];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_997_sv2v_reg <= w_data_i[425];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_996_sv2v_reg <= w_data_i[424];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_995_sv2v_reg <= w_data_i[423];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_994_sv2v_reg <= w_data_i[422];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_993_sv2v_reg <= w_data_i[421];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_992_sv2v_reg <= w_data_i[420];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_991_sv2v_reg <= w_data_i[419];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_990_sv2v_reg <= w_data_i[418];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_989_sv2v_reg <= w_data_i[417];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_988_sv2v_reg <= w_data_i[416];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_987_sv2v_reg <= w_data_i[415];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_986_sv2v_reg <= w_data_i[414];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_985_sv2v_reg <= w_data_i[413];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_984_sv2v_reg <= w_data_i[412];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_983_sv2v_reg <= w_data_i[411];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_982_sv2v_reg <= w_data_i[410];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_981_sv2v_reg <= w_data_i[409];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_980_sv2v_reg <= w_data_i[408];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_979_sv2v_reg <= w_data_i[407];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_978_sv2v_reg <= w_data_i[406];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_977_sv2v_reg <= w_data_i[405];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_976_sv2v_reg <= w_data_i[404];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_975_sv2v_reg <= w_data_i[403];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_974_sv2v_reg <= w_data_i[402];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_973_sv2v_reg <= w_data_i[401];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_972_sv2v_reg <= w_data_i[400];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_971_sv2v_reg <= w_data_i[399];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_970_sv2v_reg <= w_data_i[398];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_969_sv2v_reg <= w_data_i[397];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_968_sv2v_reg <= w_data_i[396];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_967_sv2v_reg <= w_data_i[395];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_966_sv2v_reg <= w_data_i[394];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_965_sv2v_reg <= w_data_i[393];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_964_sv2v_reg <= w_data_i[392];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_963_sv2v_reg <= w_data_i[391];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_962_sv2v_reg <= w_data_i[390];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_961_sv2v_reg <= w_data_i[389];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_960_sv2v_reg <= w_data_i[388];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_959_sv2v_reg <= w_data_i[387];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_958_sv2v_reg <= w_data_i[386];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_957_sv2v_reg <= w_data_i[385];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_956_sv2v_reg <= w_data_i[384];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_955_sv2v_reg <= w_data_i[383];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_954_sv2v_reg <= w_data_i[382];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_953_sv2v_reg <= w_data_i[381];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_952_sv2v_reg <= w_data_i[380];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_951_sv2v_reg <= w_data_i[379];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_950_sv2v_reg <= w_data_i[378];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_949_sv2v_reg <= w_data_i[377];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_948_sv2v_reg <= w_data_i[376];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_947_sv2v_reg <= w_data_i[375];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_946_sv2v_reg <= w_data_i[374];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_945_sv2v_reg <= w_data_i[373];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_944_sv2v_reg <= w_data_i[372];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_943_sv2v_reg <= w_data_i[371];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_942_sv2v_reg <= w_data_i[370];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_941_sv2v_reg <= w_data_i[369];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_940_sv2v_reg <= w_data_i[368];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_939_sv2v_reg <= w_data_i[367];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_938_sv2v_reg <= w_data_i[366];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_937_sv2v_reg <= w_data_i[365];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_936_sv2v_reg <= w_data_i[364];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_935_sv2v_reg <= w_data_i[363];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_934_sv2v_reg <= w_data_i[362];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_933_sv2v_reg <= w_data_i[361];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_932_sv2v_reg <= w_data_i[360];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_931_sv2v_reg <= w_data_i[359];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_930_sv2v_reg <= w_data_i[358];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_929_sv2v_reg <= w_data_i[357];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_928_sv2v_reg <= w_data_i[356];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_927_sv2v_reg <= w_data_i[355];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_926_sv2v_reg <= w_data_i[354];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_925_sv2v_reg <= w_data_i[353];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_924_sv2v_reg <= w_data_i[352];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_923_sv2v_reg <= w_data_i[351];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_922_sv2v_reg <= w_data_i[350];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_921_sv2v_reg <= w_data_i[349];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_920_sv2v_reg <= w_data_i[348];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_919_sv2v_reg <= w_data_i[347];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_918_sv2v_reg <= w_data_i[346];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_917_sv2v_reg <= w_data_i[345];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_916_sv2v_reg <= w_data_i[344];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_915_sv2v_reg <= w_data_i[343];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_914_sv2v_reg <= w_data_i[342];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_913_sv2v_reg <= w_data_i[341];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_912_sv2v_reg <= w_data_i[340];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_911_sv2v_reg <= w_data_i[339];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_910_sv2v_reg <= w_data_i[338];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_909_sv2v_reg <= w_data_i[337];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_908_sv2v_reg <= w_data_i[336];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_907_sv2v_reg <= w_data_i[335];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_906_sv2v_reg <= w_data_i[334];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_905_sv2v_reg <= w_data_i[333];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_904_sv2v_reg <= w_data_i[332];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_903_sv2v_reg <= w_data_i[331];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_902_sv2v_reg <= w_data_i[330];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_901_sv2v_reg <= w_data_i[329];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_900_sv2v_reg <= w_data_i[328];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_899_sv2v_reg <= w_data_i[327];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_898_sv2v_reg <= w_data_i[326];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_897_sv2v_reg <= w_data_i[325];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_896_sv2v_reg <= w_data_i[324];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_895_sv2v_reg <= w_data_i[323];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_894_sv2v_reg <= w_data_i[322];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_893_sv2v_reg <= w_data_i[321];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_892_sv2v_reg <= w_data_i[320];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_891_sv2v_reg <= w_data_i[319];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_890_sv2v_reg <= w_data_i[318];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_889_sv2v_reg <= w_data_i[317];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_888_sv2v_reg <= w_data_i[316];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_887_sv2v_reg <= w_data_i[315];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_886_sv2v_reg <= w_data_i[314];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_885_sv2v_reg <= w_data_i[313];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_884_sv2v_reg <= w_data_i[312];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_883_sv2v_reg <= w_data_i[311];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_882_sv2v_reg <= w_data_i[310];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_881_sv2v_reg <= w_data_i[309];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_880_sv2v_reg <= w_data_i[308];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_879_sv2v_reg <= w_data_i[307];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_878_sv2v_reg <= w_data_i[306];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_877_sv2v_reg <= w_data_i[305];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_876_sv2v_reg <= w_data_i[304];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_875_sv2v_reg <= w_data_i[303];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_874_sv2v_reg <= w_data_i[302];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_873_sv2v_reg <= w_data_i[301];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_872_sv2v_reg <= w_data_i[300];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_871_sv2v_reg <= w_data_i[299];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_870_sv2v_reg <= w_data_i[298];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_869_sv2v_reg <= w_data_i[297];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_868_sv2v_reg <= w_data_i[296];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_867_sv2v_reg <= w_data_i[295];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_866_sv2v_reg <= w_data_i[294];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_865_sv2v_reg <= w_data_i[293];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_864_sv2v_reg <= w_data_i[292];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_863_sv2v_reg <= w_data_i[291];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_862_sv2v_reg <= w_data_i[290];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_861_sv2v_reg <= w_data_i[289];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_860_sv2v_reg <= w_data_i[288];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_859_sv2v_reg <= w_data_i[287];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_858_sv2v_reg <= w_data_i[286];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_857_sv2v_reg <= w_data_i[285];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_856_sv2v_reg <= w_data_i[284];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_855_sv2v_reg <= w_data_i[283];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_854_sv2v_reg <= w_data_i[282];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_853_sv2v_reg <= w_data_i[281];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_852_sv2v_reg <= w_data_i[280];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_851_sv2v_reg <= w_data_i[279];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_850_sv2v_reg <= w_data_i[278];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_849_sv2v_reg <= w_data_i[277];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_848_sv2v_reg <= w_data_i[276];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_847_sv2v_reg <= w_data_i[275];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_846_sv2v_reg <= w_data_i[274];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_845_sv2v_reg <= w_data_i[273];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_844_sv2v_reg <= w_data_i[272];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_843_sv2v_reg <= w_data_i[271];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_842_sv2v_reg <= w_data_i[270];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_841_sv2v_reg <= w_data_i[269];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_840_sv2v_reg <= w_data_i[268];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_839_sv2v_reg <= w_data_i[267];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_838_sv2v_reg <= w_data_i[266];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_837_sv2v_reg <= w_data_i[265];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_836_sv2v_reg <= w_data_i[264];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_835_sv2v_reg <= w_data_i[263];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_834_sv2v_reg <= w_data_i[262];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_833_sv2v_reg <= w_data_i[261];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_832_sv2v_reg <= w_data_i[260];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_831_sv2v_reg <= w_data_i[259];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_830_sv2v_reg <= w_data_i[258];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_829_sv2v_reg <= w_data_i[257];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_828_sv2v_reg <= w_data_i[256];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_827_sv2v_reg <= w_data_i[255];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_826_sv2v_reg <= w_data_i[254];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_825_sv2v_reg <= w_data_i[253];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_824_sv2v_reg <= w_data_i[252];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_823_sv2v_reg <= w_data_i[251];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_822_sv2v_reg <= w_data_i[250];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_821_sv2v_reg <= w_data_i[249];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_820_sv2v_reg <= w_data_i[248];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_819_sv2v_reg <= w_data_i[247];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_818_sv2v_reg <= w_data_i[246];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_817_sv2v_reg <= w_data_i[245];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_816_sv2v_reg <= w_data_i[244];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_815_sv2v_reg <= w_data_i[243];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_814_sv2v_reg <= w_data_i[242];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_813_sv2v_reg <= w_data_i[241];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_812_sv2v_reg <= w_data_i[240];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_811_sv2v_reg <= w_data_i[239];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_810_sv2v_reg <= w_data_i[238];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_809_sv2v_reg <= w_data_i[237];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_808_sv2v_reg <= w_data_i[236];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_807_sv2v_reg <= w_data_i[235];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_806_sv2v_reg <= w_data_i[234];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_805_sv2v_reg <= w_data_i[233];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_804_sv2v_reg <= w_data_i[232];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_803_sv2v_reg <= w_data_i[231];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_802_sv2v_reg <= w_data_i[230];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_801_sv2v_reg <= w_data_i[229];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_800_sv2v_reg <= w_data_i[228];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_799_sv2v_reg <= w_data_i[227];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_798_sv2v_reg <= w_data_i[226];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_797_sv2v_reg <= w_data_i[225];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_796_sv2v_reg <= w_data_i[224];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_795_sv2v_reg <= w_data_i[223];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_794_sv2v_reg <= w_data_i[222];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_793_sv2v_reg <= w_data_i[221];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_792_sv2v_reg <= w_data_i[220];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_791_sv2v_reg <= w_data_i[219];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_790_sv2v_reg <= w_data_i[218];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_789_sv2v_reg <= w_data_i[217];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_788_sv2v_reg <= w_data_i[216];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_787_sv2v_reg <= w_data_i[215];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_786_sv2v_reg <= w_data_i[214];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_785_sv2v_reg <= w_data_i[213];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_784_sv2v_reg <= w_data_i[212];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_783_sv2v_reg <= w_data_i[211];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_782_sv2v_reg <= w_data_i[210];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_781_sv2v_reg <= w_data_i[209];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_780_sv2v_reg <= w_data_i[208];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_779_sv2v_reg <= w_data_i[207];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_778_sv2v_reg <= w_data_i[206];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_777_sv2v_reg <= w_data_i[205];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_776_sv2v_reg <= w_data_i[204];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_775_sv2v_reg <= w_data_i[203];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_774_sv2v_reg <= w_data_i[202];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_773_sv2v_reg <= w_data_i[201];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_772_sv2v_reg <= w_data_i[200];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_771_sv2v_reg <= w_data_i[199];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_770_sv2v_reg <= w_data_i[198];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_769_sv2v_reg <= w_data_i[197];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_768_sv2v_reg <= w_data_i[196];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_767_sv2v_reg <= w_data_i[195];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_766_sv2v_reg <= w_data_i[194];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_765_sv2v_reg <= w_data_i[193];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_764_sv2v_reg <= w_data_i[192];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_763_sv2v_reg <= w_data_i[191];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_762_sv2v_reg <= w_data_i[190];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_761_sv2v_reg <= w_data_i[189];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_760_sv2v_reg <= w_data_i[188];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_759_sv2v_reg <= w_data_i[187];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_758_sv2v_reg <= w_data_i[186];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_757_sv2v_reg <= w_data_i[185];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_756_sv2v_reg <= w_data_i[184];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_755_sv2v_reg <= w_data_i[183];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_754_sv2v_reg <= w_data_i[182];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_753_sv2v_reg <= w_data_i[181];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_752_sv2v_reg <= w_data_i[180];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_751_sv2v_reg <= w_data_i[179];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_750_sv2v_reg <= w_data_i[178];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_749_sv2v_reg <= w_data_i[177];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_748_sv2v_reg <= w_data_i[176];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_747_sv2v_reg <= w_data_i[175];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_746_sv2v_reg <= w_data_i[174];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_745_sv2v_reg <= w_data_i[173];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_744_sv2v_reg <= w_data_i[172];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_743_sv2v_reg <= w_data_i[171];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_742_sv2v_reg <= w_data_i[170];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_741_sv2v_reg <= w_data_i[169];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_740_sv2v_reg <= w_data_i[168];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_739_sv2v_reg <= w_data_i[167];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_738_sv2v_reg <= w_data_i[166];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_737_sv2v_reg <= w_data_i[165];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_736_sv2v_reg <= w_data_i[164];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_735_sv2v_reg <= w_data_i[163];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_734_sv2v_reg <= w_data_i[162];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_733_sv2v_reg <= w_data_i[161];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_732_sv2v_reg <= w_data_i[160];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_731_sv2v_reg <= w_data_i[159];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_730_sv2v_reg <= w_data_i[158];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_729_sv2v_reg <= w_data_i[157];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_728_sv2v_reg <= w_data_i[156];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_727_sv2v_reg <= w_data_i[155];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_726_sv2v_reg <= w_data_i[154];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_725_sv2v_reg <= w_data_i[153];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_724_sv2v_reg <= w_data_i[152];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_723_sv2v_reg <= w_data_i[151];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_722_sv2v_reg <= w_data_i[150];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_721_sv2v_reg <= w_data_i[149];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_720_sv2v_reg <= w_data_i[148];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_719_sv2v_reg <= w_data_i[147];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_718_sv2v_reg <= w_data_i[146];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_717_sv2v_reg <= w_data_i[145];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_716_sv2v_reg <= w_data_i[144];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_715_sv2v_reg <= w_data_i[143];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_714_sv2v_reg <= w_data_i[142];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_713_sv2v_reg <= w_data_i[141];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_712_sv2v_reg <= w_data_i[140];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_711_sv2v_reg <= w_data_i[139];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_710_sv2v_reg <= w_data_i[138];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_709_sv2v_reg <= w_data_i[137];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_708_sv2v_reg <= w_data_i[136];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_707_sv2v_reg <= w_data_i[135];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_706_sv2v_reg <= w_data_i[134];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_705_sv2v_reg <= w_data_i[133];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_704_sv2v_reg <= w_data_i[132];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_703_sv2v_reg <= w_data_i[131];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_702_sv2v_reg <= w_data_i[130];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_701_sv2v_reg <= w_data_i[129];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_700_sv2v_reg <= w_data_i[128];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_699_sv2v_reg <= w_data_i[127];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_698_sv2v_reg <= w_data_i[126];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_697_sv2v_reg <= w_data_i[125];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_696_sv2v_reg <= w_data_i[124];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_695_sv2v_reg <= w_data_i[123];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_694_sv2v_reg <= w_data_i[122];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_693_sv2v_reg <= w_data_i[121];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_692_sv2v_reg <= w_data_i[120];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_691_sv2v_reg <= w_data_i[119];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_690_sv2v_reg <= w_data_i[118];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_689_sv2v_reg <= w_data_i[117];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_688_sv2v_reg <= w_data_i[116];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_687_sv2v_reg <= w_data_i[115];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_686_sv2v_reg <= w_data_i[114];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_685_sv2v_reg <= w_data_i[113];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_684_sv2v_reg <= w_data_i[112];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_683_sv2v_reg <= w_data_i[111];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_682_sv2v_reg <= w_data_i[110];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_681_sv2v_reg <= w_data_i[109];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_680_sv2v_reg <= w_data_i[108];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_679_sv2v_reg <= w_data_i[107];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_678_sv2v_reg <= w_data_i[106];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_677_sv2v_reg <= w_data_i[105];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_676_sv2v_reg <= w_data_i[104];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_675_sv2v_reg <= w_data_i[103];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_674_sv2v_reg <= w_data_i[102];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_673_sv2v_reg <= w_data_i[101];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_672_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_671_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_670_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_669_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_668_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_667_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_666_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_665_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_664_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_663_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_662_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_661_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_660_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_659_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_658_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_657_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_656_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_655_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_654_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_653_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_652_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_651_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_650_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_649_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_648_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_647_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_646_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_645_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_644_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_643_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_642_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_641_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_640_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_639_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_638_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_637_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_636_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_635_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_634_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_633_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_632_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_631_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_630_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_629_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_628_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_627_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_626_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_625_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_624_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_623_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_622_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_621_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_620_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_619_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_618_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_617_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_616_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_615_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_614_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_613_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_612_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_611_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_610_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_609_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_608_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_607_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_606_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_605_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_604_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_603_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_602_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_601_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_600_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_599_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_598_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_597_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_596_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_595_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_594_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_593_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_592_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_591_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_590_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_589_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_588_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_587_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_586_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_585_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_584_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_583_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_582_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_581_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_580_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_579_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_578_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem_577_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem_576_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N16) begin
      mem_575_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N15) begin
      mem_574_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N14) begin
      mem_573_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N13) begin
      mem_572_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_571_sv2v_reg <= w_data_i[571];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_570_sv2v_reg <= w_data_i[570];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_569_sv2v_reg <= w_data_i[569];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_568_sv2v_reg <= w_data_i[568];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_567_sv2v_reg <= w_data_i[567];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_566_sv2v_reg <= w_data_i[566];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_565_sv2v_reg <= w_data_i[565];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_564_sv2v_reg <= w_data_i[564];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_563_sv2v_reg <= w_data_i[563];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_562_sv2v_reg <= w_data_i[562];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_561_sv2v_reg <= w_data_i[561];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_560_sv2v_reg <= w_data_i[560];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_559_sv2v_reg <= w_data_i[559];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_558_sv2v_reg <= w_data_i[558];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_557_sv2v_reg <= w_data_i[557];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_556_sv2v_reg <= w_data_i[556];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_555_sv2v_reg <= w_data_i[555];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_554_sv2v_reg <= w_data_i[554];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_553_sv2v_reg <= w_data_i[553];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_552_sv2v_reg <= w_data_i[552];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_551_sv2v_reg <= w_data_i[551];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_550_sv2v_reg <= w_data_i[550];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_549_sv2v_reg <= w_data_i[549];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_548_sv2v_reg <= w_data_i[548];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_547_sv2v_reg <= w_data_i[547];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_546_sv2v_reg <= w_data_i[546];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_545_sv2v_reg <= w_data_i[545];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_544_sv2v_reg <= w_data_i[544];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_543_sv2v_reg <= w_data_i[543];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_542_sv2v_reg <= w_data_i[542];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_541_sv2v_reg <= w_data_i[541];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_540_sv2v_reg <= w_data_i[540];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_539_sv2v_reg <= w_data_i[539];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_538_sv2v_reg <= w_data_i[538];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_537_sv2v_reg <= w_data_i[537];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_536_sv2v_reg <= w_data_i[536];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_535_sv2v_reg <= w_data_i[535];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_534_sv2v_reg <= w_data_i[534];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_533_sv2v_reg <= w_data_i[533];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_532_sv2v_reg <= w_data_i[532];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_531_sv2v_reg <= w_data_i[531];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_530_sv2v_reg <= w_data_i[530];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_529_sv2v_reg <= w_data_i[529];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_528_sv2v_reg <= w_data_i[528];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_527_sv2v_reg <= w_data_i[527];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_526_sv2v_reg <= w_data_i[526];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_525_sv2v_reg <= w_data_i[525];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_524_sv2v_reg <= w_data_i[524];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_523_sv2v_reg <= w_data_i[523];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_522_sv2v_reg <= w_data_i[522];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_521_sv2v_reg <= w_data_i[521];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_520_sv2v_reg <= w_data_i[520];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_519_sv2v_reg <= w_data_i[519];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_518_sv2v_reg <= w_data_i[518];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_517_sv2v_reg <= w_data_i[517];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_516_sv2v_reg <= w_data_i[516];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_515_sv2v_reg <= w_data_i[515];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_514_sv2v_reg <= w_data_i[514];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_513_sv2v_reg <= w_data_i[513];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_512_sv2v_reg <= w_data_i[512];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_511_sv2v_reg <= w_data_i[511];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_510_sv2v_reg <= w_data_i[510];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_509_sv2v_reg <= w_data_i[509];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_508_sv2v_reg <= w_data_i[508];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_507_sv2v_reg <= w_data_i[507];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_506_sv2v_reg <= w_data_i[506];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_505_sv2v_reg <= w_data_i[505];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_504_sv2v_reg <= w_data_i[504];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_503_sv2v_reg <= w_data_i[503];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_502_sv2v_reg <= w_data_i[502];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_501_sv2v_reg <= w_data_i[501];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_500_sv2v_reg <= w_data_i[500];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_499_sv2v_reg <= w_data_i[499];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_498_sv2v_reg <= w_data_i[498];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_497_sv2v_reg <= w_data_i[497];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_496_sv2v_reg <= w_data_i[496];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_495_sv2v_reg <= w_data_i[495];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_494_sv2v_reg <= w_data_i[494];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_493_sv2v_reg <= w_data_i[493];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_492_sv2v_reg <= w_data_i[492];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_491_sv2v_reg <= w_data_i[491];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_490_sv2v_reg <= w_data_i[490];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_489_sv2v_reg <= w_data_i[489];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_488_sv2v_reg <= w_data_i[488];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_487_sv2v_reg <= w_data_i[487];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_486_sv2v_reg <= w_data_i[486];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_485_sv2v_reg <= w_data_i[485];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_484_sv2v_reg <= w_data_i[484];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_483_sv2v_reg <= w_data_i[483];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_482_sv2v_reg <= w_data_i[482];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_481_sv2v_reg <= w_data_i[481];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_480_sv2v_reg <= w_data_i[480];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_479_sv2v_reg <= w_data_i[479];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_478_sv2v_reg <= w_data_i[478];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_477_sv2v_reg <= w_data_i[477];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_476_sv2v_reg <= w_data_i[476];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_475_sv2v_reg <= w_data_i[475];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_474_sv2v_reg <= w_data_i[474];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_473_sv2v_reg <= w_data_i[473];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_472_sv2v_reg <= w_data_i[472];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_471_sv2v_reg <= w_data_i[471];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_470_sv2v_reg <= w_data_i[470];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_469_sv2v_reg <= w_data_i[469];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_468_sv2v_reg <= w_data_i[468];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_467_sv2v_reg <= w_data_i[467];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_466_sv2v_reg <= w_data_i[466];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_465_sv2v_reg <= w_data_i[465];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_464_sv2v_reg <= w_data_i[464];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_463_sv2v_reg <= w_data_i[463];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_462_sv2v_reg <= w_data_i[462];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_461_sv2v_reg <= w_data_i[461];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_460_sv2v_reg <= w_data_i[460];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_459_sv2v_reg <= w_data_i[459];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_458_sv2v_reg <= w_data_i[458];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_457_sv2v_reg <= w_data_i[457];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_456_sv2v_reg <= w_data_i[456];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_455_sv2v_reg <= w_data_i[455];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_454_sv2v_reg <= w_data_i[454];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_453_sv2v_reg <= w_data_i[453];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_452_sv2v_reg <= w_data_i[452];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_451_sv2v_reg <= w_data_i[451];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_450_sv2v_reg <= w_data_i[450];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_449_sv2v_reg <= w_data_i[449];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_448_sv2v_reg <= w_data_i[448];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_447_sv2v_reg <= w_data_i[447];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_446_sv2v_reg <= w_data_i[446];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_445_sv2v_reg <= w_data_i[445];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_444_sv2v_reg <= w_data_i[444];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_443_sv2v_reg <= w_data_i[443];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_442_sv2v_reg <= w_data_i[442];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_441_sv2v_reg <= w_data_i[441];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_440_sv2v_reg <= w_data_i[440];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_439_sv2v_reg <= w_data_i[439];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_438_sv2v_reg <= w_data_i[438];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_437_sv2v_reg <= w_data_i[437];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_436_sv2v_reg <= w_data_i[436];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_435_sv2v_reg <= w_data_i[435];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_434_sv2v_reg <= w_data_i[434];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_433_sv2v_reg <= w_data_i[433];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_432_sv2v_reg <= w_data_i[432];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_431_sv2v_reg <= w_data_i[431];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_430_sv2v_reg <= w_data_i[430];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_429_sv2v_reg <= w_data_i[429];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_428_sv2v_reg <= w_data_i[428];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_427_sv2v_reg <= w_data_i[427];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_426_sv2v_reg <= w_data_i[426];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_425_sv2v_reg <= w_data_i[425];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_424_sv2v_reg <= w_data_i[424];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_423_sv2v_reg <= w_data_i[423];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_422_sv2v_reg <= w_data_i[422];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_421_sv2v_reg <= w_data_i[421];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_420_sv2v_reg <= w_data_i[420];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_419_sv2v_reg <= w_data_i[419];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_418_sv2v_reg <= w_data_i[418];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_417_sv2v_reg <= w_data_i[417];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_416_sv2v_reg <= w_data_i[416];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_415_sv2v_reg <= w_data_i[415];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_414_sv2v_reg <= w_data_i[414];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_413_sv2v_reg <= w_data_i[413];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_412_sv2v_reg <= w_data_i[412];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_411_sv2v_reg <= w_data_i[411];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_410_sv2v_reg <= w_data_i[410];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_409_sv2v_reg <= w_data_i[409];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_408_sv2v_reg <= w_data_i[408];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_407_sv2v_reg <= w_data_i[407];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_406_sv2v_reg <= w_data_i[406];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_405_sv2v_reg <= w_data_i[405];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_404_sv2v_reg <= w_data_i[404];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_403_sv2v_reg <= w_data_i[403];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_402_sv2v_reg <= w_data_i[402];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_401_sv2v_reg <= w_data_i[401];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_400_sv2v_reg <= w_data_i[400];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_399_sv2v_reg <= w_data_i[399];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_398_sv2v_reg <= w_data_i[398];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_397_sv2v_reg <= w_data_i[397];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_396_sv2v_reg <= w_data_i[396];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_395_sv2v_reg <= w_data_i[395];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_394_sv2v_reg <= w_data_i[394];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_393_sv2v_reg <= w_data_i[393];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_392_sv2v_reg <= w_data_i[392];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_391_sv2v_reg <= w_data_i[391];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_390_sv2v_reg <= w_data_i[390];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_389_sv2v_reg <= w_data_i[389];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_388_sv2v_reg <= w_data_i[388];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_387_sv2v_reg <= w_data_i[387];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_386_sv2v_reg <= w_data_i[386];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_385_sv2v_reg <= w_data_i[385];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_384_sv2v_reg <= w_data_i[384];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_383_sv2v_reg <= w_data_i[383];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_382_sv2v_reg <= w_data_i[382];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_381_sv2v_reg <= w_data_i[381];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_380_sv2v_reg <= w_data_i[380];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_379_sv2v_reg <= w_data_i[379];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_378_sv2v_reg <= w_data_i[378];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_377_sv2v_reg <= w_data_i[377];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_376_sv2v_reg <= w_data_i[376];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_375_sv2v_reg <= w_data_i[375];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_374_sv2v_reg <= w_data_i[374];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_373_sv2v_reg <= w_data_i[373];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_372_sv2v_reg <= w_data_i[372];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_371_sv2v_reg <= w_data_i[371];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_370_sv2v_reg <= w_data_i[370];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_369_sv2v_reg <= w_data_i[369];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_368_sv2v_reg <= w_data_i[368];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_367_sv2v_reg <= w_data_i[367];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_366_sv2v_reg <= w_data_i[366];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_365_sv2v_reg <= w_data_i[365];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_364_sv2v_reg <= w_data_i[364];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_363_sv2v_reg <= w_data_i[363];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_362_sv2v_reg <= w_data_i[362];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_361_sv2v_reg <= w_data_i[361];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_360_sv2v_reg <= w_data_i[360];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_359_sv2v_reg <= w_data_i[359];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_358_sv2v_reg <= w_data_i[358];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_357_sv2v_reg <= w_data_i[357];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_356_sv2v_reg <= w_data_i[356];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_355_sv2v_reg <= w_data_i[355];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_354_sv2v_reg <= w_data_i[354];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_353_sv2v_reg <= w_data_i[353];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_352_sv2v_reg <= w_data_i[352];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_351_sv2v_reg <= w_data_i[351];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_350_sv2v_reg <= w_data_i[350];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_349_sv2v_reg <= w_data_i[349];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_348_sv2v_reg <= w_data_i[348];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_347_sv2v_reg <= w_data_i[347];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_346_sv2v_reg <= w_data_i[346];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_345_sv2v_reg <= w_data_i[345];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_344_sv2v_reg <= w_data_i[344];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_343_sv2v_reg <= w_data_i[343];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_342_sv2v_reg <= w_data_i[342];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_341_sv2v_reg <= w_data_i[341];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_340_sv2v_reg <= w_data_i[340];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_339_sv2v_reg <= w_data_i[339];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_338_sv2v_reg <= w_data_i[338];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_337_sv2v_reg <= w_data_i[337];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_336_sv2v_reg <= w_data_i[336];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_335_sv2v_reg <= w_data_i[335];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_334_sv2v_reg <= w_data_i[334];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_333_sv2v_reg <= w_data_i[333];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_332_sv2v_reg <= w_data_i[332];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_331_sv2v_reg <= w_data_i[331];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_330_sv2v_reg <= w_data_i[330];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_329_sv2v_reg <= w_data_i[329];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_328_sv2v_reg <= w_data_i[328];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_327_sv2v_reg <= w_data_i[327];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_326_sv2v_reg <= w_data_i[326];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_325_sv2v_reg <= w_data_i[325];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_324_sv2v_reg <= w_data_i[324];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_323_sv2v_reg <= w_data_i[323];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_322_sv2v_reg <= w_data_i[322];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_321_sv2v_reg <= w_data_i[321];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_320_sv2v_reg <= w_data_i[320];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_319_sv2v_reg <= w_data_i[319];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_318_sv2v_reg <= w_data_i[318];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_317_sv2v_reg <= w_data_i[317];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_316_sv2v_reg <= w_data_i[316];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_315_sv2v_reg <= w_data_i[315];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_314_sv2v_reg <= w_data_i[314];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_313_sv2v_reg <= w_data_i[313];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_312_sv2v_reg <= w_data_i[312];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_311_sv2v_reg <= w_data_i[311];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_310_sv2v_reg <= w_data_i[310];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_309_sv2v_reg <= w_data_i[309];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_308_sv2v_reg <= w_data_i[308];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_307_sv2v_reg <= w_data_i[307];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_306_sv2v_reg <= w_data_i[306];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_305_sv2v_reg <= w_data_i[305];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_304_sv2v_reg <= w_data_i[304];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_303_sv2v_reg <= w_data_i[303];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_302_sv2v_reg <= w_data_i[302];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_301_sv2v_reg <= w_data_i[301];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_300_sv2v_reg <= w_data_i[300];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_299_sv2v_reg <= w_data_i[299];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_298_sv2v_reg <= w_data_i[298];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_297_sv2v_reg <= w_data_i[297];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_296_sv2v_reg <= w_data_i[296];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_295_sv2v_reg <= w_data_i[295];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_294_sv2v_reg <= w_data_i[294];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_293_sv2v_reg <= w_data_i[293];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_292_sv2v_reg <= w_data_i[292];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_291_sv2v_reg <= w_data_i[291];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_290_sv2v_reg <= w_data_i[290];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_289_sv2v_reg <= w_data_i[289];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_288_sv2v_reg <= w_data_i[288];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_287_sv2v_reg <= w_data_i[287];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_286_sv2v_reg <= w_data_i[286];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_285_sv2v_reg <= w_data_i[285];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_284_sv2v_reg <= w_data_i[284];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_283_sv2v_reg <= w_data_i[283];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_282_sv2v_reg <= w_data_i[282];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_281_sv2v_reg <= w_data_i[281];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_280_sv2v_reg <= w_data_i[280];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_279_sv2v_reg <= w_data_i[279];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_278_sv2v_reg <= w_data_i[278];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_277_sv2v_reg <= w_data_i[277];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_276_sv2v_reg <= w_data_i[276];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_275_sv2v_reg <= w_data_i[275];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_274_sv2v_reg <= w_data_i[274];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_273_sv2v_reg <= w_data_i[273];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_272_sv2v_reg <= w_data_i[272];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_271_sv2v_reg <= w_data_i[271];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_270_sv2v_reg <= w_data_i[270];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_269_sv2v_reg <= w_data_i[269];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_268_sv2v_reg <= w_data_i[268];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_267_sv2v_reg <= w_data_i[267];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_266_sv2v_reg <= w_data_i[266];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_265_sv2v_reg <= w_data_i[265];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_264_sv2v_reg <= w_data_i[264];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_263_sv2v_reg <= w_data_i[263];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_262_sv2v_reg <= w_data_i[262];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_261_sv2v_reg <= w_data_i[261];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_260_sv2v_reg <= w_data_i[260];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_259_sv2v_reg <= w_data_i[259];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_258_sv2v_reg <= w_data_i[258];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_257_sv2v_reg <= w_data_i[257];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_256_sv2v_reg <= w_data_i[256];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_255_sv2v_reg <= w_data_i[255];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_254_sv2v_reg <= w_data_i[254];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_253_sv2v_reg <= w_data_i[253];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_252_sv2v_reg <= w_data_i[252];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_251_sv2v_reg <= w_data_i[251];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_250_sv2v_reg <= w_data_i[250];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_249_sv2v_reg <= w_data_i[249];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_248_sv2v_reg <= w_data_i[248];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_247_sv2v_reg <= w_data_i[247];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_246_sv2v_reg <= w_data_i[246];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_245_sv2v_reg <= w_data_i[245];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_244_sv2v_reg <= w_data_i[244];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_243_sv2v_reg <= w_data_i[243];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_242_sv2v_reg <= w_data_i[242];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_241_sv2v_reg <= w_data_i[241];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_240_sv2v_reg <= w_data_i[240];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_239_sv2v_reg <= w_data_i[239];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_238_sv2v_reg <= w_data_i[238];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_237_sv2v_reg <= w_data_i[237];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_236_sv2v_reg <= w_data_i[236];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_235_sv2v_reg <= w_data_i[235];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_234_sv2v_reg <= w_data_i[234];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_233_sv2v_reg <= w_data_i[233];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_232_sv2v_reg <= w_data_i[232];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_231_sv2v_reg <= w_data_i[231];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_230_sv2v_reg <= w_data_i[230];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_229_sv2v_reg <= w_data_i[229];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_228_sv2v_reg <= w_data_i[228];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_227_sv2v_reg <= w_data_i[227];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_226_sv2v_reg <= w_data_i[226];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_225_sv2v_reg <= w_data_i[225];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_224_sv2v_reg <= w_data_i[224];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_223_sv2v_reg <= w_data_i[223];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_222_sv2v_reg <= w_data_i[222];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_221_sv2v_reg <= w_data_i[221];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_220_sv2v_reg <= w_data_i[220];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_219_sv2v_reg <= w_data_i[219];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_218_sv2v_reg <= w_data_i[218];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_217_sv2v_reg <= w_data_i[217];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_216_sv2v_reg <= w_data_i[216];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_215_sv2v_reg <= w_data_i[215];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_214_sv2v_reg <= w_data_i[214];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_213_sv2v_reg <= w_data_i[213];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_212_sv2v_reg <= w_data_i[212];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_211_sv2v_reg <= w_data_i[211];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_210_sv2v_reg <= w_data_i[210];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_209_sv2v_reg <= w_data_i[209];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_208_sv2v_reg <= w_data_i[208];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_207_sv2v_reg <= w_data_i[207];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_206_sv2v_reg <= w_data_i[206];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_205_sv2v_reg <= w_data_i[205];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_204_sv2v_reg <= w_data_i[204];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_203_sv2v_reg <= w_data_i[203];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_202_sv2v_reg <= w_data_i[202];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_201_sv2v_reg <= w_data_i[201];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_200_sv2v_reg <= w_data_i[200];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_199_sv2v_reg <= w_data_i[199];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_198_sv2v_reg <= w_data_i[198];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_197_sv2v_reg <= w_data_i[197];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_196_sv2v_reg <= w_data_i[196];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_195_sv2v_reg <= w_data_i[195];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_194_sv2v_reg <= w_data_i[194];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_193_sv2v_reg <= w_data_i[193];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_192_sv2v_reg <= w_data_i[192];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_191_sv2v_reg <= w_data_i[191];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_190_sv2v_reg <= w_data_i[190];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_189_sv2v_reg <= w_data_i[189];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_188_sv2v_reg <= w_data_i[188];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_187_sv2v_reg <= w_data_i[187];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_186_sv2v_reg <= w_data_i[186];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_185_sv2v_reg <= w_data_i[185];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_184_sv2v_reg <= w_data_i[184];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_183_sv2v_reg <= w_data_i[183];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_182_sv2v_reg <= w_data_i[182];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_181_sv2v_reg <= w_data_i[181];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_180_sv2v_reg <= w_data_i[180];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_179_sv2v_reg <= w_data_i[179];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_178_sv2v_reg <= w_data_i[178];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_177_sv2v_reg <= w_data_i[177];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_176_sv2v_reg <= w_data_i[176];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_175_sv2v_reg <= w_data_i[175];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_174_sv2v_reg <= w_data_i[174];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_173_sv2v_reg <= w_data_i[173];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_172_sv2v_reg <= w_data_i[172];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_171_sv2v_reg <= w_data_i[171];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_170_sv2v_reg <= w_data_i[170];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_169_sv2v_reg <= w_data_i[169];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_168_sv2v_reg <= w_data_i[168];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_167_sv2v_reg <= w_data_i[167];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_166_sv2v_reg <= w_data_i[166];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_165_sv2v_reg <= w_data_i[165];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_164_sv2v_reg <= w_data_i[164];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_163_sv2v_reg <= w_data_i[163];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_162_sv2v_reg <= w_data_i[162];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_161_sv2v_reg <= w_data_i[161];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_160_sv2v_reg <= w_data_i[160];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_159_sv2v_reg <= w_data_i[159];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_158_sv2v_reg <= w_data_i[158];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_157_sv2v_reg <= w_data_i[157];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_156_sv2v_reg <= w_data_i[156];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_155_sv2v_reg <= w_data_i[155];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_154_sv2v_reg <= w_data_i[154];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_153_sv2v_reg <= w_data_i[153];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_152_sv2v_reg <= w_data_i[152];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_151_sv2v_reg <= w_data_i[151];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_150_sv2v_reg <= w_data_i[150];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_149_sv2v_reg <= w_data_i[149];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_148_sv2v_reg <= w_data_i[148];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_147_sv2v_reg <= w_data_i[147];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_146_sv2v_reg <= w_data_i[146];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_145_sv2v_reg <= w_data_i[145];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_144_sv2v_reg <= w_data_i[144];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_143_sv2v_reg <= w_data_i[143];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_142_sv2v_reg <= w_data_i[142];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_141_sv2v_reg <= w_data_i[141];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_140_sv2v_reg <= w_data_i[140];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_139_sv2v_reg <= w_data_i[139];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_138_sv2v_reg <= w_data_i[138];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_137_sv2v_reg <= w_data_i[137];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_136_sv2v_reg <= w_data_i[136];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_135_sv2v_reg <= w_data_i[135];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_134_sv2v_reg <= w_data_i[134];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_133_sv2v_reg <= w_data_i[133];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_132_sv2v_reg <= w_data_i[132];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_131_sv2v_reg <= w_data_i[131];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_130_sv2v_reg <= w_data_i[130];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_129_sv2v_reg <= w_data_i[129];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_128_sv2v_reg <= w_data_i[128];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_127_sv2v_reg <= w_data_i[127];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_126_sv2v_reg <= w_data_i[126];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_125_sv2v_reg <= w_data_i[125];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_124_sv2v_reg <= w_data_i[124];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_123_sv2v_reg <= w_data_i[123];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_122_sv2v_reg <= w_data_i[122];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_121_sv2v_reg <= w_data_i[121];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_120_sv2v_reg <= w_data_i[120];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_119_sv2v_reg <= w_data_i[119];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_118_sv2v_reg <= w_data_i[118];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_117_sv2v_reg <= w_data_i[117];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_116_sv2v_reg <= w_data_i[116];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_115_sv2v_reg <= w_data_i[115];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_114_sv2v_reg <= w_data_i[114];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_113_sv2v_reg <= w_data_i[113];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_112_sv2v_reg <= w_data_i[112];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_111_sv2v_reg <= w_data_i[111];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_110_sv2v_reg <= w_data_i[110];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_109_sv2v_reg <= w_data_i[109];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_108_sv2v_reg <= w_data_i[108];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_107_sv2v_reg <= w_data_i[107];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_106_sv2v_reg <= w_data_i[106];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_105_sv2v_reg <= w_data_i[105];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_104_sv2v_reg <= w_data_i[104];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_103_sv2v_reg <= w_data_i[103];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_102_sv2v_reg <= w_data_i[102];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_101_sv2v_reg <= w_data_i[101];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_100_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_99_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_98_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_97_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_96_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_95_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_94_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_93_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_92_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_91_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_90_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_89_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_88_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_87_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_86_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_85_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_84_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_83_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_82_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_81_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_80_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_79_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_78_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_77_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_76_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_75_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_74_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_73_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_72_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_71_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_70_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_69_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_68_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_67_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_66_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_65_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_64_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_63_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_62_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_61_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_60_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_59_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_58_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_57_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_56_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_55_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_54_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_53_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_52_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_51_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_50_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_49_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_48_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_47_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_46_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_45_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_44_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_43_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_42_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_41_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_40_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_39_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_38_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_37_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_36_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_35_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_34_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_33_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_32_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_31_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_30_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_29_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_28_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_27_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_26_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_25_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_24_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_23_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_22_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_21_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_20_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_19_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_18_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_17_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_16_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_15_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_14_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_13_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_12_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_11_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_10_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_9_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_8_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_7_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_6_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_5_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_4_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_3_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_2_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_1_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end

  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } : 
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

endmodule