module bsg_parallel_in_serial_out_width_p64_els_p8
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_i
);

  input [511:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input valid_i;
  input yumi_i;
  output ready_o;
  output valid_o;
  wire [63:0] data_o;
  wire ready_o,valid_o,N0,N1,piso_done_tx_n,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39;
  wire [2:0] piso_shift_ctr_r;
  wire [0:0] piso_state_n;
  wire [511:0] piso_data_r;
  reg valid_o_sv2v_reg,piso_data_r_511_sv2v_reg,piso_data_r_510_sv2v_reg,
  piso_data_r_509_sv2v_reg,piso_data_r_508_sv2v_reg,piso_data_r_507_sv2v_reg,
  piso_data_r_506_sv2v_reg,piso_data_r_505_sv2v_reg,piso_data_r_504_sv2v_reg,
  piso_data_r_503_sv2v_reg,piso_data_r_502_sv2v_reg,piso_data_r_501_sv2v_reg,piso_data_r_500_sv2v_reg,
  piso_data_r_499_sv2v_reg,piso_data_r_498_sv2v_reg,piso_data_r_497_sv2v_reg,
  piso_data_r_496_sv2v_reg,piso_data_r_495_sv2v_reg,piso_data_r_494_sv2v_reg,
  piso_data_r_493_sv2v_reg,piso_data_r_492_sv2v_reg,piso_data_r_491_sv2v_reg,
  piso_data_r_490_sv2v_reg,piso_data_r_489_sv2v_reg,piso_data_r_488_sv2v_reg,
  piso_data_r_487_sv2v_reg,piso_data_r_486_sv2v_reg,piso_data_r_485_sv2v_reg,piso_data_r_484_sv2v_reg,
  piso_data_r_483_sv2v_reg,piso_data_r_482_sv2v_reg,piso_data_r_481_sv2v_reg,
  piso_data_r_480_sv2v_reg,piso_data_r_479_sv2v_reg,piso_data_r_478_sv2v_reg,
  piso_data_r_477_sv2v_reg,piso_data_r_476_sv2v_reg,piso_data_r_475_sv2v_reg,
  piso_data_r_474_sv2v_reg,piso_data_r_473_sv2v_reg,piso_data_r_472_sv2v_reg,
  piso_data_r_471_sv2v_reg,piso_data_r_470_sv2v_reg,piso_data_r_469_sv2v_reg,piso_data_r_468_sv2v_reg,
  piso_data_r_467_sv2v_reg,piso_data_r_466_sv2v_reg,piso_data_r_465_sv2v_reg,
  piso_data_r_464_sv2v_reg,piso_data_r_463_sv2v_reg,piso_data_r_462_sv2v_reg,
  piso_data_r_461_sv2v_reg,piso_data_r_460_sv2v_reg,piso_data_r_459_sv2v_reg,
  piso_data_r_458_sv2v_reg,piso_data_r_457_sv2v_reg,piso_data_r_456_sv2v_reg,
  piso_data_r_455_sv2v_reg,piso_data_r_454_sv2v_reg,piso_data_r_453_sv2v_reg,piso_data_r_452_sv2v_reg,
  piso_data_r_451_sv2v_reg,piso_data_r_450_sv2v_reg,piso_data_r_449_sv2v_reg,
  piso_data_r_448_sv2v_reg,piso_data_r_447_sv2v_reg,piso_data_r_446_sv2v_reg,
  piso_data_r_445_sv2v_reg,piso_data_r_444_sv2v_reg,piso_data_r_443_sv2v_reg,
  piso_data_r_442_sv2v_reg,piso_data_r_441_sv2v_reg,piso_data_r_440_sv2v_reg,
  piso_data_r_439_sv2v_reg,piso_data_r_438_sv2v_reg,piso_data_r_437_sv2v_reg,piso_data_r_436_sv2v_reg,
  piso_data_r_435_sv2v_reg,piso_data_r_434_sv2v_reg,piso_data_r_433_sv2v_reg,
  piso_data_r_432_sv2v_reg,piso_data_r_431_sv2v_reg,piso_data_r_430_sv2v_reg,
  piso_data_r_429_sv2v_reg,piso_data_r_428_sv2v_reg,piso_data_r_427_sv2v_reg,
  piso_data_r_426_sv2v_reg,piso_data_r_425_sv2v_reg,piso_data_r_424_sv2v_reg,
  piso_data_r_423_sv2v_reg,piso_data_r_422_sv2v_reg,piso_data_r_421_sv2v_reg,piso_data_r_420_sv2v_reg,
  piso_data_r_419_sv2v_reg,piso_data_r_418_sv2v_reg,piso_data_r_417_sv2v_reg,
  piso_data_r_416_sv2v_reg,piso_data_r_415_sv2v_reg,piso_data_r_414_sv2v_reg,
  piso_data_r_413_sv2v_reg,piso_data_r_412_sv2v_reg,piso_data_r_411_sv2v_reg,
  piso_data_r_410_sv2v_reg,piso_data_r_409_sv2v_reg,piso_data_r_408_sv2v_reg,
  piso_data_r_407_sv2v_reg,piso_data_r_406_sv2v_reg,piso_data_r_405_sv2v_reg,piso_data_r_404_sv2v_reg,
  piso_data_r_403_sv2v_reg,piso_data_r_402_sv2v_reg,piso_data_r_401_sv2v_reg,
  piso_data_r_400_sv2v_reg,piso_data_r_399_sv2v_reg,piso_data_r_398_sv2v_reg,
  piso_data_r_397_sv2v_reg,piso_data_r_396_sv2v_reg,piso_data_r_395_sv2v_reg,
  piso_data_r_394_sv2v_reg,piso_data_r_393_sv2v_reg,piso_data_r_392_sv2v_reg,
  piso_data_r_391_sv2v_reg,piso_data_r_390_sv2v_reg,piso_data_r_389_sv2v_reg,piso_data_r_388_sv2v_reg,
  piso_data_r_387_sv2v_reg,piso_data_r_386_sv2v_reg,piso_data_r_385_sv2v_reg,
  piso_data_r_384_sv2v_reg,piso_data_r_383_sv2v_reg,piso_data_r_382_sv2v_reg,
  piso_data_r_381_sv2v_reg,piso_data_r_380_sv2v_reg,piso_data_r_379_sv2v_reg,
  piso_data_r_378_sv2v_reg,piso_data_r_377_sv2v_reg,piso_data_r_376_sv2v_reg,
  piso_data_r_375_sv2v_reg,piso_data_r_374_sv2v_reg,piso_data_r_373_sv2v_reg,piso_data_r_372_sv2v_reg,
  piso_data_r_371_sv2v_reg,piso_data_r_370_sv2v_reg,piso_data_r_369_sv2v_reg,
  piso_data_r_368_sv2v_reg,piso_data_r_367_sv2v_reg,piso_data_r_366_sv2v_reg,
  piso_data_r_365_sv2v_reg,piso_data_r_364_sv2v_reg,piso_data_r_363_sv2v_reg,
  piso_data_r_362_sv2v_reg,piso_data_r_361_sv2v_reg,piso_data_r_360_sv2v_reg,
  piso_data_r_359_sv2v_reg,piso_data_r_358_sv2v_reg,piso_data_r_357_sv2v_reg,piso_data_r_356_sv2v_reg,
  piso_data_r_355_sv2v_reg,piso_data_r_354_sv2v_reg,piso_data_r_353_sv2v_reg,
  piso_data_r_352_sv2v_reg,piso_data_r_351_sv2v_reg,piso_data_r_350_sv2v_reg,
  piso_data_r_349_sv2v_reg,piso_data_r_348_sv2v_reg,piso_data_r_347_sv2v_reg,
  piso_data_r_346_sv2v_reg,piso_data_r_345_sv2v_reg,piso_data_r_344_sv2v_reg,
  piso_data_r_343_sv2v_reg,piso_data_r_342_sv2v_reg,piso_data_r_341_sv2v_reg,piso_data_r_340_sv2v_reg,
  piso_data_r_339_sv2v_reg,piso_data_r_338_sv2v_reg,piso_data_r_337_sv2v_reg,
  piso_data_r_336_sv2v_reg,piso_data_r_335_sv2v_reg,piso_data_r_334_sv2v_reg,
  piso_data_r_333_sv2v_reg,piso_data_r_332_sv2v_reg,piso_data_r_331_sv2v_reg,
  piso_data_r_330_sv2v_reg,piso_data_r_329_sv2v_reg,piso_data_r_328_sv2v_reg,
  piso_data_r_327_sv2v_reg,piso_data_r_326_sv2v_reg,piso_data_r_325_sv2v_reg,piso_data_r_324_sv2v_reg,
  piso_data_r_323_sv2v_reg,piso_data_r_322_sv2v_reg,piso_data_r_321_sv2v_reg,
  piso_data_r_320_sv2v_reg,piso_data_r_319_sv2v_reg,piso_data_r_318_sv2v_reg,
  piso_data_r_317_sv2v_reg,piso_data_r_316_sv2v_reg,piso_data_r_315_sv2v_reg,
  piso_data_r_314_sv2v_reg,piso_data_r_313_sv2v_reg,piso_data_r_312_sv2v_reg,
  piso_data_r_311_sv2v_reg,piso_data_r_310_sv2v_reg,piso_data_r_309_sv2v_reg,piso_data_r_308_sv2v_reg,
  piso_data_r_307_sv2v_reg,piso_data_r_306_sv2v_reg,piso_data_r_305_sv2v_reg,
  piso_data_r_304_sv2v_reg,piso_data_r_303_sv2v_reg,piso_data_r_302_sv2v_reg,
  piso_data_r_301_sv2v_reg,piso_data_r_300_sv2v_reg,piso_data_r_299_sv2v_reg,
  piso_data_r_298_sv2v_reg,piso_data_r_297_sv2v_reg,piso_data_r_296_sv2v_reg,
  piso_data_r_295_sv2v_reg,piso_data_r_294_sv2v_reg,piso_data_r_293_sv2v_reg,piso_data_r_292_sv2v_reg,
  piso_data_r_291_sv2v_reg,piso_data_r_290_sv2v_reg,piso_data_r_289_sv2v_reg,
  piso_data_r_288_sv2v_reg,piso_data_r_287_sv2v_reg,piso_data_r_286_sv2v_reg,
  piso_data_r_285_sv2v_reg,piso_data_r_284_sv2v_reg,piso_data_r_283_sv2v_reg,
  piso_data_r_282_sv2v_reg,piso_data_r_281_sv2v_reg,piso_data_r_280_sv2v_reg,
  piso_data_r_279_sv2v_reg,piso_data_r_278_sv2v_reg,piso_data_r_277_sv2v_reg,piso_data_r_276_sv2v_reg,
  piso_data_r_275_sv2v_reg,piso_data_r_274_sv2v_reg,piso_data_r_273_sv2v_reg,
  piso_data_r_272_sv2v_reg,piso_data_r_271_sv2v_reg,piso_data_r_270_sv2v_reg,
  piso_data_r_269_sv2v_reg,piso_data_r_268_sv2v_reg,piso_data_r_267_sv2v_reg,
  piso_data_r_266_sv2v_reg,piso_data_r_265_sv2v_reg,piso_data_r_264_sv2v_reg,
  piso_data_r_263_sv2v_reg,piso_data_r_262_sv2v_reg,piso_data_r_261_sv2v_reg,piso_data_r_260_sv2v_reg,
  piso_data_r_259_sv2v_reg,piso_data_r_258_sv2v_reg,piso_data_r_257_sv2v_reg,
  piso_data_r_256_sv2v_reg,piso_data_r_255_sv2v_reg,piso_data_r_254_sv2v_reg,
  piso_data_r_253_sv2v_reg,piso_data_r_252_sv2v_reg,piso_data_r_251_sv2v_reg,
  piso_data_r_250_sv2v_reg,piso_data_r_249_sv2v_reg,piso_data_r_248_sv2v_reg,
  piso_data_r_247_sv2v_reg,piso_data_r_246_sv2v_reg,piso_data_r_245_sv2v_reg,piso_data_r_244_sv2v_reg,
  piso_data_r_243_sv2v_reg,piso_data_r_242_sv2v_reg,piso_data_r_241_sv2v_reg,
  piso_data_r_240_sv2v_reg,piso_data_r_239_sv2v_reg,piso_data_r_238_sv2v_reg,
  piso_data_r_237_sv2v_reg,piso_data_r_236_sv2v_reg,piso_data_r_235_sv2v_reg,
  piso_data_r_234_sv2v_reg,piso_data_r_233_sv2v_reg,piso_data_r_232_sv2v_reg,
  piso_data_r_231_sv2v_reg,piso_data_r_230_sv2v_reg,piso_data_r_229_sv2v_reg,piso_data_r_228_sv2v_reg,
  piso_data_r_227_sv2v_reg,piso_data_r_226_sv2v_reg,piso_data_r_225_sv2v_reg,
  piso_data_r_224_sv2v_reg,piso_data_r_223_sv2v_reg,piso_data_r_222_sv2v_reg,
  piso_data_r_221_sv2v_reg,piso_data_r_220_sv2v_reg,piso_data_r_219_sv2v_reg,
  piso_data_r_218_sv2v_reg,piso_data_r_217_sv2v_reg,piso_data_r_216_sv2v_reg,
  piso_data_r_215_sv2v_reg,piso_data_r_214_sv2v_reg,piso_data_r_213_sv2v_reg,piso_data_r_212_sv2v_reg,
  piso_data_r_211_sv2v_reg,piso_data_r_210_sv2v_reg,piso_data_r_209_sv2v_reg,
  piso_data_r_208_sv2v_reg,piso_data_r_207_sv2v_reg,piso_data_r_206_sv2v_reg,
  piso_data_r_205_sv2v_reg,piso_data_r_204_sv2v_reg,piso_data_r_203_sv2v_reg,
  piso_data_r_202_sv2v_reg,piso_data_r_201_sv2v_reg,piso_data_r_200_sv2v_reg,
  piso_data_r_199_sv2v_reg,piso_data_r_198_sv2v_reg,piso_data_r_197_sv2v_reg,piso_data_r_196_sv2v_reg,
  piso_data_r_195_sv2v_reg,piso_data_r_194_sv2v_reg,piso_data_r_193_sv2v_reg,
  piso_data_r_192_sv2v_reg,piso_data_r_191_sv2v_reg,piso_data_r_190_sv2v_reg,
  piso_data_r_189_sv2v_reg,piso_data_r_188_sv2v_reg,piso_data_r_187_sv2v_reg,
  piso_data_r_186_sv2v_reg,piso_data_r_185_sv2v_reg,piso_data_r_184_sv2v_reg,
  piso_data_r_183_sv2v_reg,piso_data_r_182_sv2v_reg,piso_data_r_181_sv2v_reg,piso_data_r_180_sv2v_reg,
  piso_data_r_179_sv2v_reg,piso_data_r_178_sv2v_reg,piso_data_r_177_sv2v_reg,
  piso_data_r_176_sv2v_reg,piso_data_r_175_sv2v_reg,piso_data_r_174_sv2v_reg,
  piso_data_r_173_sv2v_reg,piso_data_r_172_sv2v_reg,piso_data_r_171_sv2v_reg,
  piso_data_r_170_sv2v_reg,piso_data_r_169_sv2v_reg,piso_data_r_168_sv2v_reg,
  piso_data_r_167_sv2v_reg,piso_data_r_166_sv2v_reg,piso_data_r_165_sv2v_reg,piso_data_r_164_sv2v_reg,
  piso_data_r_163_sv2v_reg,piso_data_r_162_sv2v_reg,piso_data_r_161_sv2v_reg,
  piso_data_r_160_sv2v_reg,piso_data_r_159_sv2v_reg,piso_data_r_158_sv2v_reg,
  piso_data_r_157_sv2v_reg,piso_data_r_156_sv2v_reg,piso_data_r_155_sv2v_reg,
  piso_data_r_154_sv2v_reg,piso_data_r_153_sv2v_reg,piso_data_r_152_sv2v_reg,
  piso_data_r_151_sv2v_reg,piso_data_r_150_sv2v_reg,piso_data_r_149_sv2v_reg,piso_data_r_148_sv2v_reg,
  piso_data_r_147_sv2v_reg,piso_data_r_146_sv2v_reg,piso_data_r_145_sv2v_reg,
  piso_data_r_144_sv2v_reg,piso_data_r_143_sv2v_reg,piso_data_r_142_sv2v_reg,
  piso_data_r_141_sv2v_reg,piso_data_r_140_sv2v_reg,piso_data_r_139_sv2v_reg,
  piso_data_r_138_sv2v_reg,piso_data_r_137_sv2v_reg,piso_data_r_136_sv2v_reg,
  piso_data_r_135_sv2v_reg,piso_data_r_134_sv2v_reg,piso_data_r_133_sv2v_reg,piso_data_r_132_sv2v_reg,
  piso_data_r_131_sv2v_reg,piso_data_r_130_sv2v_reg,piso_data_r_129_sv2v_reg,
  piso_data_r_128_sv2v_reg,piso_data_r_127_sv2v_reg,piso_data_r_126_sv2v_reg,
  piso_data_r_125_sv2v_reg,piso_data_r_124_sv2v_reg,piso_data_r_123_sv2v_reg,
  piso_data_r_122_sv2v_reg,piso_data_r_121_sv2v_reg,piso_data_r_120_sv2v_reg,
  piso_data_r_119_sv2v_reg,piso_data_r_118_sv2v_reg,piso_data_r_117_sv2v_reg,piso_data_r_116_sv2v_reg,
  piso_data_r_115_sv2v_reg,piso_data_r_114_sv2v_reg,piso_data_r_113_sv2v_reg,
  piso_data_r_112_sv2v_reg,piso_data_r_111_sv2v_reg,piso_data_r_110_sv2v_reg,
  piso_data_r_109_sv2v_reg,piso_data_r_108_sv2v_reg,piso_data_r_107_sv2v_reg,
  piso_data_r_106_sv2v_reg,piso_data_r_105_sv2v_reg,piso_data_r_104_sv2v_reg,
  piso_data_r_103_sv2v_reg,piso_data_r_102_sv2v_reg,piso_data_r_101_sv2v_reg,piso_data_r_100_sv2v_reg,
  piso_data_r_99_sv2v_reg,piso_data_r_98_sv2v_reg,piso_data_r_97_sv2v_reg,
  piso_data_r_96_sv2v_reg,piso_data_r_95_sv2v_reg,piso_data_r_94_sv2v_reg,
  piso_data_r_93_sv2v_reg,piso_data_r_92_sv2v_reg,piso_data_r_91_sv2v_reg,piso_data_r_90_sv2v_reg,
  piso_data_r_89_sv2v_reg,piso_data_r_88_sv2v_reg,piso_data_r_87_sv2v_reg,
  piso_data_r_86_sv2v_reg,piso_data_r_85_sv2v_reg,piso_data_r_84_sv2v_reg,
  piso_data_r_83_sv2v_reg,piso_data_r_82_sv2v_reg,piso_data_r_81_sv2v_reg,piso_data_r_80_sv2v_reg,
  piso_data_r_79_sv2v_reg,piso_data_r_78_sv2v_reg,piso_data_r_77_sv2v_reg,
  piso_data_r_76_sv2v_reg,piso_data_r_75_sv2v_reg,piso_data_r_74_sv2v_reg,
  piso_data_r_73_sv2v_reg,piso_data_r_72_sv2v_reg,piso_data_r_71_sv2v_reg,piso_data_r_70_sv2v_reg,
  piso_data_r_69_sv2v_reg,piso_data_r_68_sv2v_reg,piso_data_r_67_sv2v_reg,
  piso_data_r_66_sv2v_reg,piso_data_r_65_sv2v_reg,piso_data_r_64_sv2v_reg,
  piso_data_r_63_sv2v_reg,piso_data_r_62_sv2v_reg,piso_data_r_61_sv2v_reg,piso_data_r_60_sv2v_reg,
  piso_data_r_59_sv2v_reg,piso_data_r_58_sv2v_reg,piso_data_r_57_sv2v_reg,
  piso_data_r_56_sv2v_reg,piso_data_r_55_sv2v_reg,piso_data_r_54_sv2v_reg,
  piso_data_r_53_sv2v_reg,piso_data_r_52_sv2v_reg,piso_data_r_51_sv2v_reg,piso_data_r_50_sv2v_reg,
  piso_data_r_49_sv2v_reg,piso_data_r_48_sv2v_reg,piso_data_r_47_sv2v_reg,
  piso_data_r_46_sv2v_reg,piso_data_r_45_sv2v_reg,piso_data_r_44_sv2v_reg,
  piso_data_r_43_sv2v_reg,piso_data_r_42_sv2v_reg,piso_data_r_41_sv2v_reg,piso_data_r_40_sv2v_reg,
  piso_data_r_39_sv2v_reg,piso_data_r_38_sv2v_reg,piso_data_r_37_sv2v_reg,
  piso_data_r_36_sv2v_reg,piso_data_r_35_sv2v_reg,piso_data_r_34_sv2v_reg,
  piso_data_r_33_sv2v_reg,piso_data_r_32_sv2v_reg,piso_data_r_31_sv2v_reg,piso_data_r_30_sv2v_reg,
  piso_data_r_29_sv2v_reg,piso_data_r_28_sv2v_reg,piso_data_r_27_sv2v_reg,
  piso_data_r_26_sv2v_reg,piso_data_r_25_sv2v_reg,piso_data_r_24_sv2v_reg,
  piso_data_r_23_sv2v_reg,piso_data_r_22_sv2v_reg,piso_data_r_21_sv2v_reg,piso_data_r_20_sv2v_reg,
  piso_data_r_19_sv2v_reg,piso_data_r_18_sv2v_reg,piso_data_r_17_sv2v_reg,
  piso_data_r_16_sv2v_reg,piso_data_r_15_sv2v_reg,piso_data_r_14_sv2v_reg,
  piso_data_r_13_sv2v_reg,piso_data_r_12_sv2v_reg,piso_data_r_11_sv2v_reg,piso_data_r_10_sv2v_reg,
  piso_data_r_9_sv2v_reg,piso_data_r_8_sv2v_reg,piso_data_r_7_sv2v_reg,
  piso_data_r_6_sv2v_reg,piso_data_r_5_sv2v_reg,piso_data_r_4_sv2v_reg,piso_data_r_3_sv2v_reg,
  piso_data_r_2_sv2v_reg,piso_data_r_1_sv2v_reg,piso_data_r_0_sv2v_reg,
  piso_shift_ctr_r_2_sv2v_reg,piso_shift_ctr_r_1_sv2v_reg,piso_shift_ctr_r_0_sv2v_reg;
  assign valid_o = valid_o_sv2v_reg;
  assign piso_data_r[511] = piso_data_r_511_sv2v_reg;
  assign piso_data_r[510] = piso_data_r_510_sv2v_reg;
  assign piso_data_r[509] = piso_data_r_509_sv2v_reg;
  assign piso_data_r[508] = piso_data_r_508_sv2v_reg;
  assign piso_data_r[507] = piso_data_r_507_sv2v_reg;
  assign piso_data_r[506] = piso_data_r_506_sv2v_reg;
  assign piso_data_r[505] = piso_data_r_505_sv2v_reg;
  assign piso_data_r[504] = piso_data_r_504_sv2v_reg;
  assign piso_data_r[503] = piso_data_r_503_sv2v_reg;
  assign piso_data_r[502] = piso_data_r_502_sv2v_reg;
  assign piso_data_r[501] = piso_data_r_501_sv2v_reg;
  assign piso_data_r[500] = piso_data_r_500_sv2v_reg;
  assign piso_data_r[499] = piso_data_r_499_sv2v_reg;
  assign piso_data_r[498] = piso_data_r_498_sv2v_reg;
  assign piso_data_r[497] = piso_data_r_497_sv2v_reg;
  assign piso_data_r[496] = piso_data_r_496_sv2v_reg;
  assign piso_data_r[495] = piso_data_r_495_sv2v_reg;
  assign piso_data_r[494] = piso_data_r_494_sv2v_reg;
  assign piso_data_r[493] = piso_data_r_493_sv2v_reg;
  assign piso_data_r[492] = piso_data_r_492_sv2v_reg;
  assign piso_data_r[491] = piso_data_r_491_sv2v_reg;
  assign piso_data_r[490] = piso_data_r_490_sv2v_reg;
  assign piso_data_r[489] = piso_data_r_489_sv2v_reg;
  assign piso_data_r[488] = piso_data_r_488_sv2v_reg;
  assign piso_data_r[487] = piso_data_r_487_sv2v_reg;
  assign piso_data_r[486] = piso_data_r_486_sv2v_reg;
  assign piso_data_r[485] = piso_data_r_485_sv2v_reg;
  assign piso_data_r[484] = piso_data_r_484_sv2v_reg;
  assign piso_data_r[483] = piso_data_r_483_sv2v_reg;
  assign piso_data_r[482] = piso_data_r_482_sv2v_reg;
  assign piso_data_r[481] = piso_data_r_481_sv2v_reg;
  assign piso_data_r[480] = piso_data_r_480_sv2v_reg;
  assign piso_data_r[479] = piso_data_r_479_sv2v_reg;
  assign piso_data_r[478] = piso_data_r_478_sv2v_reg;
  assign piso_data_r[477] = piso_data_r_477_sv2v_reg;
  assign piso_data_r[476] = piso_data_r_476_sv2v_reg;
  assign piso_data_r[475] = piso_data_r_475_sv2v_reg;
  assign piso_data_r[474] = piso_data_r_474_sv2v_reg;
  assign piso_data_r[473] = piso_data_r_473_sv2v_reg;
  assign piso_data_r[472] = piso_data_r_472_sv2v_reg;
  assign piso_data_r[471] = piso_data_r_471_sv2v_reg;
  assign piso_data_r[470] = piso_data_r_470_sv2v_reg;
  assign piso_data_r[469] = piso_data_r_469_sv2v_reg;
  assign piso_data_r[468] = piso_data_r_468_sv2v_reg;
  assign piso_data_r[467] = piso_data_r_467_sv2v_reg;
  assign piso_data_r[466] = piso_data_r_466_sv2v_reg;
  assign piso_data_r[465] = piso_data_r_465_sv2v_reg;
  assign piso_data_r[464] = piso_data_r_464_sv2v_reg;
  assign piso_data_r[463] = piso_data_r_463_sv2v_reg;
  assign piso_data_r[462] = piso_data_r_462_sv2v_reg;
  assign piso_data_r[461] = piso_data_r_461_sv2v_reg;
  assign piso_data_r[460] = piso_data_r_460_sv2v_reg;
  assign piso_data_r[459] = piso_data_r_459_sv2v_reg;
  assign piso_data_r[458] = piso_data_r_458_sv2v_reg;
  assign piso_data_r[457] = piso_data_r_457_sv2v_reg;
  assign piso_data_r[456] = piso_data_r_456_sv2v_reg;
  assign piso_data_r[455] = piso_data_r_455_sv2v_reg;
  assign piso_data_r[454] = piso_data_r_454_sv2v_reg;
  assign piso_data_r[453] = piso_data_r_453_sv2v_reg;
  assign piso_data_r[452] = piso_data_r_452_sv2v_reg;
  assign piso_data_r[451] = piso_data_r_451_sv2v_reg;
  assign piso_data_r[450] = piso_data_r_450_sv2v_reg;
  assign piso_data_r[449] = piso_data_r_449_sv2v_reg;
  assign piso_data_r[448] = piso_data_r_448_sv2v_reg;
  assign piso_data_r[447] = piso_data_r_447_sv2v_reg;
  assign piso_data_r[446] = piso_data_r_446_sv2v_reg;
  assign piso_data_r[445] = piso_data_r_445_sv2v_reg;
  assign piso_data_r[444] = piso_data_r_444_sv2v_reg;
  assign piso_data_r[443] = piso_data_r_443_sv2v_reg;
  assign piso_data_r[442] = piso_data_r_442_sv2v_reg;
  assign piso_data_r[441] = piso_data_r_441_sv2v_reg;
  assign piso_data_r[440] = piso_data_r_440_sv2v_reg;
  assign piso_data_r[439] = piso_data_r_439_sv2v_reg;
  assign piso_data_r[438] = piso_data_r_438_sv2v_reg;
  assign piso_data_r[437] = piso_data_r_437_sv2v_reg;
  assign piso_data_r[436] = piso_data_r_436_sv2v_reg;
  assign piso_data_r[435] = piso_data_r_435_sv2v_reg;
  assign piso_data_r[434] = piso_data_r_434_sv2v_reg;
  assign piso_data_r[433] = piso_data_r_433_sv2v_reg;
  assign piso_data_r[432] = piso_data_r_432_sv2v_reg;
  assign piso_data_r[431] = piso_data_r_431_sv2v_reg;
  assign piso_data_r[430] = piso_data_r_430_sv2v_reg;
  assign piso_data_r[429] = piso_data_r_429_sv2v_reg;
  assign piso_data_r[428] = piso_data_r_428_sv2v_reg;
  assign piso_data_r[427] = piso_data_r_427_sv2v_reg;
  assign piso_data_r[426] = piso_data_r_426_sv2v_reg;
  assign piso_data_r[425] = piso_data_r_425_sv2v_reg;
  assign piso_data_r[424] = piso_data_r_424_sv2v_reg;
  assign piso_data_r[423] = piso_data_r_423_sv2v_reg;
  assign piso_data_r[422] = piso_data_r_422_sv2v_reg;
  assign piso_data_r[421] = piso_data_r_421_sv2v_reg;
  assign piso_data_r[420] = piso_data_r_420_sv2v_reg;
  assign piso_data_r[419] = piso_data_r_419_sv2v_reg;
  assign piso_data_r[418] = piso_data_r_418_sv2v_reg;
  assign piso_data_r[417] = piso_data_r_417_sv2v_reg;
  assign piso_data_r[416] = piso_data_r_416_sv2v_reg;
  assign piso_data_r[415] = piso_data_r_415_sv2v_reg;
  assign piso_data_r[414] = piso_data_r_414_sv2v_reg;
  assign piso_data_r[413] = piso_data_r_413_sv2v_reg;
  assign piso_data_r[412] = piso_data_r_412_sv2v_reg;
  assign piso_data_r[411] = piso_data_r_411_sv2v_reg;
  assign piso_data_r[410] = piso_data_r_410_sv2v_reg;
  assign piso_data_r[409] = piso_data_r_409_sv2v_reg;
  assign piso_data_r[408] = piso_data_r_408_sv2v_reg;
  assign piso_data_r[407] = piso_data_r_407_sv2v_reg;
  assign piso_data_r[406] = piso_data_r_406_sv2v_reg;
  assign piso_data_r[405] = piso_data_r_405_sv2v_reg;
  assign piso_data_r[404] = piso_data_r_404_sv2v_reg;
  assign piso_data_r[403] = piso_data_r_403_sv2v_reg;
  assign piso_data_r[402] = piso_data_r_402_sv2v_reg;
  assign piso_data_r[401] = piso_data_r_401_sv2v_reg;
  assign piso_data_r[400] = piso_data_r_400_sv2v_reg;
  assign piso_data_r[399] = piso_data_r_399_sv2v_reg;
  assign piso_data_r[398] = piso_data_r_398_sv2v_reg;
  assign piso_data_r[397] = piso_data_r_397_sv2v_reg;
  assign piso_data_r[396] = piso_data_r_396_sv2v_reg;
  assign piso_data_r[395] = piso_data_r_395_sv2v_reg;
  assign piso_data_r[394] = piso_data_r_394_sv2v_reg;
  assign piso_data_r[393] = piso_data_r_393_sv2v_reg;
  assign piso_data_r[392] = piso_data_r_392_sv2v_reg;
  assign piso_data_r[391] = piso_data_r_391_sv2v_reg;
  assign piso_data_r[390] = piso_data_r_390_sv2v_reg;
  assign piso_data_r[389] = piso_data_r_389_sv2v_reg;
  assign piso_data_r[388] = piso_data_r_388_sv2v_reg;
  assign piso_data_r[387] = piso_data_r_387_sv2v_reg;
  assign piso_data_r[386] = piso_data_r_386_sv2v_reg;
  assign piso_data_r[385] = piso_data_r_385_sv2v_reg;
  assign piso_data_r[384] = piso_data_r_384_sv2v_reg;
  assign piso_data_r[383] = piso_data_r_383_sv2v_reg;
  assign piso_data_r[382] = piso_data_r_382_sv2v_reg;
  assign piso_data_r[381] = piso_data_r_381_sv2v_reg;
  assign piso_data_r[380] = piso_data_r_380_sv2v_reg;
  assign piso_data_r[379] = piso_data_r_379_sv2v_reg;
  assign piso_data_r[378] = piso_data_r_378_sv2v_reg;
  assign piso_data_r[377] = piso_data_r_377_sv2v_reg;
  assign piso_data_r[376] = piso_data_r_376_sv2v_reg;
  assign piso_data_r[375] = piso_data_r_375_sv2v_reg;
  assign piso_data_r[374] = piso_data_r_374_sv2v_reg;
  assign piso_data_r[373] = piso_data_r_373_sv2v_reg;
  assign piso_data_r[372] = piso_data_r_372_sv2v_reg;
  assign piso_data_r[371] = piso_data_r_371_sv2v_reg;
  assign piso_data_r[370] = piso_data_r_370_sv2v_reg;
  assign piso_data_r[369] = piso_data_r_369_sv2v_reg;
  assign piso_data_r[368] = piso_data_r_368_sv2v_reg;
  assign piso_data_r[367] = piso_data_r_367_sv2v_reg;
  assign piso_data_r[366] = piso_data_r_366_sv2v_reg;
  assign piso_data_r[365] = piso_data_r_365_sv2v_reg;
  assign piso_data_r[364] = piso_data_r_364_sv2v_reg;
  assign piso_data_r[363] = piso_data_r_363_sv2v_reg;
  assign piso_data_r[362] = piso_data_r_362_sv2v_reg;
  assign piso_data_r[361] = piso_data_r_361_sv2v_reg;
  assign piso_data_r[360] = piso_data_r_360_sv2v_reg;
  assign piso_data_r[359] = piso_data_r_359_sv2v_reg;
  assign piso_data_r[358] = piso_data_r_358_sv2v_reg;
  assign piso_data_r[357] = piso_data_r_357_sv2v_reg;
  assign piso_data_r[356] = piso_data_r_356_sv2v_reg;
  assign piso_data_r[355] = piso_data_r_355_sv2v_reg;
  assign piso_data_r[354] = piso_data_r_354_sv2v_reg;
  assign piso_data_r[353] = piso_data_r_353_sv2v_reg;
  assign piso_data_r[352] = piso_data_r_352_sv2v_reg;
  assign piso_data_r[351] = piso_data_r_351_sv2v_reg;
  assign piso_data_r[350] = piso_data_r_350_sv2v_reg;
  assign piso_data_r[349] = piso_data_r_349_sv2v_reg;
  assign piso_data_r[348] = piso_data_r_348_sv2v_reg;
  assign piso_data_r[347] = piso_data_r_347_sv2v_reg;
  assign piso_data_r[346] = piso_data_r_346_sv2v_reg;
  assign piso_data_r[345] = piso_data_r_345_sv2v_reg;
  assign piso_data_r[344] = piso_data_r_344_sv2v_reg;
  assign piso_data_r[343] = piso_data_r_343_sv2v_reg;
  assign piso_data_r[342] = piso_data_r_342_sv2v_reg;
  assign piso_data_r[341] = piso_data_r_341_sv2v_reg;
  assign piso_data_r[340] = piso_data_r_340_sv2v_reg;
  assign piso_data_r[339] = piso_data_r_339_sv2v_reg;
  assign piso_data_r[338] = piso_data_r_338_sv2v_reg;
  assign piso_data_r[337] = piso_data_r_337_sv2v_reg;
  assign piso_data_r[336] = piso_data_r_336_sv2v_reg;
  assign piso_data_r[335] = piso_data_r_335_sv2v_reg;
  assign piso_data_r[334] = piso_data_r_334_sv2v_reg;
  assign piso_data_r[333] = piso_data_r_333_sv2v_reg;
  assign piso_data_r[332] = piso_data_r_332_sv2v_reg;
  assign piso_data_r[331] = piso_data_r_331_sv2v_reg;
  assign piso_data_r[330] = piso_data_r_330_sv2v_reg;
  assign piso_data_r[329] = piso_data_r_329_sv2v_reg;
  assign piso_data_r[328] = piso_data_r_328_sv2v_reg;
  assign piso_data_r[327] = piso_data_r_327_sv2v_reg;
  assign piso_data_r[326] = piso_data_r_326_sv2v_reg;
  assign piso_data_r[325] = piso_data_r_325_sv2v_reg;
  assign piso_data_r[324] = piso_data_r_324_sv2v_reg;
  assign piso_data_r[323] = piso_data_r_323_sv2v_reg;
  assign piso_data_r[322] = piso_data_r_322_sv2v_reg;
  assign piso_data_r[321] = piso_data_r_321_sv2v_reg;
  assign piso_data_r[320] = piso_data_r_320_sv2v_reg;
  assign piso_data_r[319] = piso_data_r_319_sv2v_reg;
  assign piso_data_r[318] = piso_data_r_318_sv2v_reg;
  assign piso_data_r[317] = piso_data_r_317_sv2v_reg;
  assign piso_data_r[316] = piso_data_r_316_sv2v_reg;
  assign piso_data_r[315] = piso_data_r_315_sv2v_reg;
  assign piso_data_r[314] = piso_data_r_314_sv2v_reg;
  assign piso_data_r[313] = piso_data_r_313_sv2v_reg;
  assign piso_data_r[312] = piso_data_r_312_sv2v_reg;
  assign piso_data_r[311] = piso_data_r_311_sv2v_reg;
  assign piso_data_r[310] = piso_data_r_310_sv2v_reg;
  assign piso_data_r[309] = piso_data_r_309_sv2v_reg;
  assign piso_data_r[308] = piso_data_r_308_sv2v_reg;
  assign piso_data_r[307] = piso_data_r_307_sv2v_reg;
  assign piso_data_r[306] = piso_data_r_306_sv2v_reg;
  assign piso_data_r[305] = piso_data_r_305_sv2v_reg;
  assign piso_data_r[304] = piso_data_r_304_sv2v_reg;
  assign piso_data_r[303] = piso_data_r_303_sv2v_reg;
  assign piso_data_r[302] = piso_data_r_302_sv2v_reg;
  assign piso_data_r[301] = piso_data_r_301_sv2v_reg;
  assign piso_data_r[300] = piso_data_r_300_sv2v_reg;
  assign piso_data_r[299] = piso_data_r_299_sv2v_reg;
  assign piso_data_r[298] = piso_data_r_298_sv2v_reg;
  assign piso_data_r[297] = piso_data_r_297_sv2v_reg;
  assign piso_data_r[296] = piso_data_r_296_sv2v_reg;
  assign piso_data_r[295] = piso_data_r_295_sv2v_reg;
  assign piso_data_r[294] = piso_data_r_294_sv2v_reg;
  assign piso_data_r[293] = piso_data_r_293_sv2v_reg;
  assign piso_data_r[292] = piso_data_r_292_sv2v_reg;
  assign piso_data_r[291] = piso_data_r_291_sv2v_reg;
  assign piso_data_r[290] = piso_data_r_290_sv2v_reg;
  assign piso_data_r[289] = piso_data_r_289_sv2v_reg;
  assign piso_data_r[288] = piso_data_r_288_sv2v_reg;
  assign piso_data_r[287] = piso_data_r_287_sv2v_reg;
  assign piso_data_r[286] = piso_data_r_286_sv2v_reg;
  assign piso_data_r[285] = piso_data_r_285_sv2v_reg;
  assign piso_data_r[284] = piso_data_r_284_sv2v_reg;
  assign piso_data_r[283] = piso_data_r_283_sv2v_reg;
  assign piso_data_r[282] = piso_data_r_282_sv2v_reg;
  assign piso_data_r[281] = piso_data_r_281_sv2v_reg;
  assign piso_data_r[280] = piso_data_r_280_sv2v_reg;
  assign piso_data_r[279] = piso_data_r_279_sv2v_reg;
  assign piso_data_r[278] = piso_data_r_278_sv2v_reg;
  assign piso_data_r[277] = piso_data_r_277_sv2v_reg;
  assign piso_data_r[276] = piso_data_r_276_sv2v_reg;
  assign piso_data_r[275] = piso_data_r_275_sv2v_reg;
  assign piso_data_r[274] = piso_data_r_274_sv2v_reg;
  assign piso_data_r[273] = piso_data_r_273_sv2v_reg;
  assign piso_data_r[272] = piso_data_r_272_sv2v_reg;
  assign piso_data_r[271] = piso_data_r_271_sv2v_reg;
  assign piso_data_r[270] = piso_data_r_270_sv2v_reg;
  assign piso_data_r[269] = piso_data_r_269_sv2v_reg;
  assign piso_data_r[268] = piso_data_r_268_sv2v_reg;
  assign piso_data_r[267] = piso_data_r_267_sv2v_reg;
  assign piso_data_r[266] = piso_data_r_266_sv2v_reg;
  assign piso_data_r[265] = piso_data_r_265_sv2v_reg;
  assign piso_data_r[264] = piso_data_r_264_sv2v_reg;
  assign piso_data_r[263] = piso_data_r_263_sv2v_reg;
  assign piso_data_r[262] = piso_data_r_262_sv2v_reg;
  assign piso_data_r[261] = piso_data_r_261_sv2v_reg;
  assign piso_data_r[260] = piso_data_r_260_sv2v_reg;
  assign piso_data_r[259] = piso_data_r_259_sv2v_reg;
  assign piso_data_r[258] = piso_data_r_258_sv2v_reg;
  assign piso_data_r[257] = piso_data_r_257_sv2v_reg;
  assign piso_data_r[256] = piso_data_r_256_sv2v_reg;
  assign piso_data_r[255] = piso_data_r_255_sv2v_reg;
  assign piso_data_r[254] = piso_data_r_254_sv2v_reg;
  assign piso_data_r[253] = piso_data_r_253_sv2v_reg;
  assign piso_data_r[252] = piso_data_r_252_sv2v_reg;
  assign piso_data_r[251] = piso_data_r_251_sv2v_reg;
  assign piso_data_r[250] = piso_data_r_250_sv2v_reg;
  assign piso_data_r[249] = piso_data_r_249_sv2v_reg;
  assign piso_data_r[248] = piso_data_r_248_sv2v_reg;
  assign piso_data_r[247] = piso_data_r_247_sv2v_reg;
  assign piso_data_r[246] = piso_data_r_246_sv2v_reg;
  assign piso_data_r[245] = piso_data_r_245_sv2v_reg;
  assign piso_data_r[244] = piso_data_r_244_sv2v_reg;
  assign piso_data_r[243] = piso_data_r_243_sv2v_reg;
  assign piso_data_r[242] = piso_data_r_242_sv2v_reg;
  assign piso_data_r[241] = piso_data_r_241_sv2v_reg;
  assign piso_data_r[240] = piso_data_r_240_sv2v_reg;
  assign piso_data_r[239] = piso_data_r_239_sv2v_reg;
  assign piso_data_r[238] = piso_data_r_238_sv2v_reg;
  assign piso_data_r[237] = piso_data_r_237_sv2v_reg;
  assign piso_data_r[236] = piso_data_r_236_sv2v_reg;
  assign piso_data_r[235] = piso_data_r_235_sv2v_reg;
  assign piso_data_r[234] = piso_data_r_234_sv2v_reg;
  assign piso_data_r[233] = piso_data_r_233_sv2v_reg;
  assign piso_data_r[232] = piso_data_r_232_sv2v_reg;
  assign piso_data_r[231] = piso_data_r_231_sv2v_reg;
  assign piso_data_r[230] = piso_data_r_230_sv2v_reg;
  assign piso_data_r[229] = piso_data_r_229_sv2v_reg;
  assign piso_data_r[228] = piso_data_r_228_sv2v_reg;
  assign piso_data_r[227] = piso_data_r_227_sv2v_reg;
  assign piso_data_r[226] = piso_data_r_226_sv2v_reg;
  assign piso_data_r[225] = piso_data_r_225_sv2v_reg;
  assign piso_data_r[224] = piso_data_r_224_sv2v_reg;
  assign piso_data_r[223] = piso_data_r_223_sv2v_reg;
  assign piso_data_r[222] = piso_data_r_222_sv2v_reg;
  assign piso_data_r[221] = piso_data_r_221_sv2v_reg;
  assign piso_data_r[220] = piso_data_r_220_sv2v_reg;
  assign piso_data_r[219] = piso_data_r_219_sv2v_reg;
  assign piso_data_r[218] = piso_data_r_218_sv2v_reg;
  assign piso_data_r[217] = piso_data_r_217_sv2v_reg;
  assign piso_data_r[216] = piso_data_r_216_sv2v_reg;
  assign piso_data_r[215] = piso_data_r_215_sv2v_reg;
  assign piso_data_r[214] = piso_data_r_214_sv2v_reg;
  assign piso_data_r[213] = piso_data_r_213_sv2v_reg;
  assign piso_data_r[212] = piso_data_r_212_sv2v_reg;
  assign piso_data_r[211] = piso_data_r_211_sv2v_reg;
  assign piso_data_r[210] = piso_data_r_210_sv2v_reg;
  assign piso_data_r[209] = piso_data_r_209_sv2v_reg;
  assign piso_data_r[208] = piso_data_r_208_sv2v_reg;
  assign piso_data_r[207] = piso_data_r_207_sv2v_reg;
  assign piso_data_r[206] = piso_data_r_206_sv2v_reg;
  assign piso_data_r[205] = piso_data_r_205_sv2v_reg;
  assign piso_data_r[204] = piso_data_r_204_sv2v_reg;
  assign piso_data_r[203] = piso_data_r_203_sv2v_reg;
  assign piso_data_r[202] = piso_data_r_202_sv2v_reg;
  assign piso_data_r[201] = piso_data_r_201_sv2v_reg;
  assign piso_data_r[200] = piso_data_r_200_sv2v_reg;
  assign piso_data_r[199] = piso_data_r_199_sv2v_reg;
  assign piso_data_r[198] = piso_data_r_198_sv2v_reg;
  assign piso_data_r[197] = piso_data_r_197_sv2v_reg;
  assign piso_data_r[196] = piso_data_r_196_sv2v_reg;
  assign piso_data_r[195] = piso_data_r_195_sv2v_reg;
  assign piso_data_r[194] = piso_data_r_194_sv2v_reg;
  assign piso_data_r[193] = piso_data_r_193_sv2v_reg;
  assign piso_data_r[192] = piso_data_r_192_sv2v_reg;
  assign piso_data_r[191] = piso_data_r_191_sv2v_reg;
  assign piso_data_r[190] = piso_data_r_190_sv2v_reg;
  assign piso_data_r[189] = piso_data_r_189_sv2v_reg;
  assign piso_data_r[188] = piso_data_r_188_sv2v_reg;
  assign piso_data_r[187] = piso_data_r_187_sv2v_reg;
  assign piso_data_r[186] = piso_data_r_186_sv2v_reg;
  assign piso_data_r[185] = piso_data_r_185_sv2v_reg;
  assign piso_data_r[184] = piso_data_r_184_sv2v_reg;
  assign piso_data_r[183] = piso_data_r_183_sv2v_reg;
  assign piso_data_r[182] = piso_data_r_182_sv2v_reg;
  assign piso_data_r[181] = piso_data_r_181_sv2v_reg;
  assign piso_data_r[180] = piso_data_r_180_sv2v_reg;
  assign piso_data_r[179] = piso_data_r_179_sv2v_reg;
  assign piso_data_r[178] = piso_data_r_178_sv2v_reg;
  assign piso_data_r[177] = piso_data_r_177_sv2v_reg;
  assign piso_data_r[176] = piso_data_r_176_sv2v_reg;
  assign piso_data_r[175] = piso_data_r_175_sv2v_reg;
  assign piso_data_r[174] = piso_data_r_174_sv2v_reg;
  assign piso_data_r[173] = piso_data_r_173_sv2v_reg;
  assign piso_data_r[172] = piso_data_r_172_sv2v_reg;
  assign piso_data_r[171] = piso_data_r_171_sv2v_reg;
  assign piso_data_r[170] = piso_data_r_170_sv2v_reg;
  assign piso_data_r[169] = piso_data_r_169_sv2v_reg;
  assign piso_data_r[168] = piso_data_r_168_sv2v_reg;
  assign piso_data_r[167] = piso_data_r_167_sv2v_reg;
  assign piso_data_r[166] = piso_data_r_166_sv2v_reg;
  assign piso_data_r[165] = piso_data_r_165_sv2v_reg;
  assign piso_data_r[164] = piso_data_r_164_sv2v_reg;
  assign piso_data_r[163] = piso_data_r_163_sv2v_reg;
  assign piso_data_r[162] = piso_data_r_162_sv2v_reg;
  assign piso_data_r[161] = piso_data_r_161_sv2v_reg;
  assign piso_data_r[160] = piso_data_r_160_sv2v_reg;
  assign piso_data_r[159] = piso_data_r_159_sv2v_reg;
  assign piso_data_r[158] = piso_data_r_158_sv2v_reg;
  assign piso_data_r[157] = piso_data_r_157_sv2v_reg;
  assign piso_data_r[156] = piso_data_r_156_sv2v_reg;
  assign piso_data_r[155] = piso_data_r_155_sv2v_reg;
  assign piso_data_r[154] = piso_data_r_154_sv2v_reg;
  assign piso_data_r[153] = piso_data_r_153_sv2v_reg;
  assign piso_data_r[152] = piso_data_r_152_sv2v_reg;
  assign piso_data_r[151] = piso_data_r_151_sv2v_reg;
  assign piso_data_r[150] = piso_data_r_150_sv2v_reg;
  assign piso_data_r[149] = piso_data_r_149_sv2v_reg;
  assign piso_data_r[148] = piso_data_r_148_sv2v_reg;
  assign piso_data_r[147] = piso_data_r_147_sv2v_reg;
  assign piso_data_r[146] = piso_data_r_146_sv2v_reg;
  assign piso_data_r[145] = piso_data_r_145_sv2v_reg;
  assign piso_data_r[144] = piso_data_r_144_sv2v_reg;
  assign piso_data_r[143] = piso_data_r_143_sv2v_reg;
  assign piso_data_r[142] = piso_data_r_142_sv2v_reg;
  assign piso_data_r[141] = piso_data_r_141_sv2v_reg;
  assign piso_data_r[140] = piso_data_r_140_sv2v_reg;
  assign piso_data_r[139] = piso_data_r_139_sv2v_reg;
  assign piso_data_r[138] = piso_data_r_138_sv2v_reg;
  assign piso_data_r[137] = piso_data_r_137_sv2v_reg;
  assign piso_data_r[136] = piso_data_r_136_sv2v_reg;
  assign piso_data_r[135] = piso_data_r_135_sv2v_reg;
  assign piso_data_r[134] = piso_data_r_134_sv2v_reg;
  assign piso_data_r[133] = piso_data_r_133_sv2v_reg;
  assign piso_data_r[132] = piso_data_r_132_sv2v_reg;
  assign piso_data_r[131] = piso_data_r_131_sv2v_reg;
  assign piso_data_r[130] = piso_data_r_130_sv2v_reg;
  assign piso_data_r[129] = piso_data_r_129_sv2v_reg;
  assign piso_data_r[128] = piso_data_r_128_sv2v_reg;
  assign piso_data_r[127] = piso_data_r_127_sv2v_reg;
  assign piso_data_r[126] = piso_data_r_126_sv2v_reg;
  assign piso_data_r[125] = piso_data_r_125_sv2v_reg;
  assign piso_data_r[124] = piso_data_r_124_sv2v_reg;
  assign piso_data_r[123] = piso_data_r_123_sv2v_reg;
  assign piso_data_r[122] = piso_data_r_122_sv2v_reg;
  assign piso_data_r[121] = piso_data_r_121_sv2v_reg;
  assign piso_data_r[120] = piso_data_r_120_sv2v_reg;
  assign piso_data_r[119] = piso_data_r_119_sv2v_reg;
  assign piso_data_r[118] = piso_data_r_118_sv2v_reg;
  assign piso_data_r[117] = piso_data_r_117_sv2v_reg;
  assign piso_data_r[116] = piso_data_r_116_sv2v_reg;
  assign piso_data_r[115] = piso_data_r_115_sv2v_reg;
  assign piso_data_r[114] = piso_data_r_114_sv2v_reg;
  assign piso_data_r[113] = piso_data_r_113_sv2v_reg;
  assign piso_data_r[112] = piso_data_r_112_sv2v_reg;
  assign piso_data_r[111] = piso_data_r_111_sv2v_reg;
  assign piso_data_r[110] = piso_data_r_110_sv2v_reg;
  assign piso_data_r[109] = piso_data_r_109_sv2v_reg;
  assign piso_data_r[108] = piso_data_r_108_sv2v_reg;
  assign piso_data_r[107] = piso_data_r_107_sv2v_reg;
  assign piso_data_r[106] = piso_data_r_106_sv2v_reg;
  assign piso_data_r[105] = piso_data_r_105_sv2v_reg;
  assign piso_data_r[104] = piso_data_r_104_sv2v_reg;
  assign piso_data_r[103] = piso_data_r_103_sv2v_reg;
  assign piso_data_r[102] = piso_data_r_102_sv2v_reg;
  assign piso_data_r[101] = piso_data_r_101_sv2v_reg;
  assign piso_data_r[100] = piso_data_r_100_sv2v_reg;
  assign piso_data_r[99] = piso_data_r_99_sv2v_reg;
  assign piso_data_r[98] = piso_data_r_98_sv2v_reg;
  assign piso_data_r[97] = piso_data_r_97_sv2v_reg;
  assign piso_data_r[96] = piso_data_r_96_sv2v_reg;
  assign piso_data_r[95] = piso_data_r_95_sv2v_reg;
  assign piso_data_r[94] = piso_data_r_94_sv2v_reg;
  assign piso_data_r[93] = piso_data_r_93_sv2v_reg;
  assign piso_data_r[92] = piso_data_r_92_sv2v_reg;
  assign piso_data_r[91] = piso_data_r_91_sv2v_reg;
  assign piso_data_r[90] = piso_data_r_90_sv2v_reg;
  assign piso_data_r[89] = piso_data_r_89_sv2v_reg;
  assign piso_data_r[88] = piso_data_r_88_sv2v_reg;
  assign piso_data_r[87] = piso_data_r_87_sv2v_reg;
  assign piso_data_r[86] = piso_data_r_86_sv2v_reg;
  assign piso_data_r[85] = piso_data_r_85_sv2v_reg;
  assign piso_data_r[84] = piso_data_r_84_sv2v_reg;
  assign piso_data_r[83] = piso_data_r_83_sv2v_reg;
  assign piso_data_r[82] = piso_data_r_82_sv2v_reg;
  assign piso_data_r[81] = piso_data_r_81_sv2v_reg;
  assign piso_data_r[80] = piso_data_r_80_sv2v_reg;
  assign piso_data_r[79] = piso_data_r_79_sv2v_reg;
  assign piso_data_r[78] = piso_data_r_78_sv2v_reg;
  assign piso_data_r[77] = piso_data_r_77_sv2v_reg;
  assign piso_data_r[76] = piso_data_r_76_sv2v_reg;
  assign piso_data_r[75] = piso_data_r_75_sv2v_reg;
  assign piso_data_r[74] = piso_data_r_74_sv2v_reg;
  assign piso_data_r[73] = piso_data_r_73_sv2v_reg;
  assign piso_data_r[72] = piso_data_r_72_sv2v_reg;
  assign piso_data_r[71] = piso_data_r_71_sv2v_reg;
  assign piso_data_r[70] = piso_data_r_70_sv2v_reg;
  assign piso_data_r[69] = piso_data_r_69_sv2v_reg;
  assign piso_data_r[68] = piso_data_r_68_sv2v_reg;
  assign piso_data_r[67] = piso_data_r_67_sv2v_reg;
  assign piso_data_r[66] = piso_data_r_66_sv2v_reg;
  assign piso_data_r[65] = piso_data_r_65_sv2v_reg;
  assign piso_data_r[64] = piso_data_r_64_sv2v_reg;
  assign piso_data_r[63] = piso_data_r_63_sv2v_reg;
  assign piso_data_r[62] = piso_data_r_62_sv2v_reg;
  assign piso_data_r[61] = piso_data_r_61_sv2v_reg;
  assign piso_data_r[60] = piso_data_r_60_sv2v_reg;
  assign piso_data_r[59] = piso_data_r_59_sv2v_reg;
  assign piso_data_r[58] = piso_data_r_58_sv2v_reg;
  assign piso_data_r[57] = piso_data_r_57_sv2v_reg;
  assign piso_data_r[56] = piso_data_r_56_sv2v_reg;
  assign piso_data_r[55] = piso_data_r_55_sv2v_reg;
  assign piso_data_r[54] = piso_data_r_54_sv2v_reg;
  assign piso_data_r[53] = piso_data_r_53_sv2v_reg;
  assign piso_data_r[52] = piso_data_r_52_sv2v_reg;
  assign piso_data_r[51] = piso_data_r_51_sv2v_reg;
  assign piso_data_r[50] = piso_data_r_50_sv2v_reg;
  assign piso_data_r[49] = piso_data_r_49_sv2v_reg;
  assign piso_data_r[48] = piso_data_r_48_sv2v_reg;
  assign piso_data_r[47] = piso_data_r_47_sv2v_reg;
  assign piso_data_r[46] = piso_data_r_46_sv2v_reg;
  assign piso_data_r[45] = piso_data_r_45_sv2v_reg;
  assign piso_data_r[44] = piso_data_r_44_sv2v_reg;
  assign piso_data_r[43] = piso_data_r_43_sv2v_reg;
  assign piso_data_r[42] = piso_data_r_42_sv2v_reg;
  assign piso_data_r[41] = piso_data_r_41_sv2v_reg;
  assign piso_data_r[40] = piso_data_r_40_sv2v_reg;
  assign piso_data_r[39] = piso_data_r_39_sv2v_reg;
  assign piso_data_r[38] = piso_data_r_38_sv2v_reg;
  assign piso_data_r[37] = piso_data_r_37_sv2v_reg;
  assign piso_data_r[36] = piso_data_r_36_sv2v_reg;
  assign piso_data_r[35] = piso_data_r_35_sv2v_reg;
  assign piso_data_r[34] = piso_data_r_34_sv2v_reg;
  assign piso_data_r[33] = piso_data_r_33_sv2v_reg;
  assign piso_data_r[32] = piso_data_r_32_sv2v_reg;
  assign piso_data_r[31] = piso_data_r_31_sv2v_reg;
  assign piso_data_r[30] = piso_data_r_30_sv2v_reg;
  assign piso_data_r[29] = piso_data_r_29_sv2v_reg;
  assign piso_data_r[28] = piso_data_r_28_sv2v_reg;
  assign piso_data_r[27] = piso_data_r_27_sv2v_reg;
  assign piso_data_r[26] = piso_data_r_26_sv2v_reg;
  assign piso_data_r[25] = piso_data_r_25_sv2v_reg;
  assign piso_data_r[24] = piso_data_r_24_sv2v_reg;
  assign piso_data_r[23] = piso_data_r_23_sv2v_reg;
  assign piso_data_r[22] = piso_data_r_22_sv2v_reg;
  assign piso_data_r[21] = piso_data_r_21_sv2v_reg;
  assign piso_data_r[20] = piso_data_r_20_sv2v_reg;
  assign piso_data_r[19] = piso_data_r_19_sv2v_reg;
  assign piso_data_r[18] = piso_data_r_18_sv2v_reg;
  assign piso_data_r[17] = piso_data_r_17_sv2v_reg;
  assign piso_data_r[16] = piso_data_r_16_sv2v_reg;
  assign piso_data_r[15] = piso_data_r_15_sv2v_reg;
  assign piso_data_r[14] = piso_data_r_14_sv2v_reg;
  assign piso_data_r[13] = piso_data_r_13_sv2v_reg;
  assign piso_data_r[12] = piso_data_r_12_sv2v_reg;
  assign piso_data_r[11] = piso_data_r_11_sv2v_reg;
  assign piso_data_r[10] = piso_data_r_10_sv2v_reg;
  assign piso_data_r[9] = piso_data_r_9_sv2v_reg;
  assign piso_data_r[8] = piso_data_r_8_sv2v_reg;
  assign piso_data_r[7] = piso_data_r_7_sv2v_reg;
  assign piso_data_r[6] = piso_data_r_6_sv2v_reg;
  assign piso_data_r[5] = piso_data_r_5_sv2v_reg;
  assign piso_data_r[4] = piso_data_r_4_sv2v_reg;
  assign piso_data_r[3] = piso_data_r_3_sv2v_reg;
  assign piso_data_r[2] = piso_data_r_2_sv2v_reg;
  assign piso_data_r[1] = piso_data_r_1_sv2v_reg;
  assign piso_data_r[0] = piso_data_r_0_sv2v_reg;
  assign piso_shift_ctr_r[2] = piso_shift_ctr_r_2_sv2v_reg;
  assign piso_shift_ctr_r[1] = piso_shift_ctr_r_1_sv2v_reg;
  assign piso_shift_ctr_r[0] = piso_shift_ctr_r_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(reset_i) begin
      valid_o_sv2v_reg <= 1'b0;
    end else if(N3) begin
      valid_o_sv2v_reg <= piso_state_n[0];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_511_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_511_sv2v_reg <= data_i[511];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_510_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_510_sv2v_reg <= data_i[510];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_509_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_509_sv2v_reg <= data_i[509];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_508_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_508_sv2v_reg <= data_i[508];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_507_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_507_sv2v_reg <= data_i[507];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_506_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_506_sv2v_reg <= data_i[506];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_505_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_505_sv2v_reg <= data_i[505];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_504_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_504_sv2v_reg <= data_i[504];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_503_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_503_sv2v_reg <= data_i[503];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_502_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_502_sv2v_reg <= data_i[502];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_501_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_501_sv2v_reg <= data_i[501];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_500_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_500_sv2v_reg <= data_i[500];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_499_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_499_sv2v_reg <= data_i[499];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_498_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_498_sv2v_reg <= data_i[498];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_497_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_497_sv2v_reg <= data_i[497];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_496_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_496_sv2v_reg <= data_i[496];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_495_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_495_sv2v_reg <= data_i[495];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_494_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_494_sv2v_reg <= data_i[494];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_493_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_493_sv2v_reg <= data_i[493];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_492_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_492_sv2v_reg <= data_i[492];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_491_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_491_sv2v_reg <= data_i[491];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_490_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_490_sv2v_reg <= data_i[490];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_489_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_489_sv2v_reg <= data_i[489];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_488_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_488_sv2v_reg <= data_i[488];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_487_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_487_sv2v_reg <= data_i[487];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_486_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_486_sv2v_reg <= data_i[486];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_485_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_485_sv2v_reg <= data_i[485];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_484_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_484_sv2v_reg <= data_i[484];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_483_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_483_sv2v_reg <= data_i[483];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_482_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_482_sv2v_reg <= data_i[482];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_481_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_481_sv2v_reg <= data_i[481];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_480_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_480_sv2v_reg <= data_i[480];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_479_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_479_sv2v_reg <= data_i[479];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_478_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_478_sv2v_reg <= data_i[478];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_477_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_477_sv2v_reg <= data_i[477];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_476_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_476_sv2v_reg <= data_i[476];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_475_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_475_sv2v_reg <= data_i[475];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_474_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_474_sv2v_reg <= data_i[474];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_473_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_473_sv2v_reg <= data_i[473];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_472_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_472_sv2v_reg <= data_i[472];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_471_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_471_sv2v_reg <= data_i[471];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_470_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_470_sv2v_reg <= data_i[470];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_469_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_469_sv2v_reg <= data_i[469];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_468_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_468_sv2v_reg <= data_i[468];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_467_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_467_sv2v_reg <= data_i[467];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_466_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_466_sv2v_reg <= data_i[466];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_465_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_465_sv2v_reg <= data_i[465];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_464_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_464_sv2v_reg <= data_i[464];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_463_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_463_sv2v_reg <= data_i[463];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_462_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_462_sv2v_reg <= data_i[462];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_461_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_461_sv2v_reg <= data_i[461];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_460_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_460_sv2v_reg <= data_i[460];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_459_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_459_sv2v_reg <= data_i[459];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_458_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_458_sv2v_reg <= data_i[458];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_457_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_457_sv2v_reg <= data_i[457];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_456_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_456_sv2v_reg <= data_i[456];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_455_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_455_sv2v_reg <= data_i[455];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_454_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_454_sv2v_reg <= data_i[454];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_453_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_453_sv2v_reg <= data_i[453];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_452_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_452_sv2v_reg <= data_i[452];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_451_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_451_sv2v_reg <= data_i[451];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_450_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_450_sv2v_reg <= data_i[450];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_449_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_449_sv2v_reg <= data_i[449];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_448_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_448_sv2v_reg <= data_i[448];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_447_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_447_sv2v_reg <= data_i[447];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_446_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_446_sv2v_reg <= data_i[446];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_445_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_445_sv2v_reg <= data_i[445];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_444_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_444_sv2v_reg <= data_i[444];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_443_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_443_sv2v_reg <= data_i[443];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_442_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_442_sv2v_reg <= data_i[442];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_441_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_441_sv2v_reg <= data_i[441];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_440_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_440_sv2v_reg <= data_i[440];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_439_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_439_sv2v_reg <= data_i[439];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_438_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_438_sv2v_reg <= data_i[438];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_437_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_437_sv2v_reg <= data_i[437];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_436_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_436_sv2v_reg <= data_i[436];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_435_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_435_sv2v_reg <= data_i[435];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_434_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_434_sv2v_reg <= data_i[434];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_433_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_433_sv2v_reg <= data_i[433];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_432_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_432_sv2v_reg <= data_i[432];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_431_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_431_sv2v_reg <= data_i[431];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_430_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_430_sv2v_reg <= data_i[430];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_429_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_429_sv2v_reg <= data_i[429];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_428_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_428_sv2v_reg <= data_i[428];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_427_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_427_sv2v_reg <= data_i[427];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_426_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_426_sv2v_reg <= data_i[426];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_425_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_425_sv2v_reg <= data_i[425];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_424_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_424_sv2v_reg <= data_i[424];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_423_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_423_sv2v_reg <= data_i[423];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_422_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_422_sv2v_reg <= data_i[422];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_421_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_421_sv2v_reg <= data_i[421];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_420_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_420_sv2v_reg <= data_i[420];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_419_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_419_sv2v_reg <= data_i[419];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_418_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_418_sv2v_reg <= data_i[418];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_417_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_417_sv2v_reg <= data_i[417];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_416_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_416_sv2v_reg <= data_i[416];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_415_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_415_sv2v_reg <= data_i[415];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_414_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_414_sv2v_reg <= data_i[414];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_413_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_413_sv2v_reg <= data_i[413];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_412_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_412_sv2v_reg <= data_i[412];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_411_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_411_sv2v_reg <= data_i[411];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_410_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_410_sv2v_reg <= data_i[410];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_409_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_409_sv2v_reg <= data_i[409];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_408_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_408_sv2v_reg <= data_i[408];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_407_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_407_sv2v_reg <= data_i[407];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_406_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_406_sv2v_reg <= data_i[406];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_405_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_405_sv2v_reg <= data_i[405];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_404_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_404_sv2v_reg <= data_i[404];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_403_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_403_sv2v_reg <= data_i[403];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_402_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_402_sv2v_reg <= data_i[402];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_401_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_401_sv2v_reg <= data_i[401];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_400_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_400_sv2v_reg <= data_i[400];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_399_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_399_sv2v_reg <= data_i[399];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_398_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_398_sv2v_reg <= data_i[398];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_397_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_397_sv2v_reg <= data_i[397];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_396_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_396_sv2v_reg <= data_i[396];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_395_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_395_sv2v_reg <= data_i[395];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_394_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_394_sv2v_reg <= data_i[394];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_393_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_393_sv2v_reg <= data_i[393];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_392_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_392_sv2v_reg <= data_i[392];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_391_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_391_sv2v_reg <= data_i[391];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_390_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_390_sv2v_reg <= data_i[390];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_389_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_389_sv2v_reg <= data_i[389];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_388_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_388_sv2v_reg <= data_i[388];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_387_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_387_sv2v_reg <= data_i[387];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_386_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_386_sv2v_reg <= data_i[386];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_385_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_385_sv2v_reg <= data_i[385];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_384_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_384_sv2v_reg <= data_i[384];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_383_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_383_sv2v_reg <= data_i[383];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_382_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_382_sv2v_reg <= data_i[382];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_381_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_381_sv2v_reg <= data_i[381];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_380_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_380_sv2v_reg <= data_i[380];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_379_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_379_sv2v_reg <= data_i[379];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_378_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_378_sv2v_reg <= data_i[378];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_377_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_377_sv2v_reg <= data_i[377];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_376_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_376_sv2v_reg <= data_i[376];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_375_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_375_sv2v_reg <= data_i[375];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_374_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_374_sv2v_reg <= data_i[374];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_373_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_373_sv2v_reg <= data_i[373];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_372_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_372_sv2v_reg <= data_i[372];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_371_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_371_sv2v_reg <= data_i[371];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_370_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_370_sv2v_reg <= data_i[370];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_369_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_369_sv2v_reg <= data_i[369];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_368_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_368_sv2v_reg <= data_i[368];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_367_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_367_sv2v_reg <= data_i[367];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_366_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_366_sv2v_reg <= data_i[366];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_365_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_365_sv2v_reg <= data_i[365];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_364_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_364_sv2v_reg <= data_i[364];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_363_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_363_sv2v_reg <= data_i[363];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_362_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_362_sv2v_reg <= data_i[362];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_361_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_361_sv2v_reg <= data_i[361];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_360_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_360_sv2v_reg <= data_i[360];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_359_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_359_sv2v_reg <= data_i[359];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_358_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_358_sv2v_reg <= data_i[358];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_357_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_357_sv2v_reg <= data_i[357];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_356_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_356_sv2v_reg <= data_i[356];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_355_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_355_sv2v_reg <= data_i[355];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_354_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_354_sv2v_reg <= data_i[354];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_353_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_353_sv2v_reg <= data_i[353];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_352_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_352_sv2v_reg <= data_i[352];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_351_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_351_sv2v_reg <= data_i[351];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_350_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_350_sv2v_reg <= data_i[350];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_349_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_349_sv2v_reg <= data_i[349];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_348_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_348_sv2v_reg <= data_i[348];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_347_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_347_sv2v_reg <= data_i[347];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_346_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_346_sv2v_reg <= data_i[346];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_345_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_345_sv2v_reg <= data_i[345];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_344_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_344_sv2v_reg <= data_i[344];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_343_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_343_sv2v_reg <= data_i[343];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_342_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_342_sv2v_reg <= data_i[342];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_341_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_341_sv2v_reg <= data_i[341];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_340_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_340_sv2v_reg <= data_i[340];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_339_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_339_sv2v_reg <= data_i[339];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_338_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_338_sv2v_reg <= data_i[338];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_337_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_337_sv2v_reg <= data_i[337];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_336_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_336_sv2v_reg <= data_i[336];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_335_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_335_sv2v_reg <= data_i[335];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_334_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_334_sv2v_reg <= data_i[334];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_333_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_333_sv2v_reg <= data_i[333];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_332_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_332_sv2v_reg <= data_i[332];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_331_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_331_sv2v_reg <= data_i[331];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_330_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_330_sv2v_reg <= data_i[330];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_329_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_329_sv2v_reg <= data_i[329];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_328_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_328_sv2v_reg <= data_i[328];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_327_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_327_sv2v_reg <= data_i[327];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_326_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_326_sv2v_reg <= data_i[326];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_325_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_325_sv2v_reg <= data_i[325];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_324_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_324_sv2v_reg <= data_i[324];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_323_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_323_sv2v_reg <= data_i[323];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_322_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_322_sv2v_reg <= data_i[322];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_321_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_321_sv2v_reg <= data_i[321];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_320_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_320_sv2v_reg <= data_i[320];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_319_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_319_sv2v_reg <= data_i[319];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_318_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_318_sv2v_reg <= data_i[318];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_317_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_317_sv2v_reg <= data_i[317];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_316_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_316_sv2v_reg <= data_i[316];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_315_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_315_sv2v_reg <= data_i[315];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_314_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_314_sv2v_reg <= data_i[314];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_313_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_313_sv2v_reg <= data_i[313];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_312_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_312_sv2v_reg <= data_i[312];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_311_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_311_sv2v_reg <= data_i[311];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_310_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_310_sv2v_reg <= data_i[310];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_309_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_309_sv2v_reg <= data_i[309];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_308_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_308_sv2v_reg <= data_i[308];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_307_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_307_sv2v_reg <= data_i[307];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_306_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_306_sv2v_reg <= data_i[306];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_305_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_305_sv2v_reg <= data_i[305];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_304_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_304_sv2v_reg <= data_i[304];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_303_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_303_sv2v_reg <= data_i[303];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_302_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_302_sv2v_reg <= data_i[302];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_301_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_301_sv2v_reg <= data_i[301];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_300_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_300_sv2v_reg <= data_i[300];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_299_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_299_sv2v_reg <= data_i[299];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_298_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_298_sv2v_reg <= data_i[298];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_297_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_297_sv2v_reg <= data_i[297];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_296_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_296_sv2v_reg <= data_i[296];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_295_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_295_sv2v_reg <= data_i[295];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_294_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_294_sv2v_reg <= data_i[294];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_293_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_293_sv2v_reg <= data_i[293];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_292_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_292_sv2v_reg <= data_i[292];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_291_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_291_sv2v_reg <= data_i[291];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_290_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_290_sv2v_reg <= data_i[290];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_289_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_289_sv2v_reg <= data_i[289];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_288_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_288_sv2v_reg <= data_i[288];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_287_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_287_sv2v_reg <= data_i[287];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_286_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_286_sv2v_reg <= data_i[286];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_285_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_285_sv2v_reg <= data_i[285];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_284_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_284_sv2v_reg <= data_i[284];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_283_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_283_sv2v_reg <= data_i[283];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_282_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_282_sv2v_reg <= data_i[282];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_281_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_281_sv2v_reg <= data_i[281];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_280_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_280_sv2v_reg <= data_i[280];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_279_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_279_sv2v_reg <= data_i[279];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_278_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_278_sv2v_reg <= data_i[278];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_277_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_277_sv2v_reg <= data_i[277];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_276_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_276_sv2v_reg <= data_i[276];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_275_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_275_sv2v_reg <= data_i[275];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_274_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_274_sv2v_reg <= data_i[274];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_273_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_273_sv2v_reg <= data_i[273];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_272_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_272_sv2v_reg <= data_i[272];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_271_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_271_sv2v_reg <= data_i[271];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_270_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_270_sv2v_reg <= data_i[270];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_269_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_269_sv2v_reg <= data_i[269];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_268_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_268_sv2v_reg <= data_i[268];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_267_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_267_sv2v_reg <= data_i[267];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_266_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_266_sv2v_reg <= data_i[266];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_265_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_265_sv2v_reg <= data_i[265];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_264_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_264_sv2v_reg <= data_i[264];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_263_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_263_sv2v_reg <= data_i[263];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_262_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_262_sv2v_reg <= data_i[262];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_261_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_261_sv2v_reg <= data_i[261];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_260_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_260_sv2v_reg <= data_i[260];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_259_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_259_sv2v_reg <= data_i[259];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_258_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_258_sv2v_reg <= data_i[258];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_257_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_257_sv2v_reg <= data_i[257];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_256_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_256_sv2v_reg <= data_i[256];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_255_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_255_sv2v_reg <= data_i[255];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_254_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_254_sv2v_reg <= data_i[254];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_253_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_253_sv2v_reg <= data_i[253];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_252_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_252_sv2v_reg <= data_i[252];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_251_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_251_sv2v_reg <= data_i[251];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_250_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_250_sv2v_reg <= data_i[250];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_249_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_249_sv2v_reg <= data_i[249];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_248_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_248_sv2v_reg <= data_i[248];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_247_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_247_sv2v_reg <= data_i[247];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_246_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_246_sv2v_reg <= data_i[246];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_245_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_245_sv2v_reg <= data_i[245];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_244_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_244_sv2v_reg <= data_i[244];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_243_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_243_sv2v_reg <= data_i[243];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_242_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_242_sv2v_reg <= data_i[242];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_241_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_241_sv2v_reg <= data_i[241];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_240_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_240_sv2v_reg <= data_i[240];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_239_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_239_sv2v_reg <= data_i[239];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_238_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_238_sv2v_reg <= data_i[238];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_237_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_237_sv2v_reg <= data_i[237];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_236_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_236_sv2v_reg <= data_i[236];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_235_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_235_sv2v_reg <= data_i[235];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_234_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_234_sv2v_reg <= data_i[234];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_233_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_233_sv2v_reg <= data_i[233];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_232_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_232_sv2v_reg <= data_i[232];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_231_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_231_sv2v_reg <= data_i[231];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_230_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_230_sv2v_reg <= data_i[230];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_229_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_229_sv2v_reg <= data_i[229];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_228_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_228_sv2v_reg <= data_i[228];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_227_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_227_sv2v_reg <= data_i[227];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_226_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_226_sv2v_reg <= data_i[226];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_225_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_225_sv2v_reg <= data_i[225];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_224_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_224_sv2v_reg <= data_i[224];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_223_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_223_sv2v_reg <= data_i[223];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_222_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_222_sv2v_reg <= data_i[222];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_221_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_221_sv2v_reg <= data_i[221];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_220_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_220_sv2v_reg <= data_i[220];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_219_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_219_sv2v_reg <= data_i[219];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_218_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_218_sv2v_reg <= data_i[218];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_217_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_217_sv2v_reg <= data_i[217];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_216_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_216_sv2v_reg <= data_i[216];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_215_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_215_sv2v_reg <= data_i[215];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_214_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_214_sv2v_reg <= data_i[214];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_213_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_213_sv2v_reg <= data_i[213];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_212_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_212_sv2v_reg <= data_i[212];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_211_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_211_sv2v_reg <= data_i[211];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_210_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_210_sv2v_reg <= data_i[210];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_209_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_209_sv2v_reg <= data_i[209];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_208_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_208_sv2v_reg <= data_i[208];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_207_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_207_sv2v_reg <= data_i[207];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_206_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_206_sv2v_reg <= data_i[206];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_205_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_205_sv2v_reg <= data_i[205];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_204_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_204_sv2v_reg <= data_i[204];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_203_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_203_sv2v_reg <= data_i[203];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_202_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_202_sv2v_reg <= data_i[202];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_201_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_201_sv2v_reg <= data_i[201];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_200_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_200_sv2v_reg <= data_i[200];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_199_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_199_sv2v_reg <= data_i[199];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_198_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_198_sv2v_reg <= data_i[198];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_197_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_197_sv2v_reg <= data_i[197];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_196_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_196_sv2v_reg <= data_i[196];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_195_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_195_sv2v_reg <= data_i[195];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_194_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_194_sv2v_reg <= data_i[194];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_193_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_193_sv2v_reg <= data_i[193];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_192_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_192_sv2v_reg <= data_i[192];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_191_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_191_sv2v_reg <= data_i[191];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_190_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_190_sv2v_reg <= data_i[190];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_189_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_189_sv2v_reg <= data_i[189];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_188_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_188_sv2v_reg <= data_i[188];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_187_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_187_sv2v_reg <= data_i[187];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_186_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_186_sv2v_reg <= data_i[186];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_185_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_185_sv2v_reg <= data_i[185];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_184_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_184_sv2v_reg <= data_i[184];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_183_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_183_sv2v_reg <= data_i[183];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_182_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_182_sv2v_reg <= data_i[182];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_181_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_181_sv2v_reg <= data_i[181];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_180_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_180_sv2v_reg <= data_i[180];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_179_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_179_sv2v_reg <= data_i[179];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_178_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_178_sv2v_reg <= data_i[178];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_177_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_177_sv2v_reg <= data_i[177];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_176_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_176_sv2v_reg <= data_i[176];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_175_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_175_sv2v_reg <= data_i[175];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_174_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_174_sv2v_reg <= data_i[174];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_173_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_173_sv2v_reg <= data_i[173];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_172_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_172_sv2v_reg <= data_i[172];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_171_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_171_sv2v_reg <= data_i[171];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_170_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_170_sv2v_reg <= data_i[170];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_169_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_169_sv2v_reg <= data_i[169];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_168_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_168_sv2v_reg <= data_i[168];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_167_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_167_sv2v_reg <= data_i[167];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_166_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_166_sv2v_reg <= data_i[166];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_165_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_165_sv2v_reg <= data_i[165];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_164_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_164_sv2v_reg <= data_i[164];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_163_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_163_sv2v_reg <= data_i[163];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_162_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_162_sv2v_reg <= data_i[162];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_161_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_161_sv2v_reg <= data_i[161];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_160_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_160_sv2v_reg <= data_i[160];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_159_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_159_sv2v_reg <= data_i[159];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_158_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_158_sv2v_reg <= data_i[158];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_157_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_157_sv2v_reg <= data_i[157];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_156_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_156_sv2v_reg <= data_i[156];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_155_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_155_sv2v_reg <= data_i[155];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_154_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_154_sv2v_reg <= data_i[154];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_153_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_153_sv2v_reg <= data_i[153];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_152_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_152_sv2v_reg <= data_i[152];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_151_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_151_sv2v_reg <= data_i[151];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_150_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_150_sv2v_reg <= data_i[150];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_149_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_149_sv2v_reg <= data_i[149];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_148_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_148_sv2v_reg <= data_i[148];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_147_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_147_sv2v_reg <= data_i[147];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_146_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_146_sv2v_reg <= data_i[146];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_145_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_145_sv2v_reg <= data_i[145];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_144_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_144_sv2v_reg <= data_i[144];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_143_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_143_sv2v_reg <= data_i[143];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_142_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_142_sv2v_reg <= data_i[142];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_141_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_141_sv2v_reg <= data_i[141];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_140_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_140_sv2v_reg <= data_i[140];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_139_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_139_sv2v_reg <= data_i[139];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_138_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_138_sv2v_reg <= data_i[138];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_137_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_137_sv2v_reg <= data_i[137];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_136_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_136_sv2v_reg <= data_i[136];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_135_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_135_sv2v_reg <= data_i[135];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_134_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_134_sv2v_reg <= data_i[134];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_133_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_133_sv2v_reg <= data_i[133];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_132_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_132_sv2v_reg <= data_i[132];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_131_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_131_sv2v_reg <= data_i[131];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_130_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_130_sv2v_reg <= data_i[130];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_129_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_129_sv2v_reg <= data_i[129];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_128_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_128_sv2v_reg <= data_i[128];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_127_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_127_sv2v_reg <= data_i[127];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_126_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_126_sv2v_reg <= data_i[126];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_125_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_125_sv2v_reg <= data_i[125];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_124_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_124_sv2v_reg <= data_i[124];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_123_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_123_sv2v_reg <= data_i[123];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_122_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_122_sv2v_reg <= data_i[122];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_121_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_121_sv2v_reg <= data_i[121];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_120_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_120_sv2v_reg <= data_i[120];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_119_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_119_sv2v_reg <= data_i[119];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_118_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_118_sv2v_reg <= data_i[118];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_117_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_117_sv2v_reg <= data_i[117];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_116_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_116_sv2v_reg <= data_i[116];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_115_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_115_sv2v_reg <= data_i[115];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_114_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_114_sv2v_reg <= data_i[114];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_113_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_113_sv2v_reg <= data_i[113];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_112_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_112_sv2v_reg <= data_i[112];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_111_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_111_sv2v_reg <= data_i[111];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_110_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_110_sv2v_reg <= data_i[110];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_109_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_109_sv2v_reg <= data_i[109];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_108_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_108_sv2v_reg <= data_i[108];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_107_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_107_sv2v_reg <= data_i[107];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_106_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_106_sv2v_reg <= data_i[106];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_105_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_105_sv2v_reg <= data_i[105];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_104_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_104_sv2v_reg <= data_i[104];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_103_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_103_sv2v_reg <= data_i[103];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_102_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_102_sv2v_reg <= data_i[102];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_101_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_101_sv2v_reg <= data_i[101];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_100_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_100_sv2v_reg <= data_i[100];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_99_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_99_sv2v_reg <= data_i[99];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_98_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_98_sv2v_reg <= data_i[98];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_97_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_97_sv2v_reg <= data_i[97];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_96_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_96_sv2v_reg <= data_i[96];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_95_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_95_sv2v_reg <= data_i[95];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_94_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_94_sv2v_reg <= data_i[94];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_93_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_93_sv2v_reg <= data_i[93];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_92_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_92_sv2v_reg <= data_i[92];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_91_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_91_sv2v_reg <= data_i[91];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_90_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_90_sv2v_reg <= data_i[90];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_89_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_89_sv2v_reg <= data_i[89];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_88_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_88_sv2v_reg <= data_i[88];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_87_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_87_sv2v_reg <= data_i[87];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_86_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_86_sv2v_reg <= data_i[86];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_85_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_85_sv2v_reg <= data_i[85];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_84_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_84_sv2v_reg <= data_i[84];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_83_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_83_sv2v_reg <= data_i[83];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_82_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_82_sv2v_reg <= data_i[82];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_81_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_81_sv2v_reg <= data_i[81];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_80_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_80_sv2v_reg <= data_i[80];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_79_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_79_sv2v_reg <= data_i[79];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_78_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_78_sv2v_reg <= data_i[78];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_77_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_77_sv2v_reg <= data_i[77];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_76_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_76_sv2v_reg <= data_i[76];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_75_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_75_sv2v_reg <= data_i[75];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_74_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_74_sv2v_reg <= data_i[74];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_73_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_73_sv2v_reg <= data_i[73];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_72_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_72_sv2v_reg <= data_i[72];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_71_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_71_sv2v_reg <= data_i[71];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_70_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_70_sv2v_reg <= data_i[70];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_69_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_69_sv2v_reg <= data_i[69];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_68_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_68_sv2v_reg <= data_i[68];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_67_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_67_sv2v_reg <= data_i[67];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_66_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_66_sv2v_reg <= data_i[66];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_65_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_65_sv2v_reg <= data_i[65];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_64_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_64_sv2v_reg <= data_i[64];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_63_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_63_sv2v_reg <= data_i[63];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_62_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_62_sv2v_reg <= data_i[62];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_61_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_61_sv2v_reg <= data_i[61];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_60_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_60_sv2v_reg <= data_i[60];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_59_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_59_sv2v_reg <= data_i[59];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_58_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_58_sv2v_reg <= data_i[58];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_57_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_57_sv2v_reg <= data_i[57];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_56_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_56_sv2v_reg <= data_i[56];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_55_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_55_sv2v_reg <= data_i[55];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_54_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_54_sv2v_reg <= data_i[54];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_53_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_53_sv2v_reg <= data_i[53];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_52_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_52_sv2v_reg <= data_i[52];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_51_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_51_sv2v_reg <= data_i[51];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_50_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_50_sv2v_reg <= data_i[50];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_49_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_49_sv2v_reg <= data_i[49];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_48_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_48_sv2v_reg <= data_i[48];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_47_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_47_sv2v_reg <= data_i[47];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_46_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_46_sv2v_reg <= data_i[46];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_45_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_45_sv2v_reg <= data_i[45];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_44_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_44_sv2v_reg <= data_i[44];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_43_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_43_sv2v_reg <= data_i[43];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_42_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_42_sv2v_reg <= data_i[42];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_41_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_41_sv2v_reg <= data_i[41];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_40_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_40_sv2v_reg <= data_i[40];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_39_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_39_sv2v_reg <= data_i[39];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_38_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_38_sv2v_reg <= data_i[38];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_37_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_37_sv2v_reg <= data_i[37];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_36_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_36_sv2v_reg <= data_i[36];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_35_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_35_sv2v_reg <= data_i[35];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_34_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_34_sv2v_reg <= data_i[34];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_33_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_33_sv2v_reg <= data_i[33];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_32_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_32_sv2v_reg <= data_i[32];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_31_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_31_sv2v_reg <= data_i[31];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_30_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_30_sv2v_reg <= data_i[30];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_29_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_29_sv2v_reg <= data_i[29];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_28_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_28_sv2v_reg <= data_i[28];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_27_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_27_sv2v_reg <= data_i[27];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_26_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_26_sv2v_reg <= data_i[26];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_25_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_25_sv2v_reg <= data_i[25];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_24_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_24_sv2v_reg <= data_i[24];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_23_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_23_sv2v_reg <= data_i[23];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_22_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_22_sv2v_reg <= data_i[22];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_21_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_21_sv2v_reg <= data_i[21];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_20_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_20_sv2v_reg <= data_i[20];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_19_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_19_sv2v_reg <= data_i[19];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_18_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_18_sv2v_reg <= data_i[18];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_17_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_17_sv2v_reg <= data_i[17];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_16_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_16_sv2v_reg <= data_i[16];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_15_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_15_sv2v_reg <= data_i[15];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_14_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_14_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_13_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_13_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_12_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_12_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_11_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_11_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_10_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_10_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_9_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_9_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_8_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_8_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_7_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_7_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_6_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_6_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_5_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_5_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_4_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_4_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_3_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_3_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_2_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_2_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_1_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_1_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_data_r_0_sv2v_reg <= 1'b0;
    end else if(N6) begin
      piso_data_r_0_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_shift_ctr_r_2_sv2v_reg <= 1'b0;
    end else if(N33) begin
      piso_shift_ctr_r_2_sv2v_reg <= N11;
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_shift_ctr_r_1_sv2v_reg <= 1'b0;
    end else if(N33) begin
      piso_shift_ctr_r_1_sv2v_reg <= N10;
    end 
  end


  always @(posedge clk_i) begin
    if(reset_i) begin
      piso_shift_ctr_r_0_sv2v_reg <= 1'b0;
    end else if(N33) begin
      piso_shift_ctr_r_0_sv2v_reg <= N9;
    end 
  end

  assign data_o[63] = (N24)? piso_data_r[63] : 
                      (N26)? piso_data_r[127] : 
                      (N28)? piso_data_r[191] : 
                      (N30)? piso_data_r[255] : 
                      (N25)? piso_data_r[319] : 
                      (N27)? piso_data_r[383] : 
                      (N29)? piso_data_r[447] : 
                      (N31)? piso_data_r[511] : 1'b0;
  assign data_o[62] = (N24)? piso_data_r[62] : 
                      (N26)? piso_data_r[126] : 
                      (N28)? piso_data_r[190] : 
                      (N30)? piso_data_r[254] : 
                      (N25)? piso_data_r[318] : 
                      (N27)? piso_data_r[382] : 
                      (N29)? piso_data_r[446] : 
                      (N31)? piso_data_r[510] : 1'b0;
  assign data_o[61] = (N24)? piso_data_r[61] : 
                      (N26)? piso_data_r[125] : 
                      (N28)? piso_data_r[189] : 
                      (N30)? piso_data_r[253] : 
                      (N25)? piso_data_r[317] : 
                      (N27)? piso_data_r[381] : 
                      (N29)? piso_data_r[445] : 
                      (N31)? piso_data_r[509] : 1'b0;
  assign data_o[60] = (N24)? piso_data_r[60] : 
                      (N26)? piso_data_r[124] : 
                      (N28)? piso_data_r[188] : 
                      (N30)? piso_data_r[252] : 
                      (N25)? piso_data_r[316] : 
                      (N27)? piso_data_r[380] : 
                      (N29)? piso_data_r[444] : 
                      (N31)? piso_data_r[508] : 1'b0;
  assign data_o[59] = (N24)? piso_data_r[59] : 
                      (N26)? piso_data_r[123] : 
                      (N28)? piso_data_r[187] : 
                      (N30)? piso_data_r[251] : 
                      (N25)? piso_data_r[315] : 
                      (N27)? piso_data_r[379] : 
                      (N29)? piso_data_r[443] : 
                      (N31)? piso_data_r[507] : 1'b0;
  assign data_o[58] = (N24)? piso_data_r[58] : 
                      (N26)? piso_data_r[122] : 
                      (N28)? piso_data_r[186] : 
                      (N30)? piso_data_r[250] : 
                      (N25)? piso_data_r[314] : 
                      (N27)? piso_data_r[378] : 
                      (N29)? piso_data_r[442] : 
                      (N31)? piso_data_r[506] : 1'b0;
  assign data_o[57] = (N24)? piso_data_r[57] : 
                      (N26)? piso_data_r[121] : 
                      (N28)? piso_data_r[185] : 
                      (N30)? piso_data_r[249] : 
                      (N25)? piso_data_r[313] : 
                      (N27)? piso_data_r[377] : 
                      (N29)? piso_data_r[441] : 
                      (N31)? piso_data_r[505] : 1'b0;
  assign data_o[56] = (N24)? piso_data_r[56] : 
                      (N26)? piso_data_r[120] : 
                      (N28)? piso_data_r[184] : 
                      (N30)? piso_data_r[248] : 
                      (N25)? piso_data_r[312] : 
                      (N27)? piso_data_r[376] : 
                      (N29)? piso_data_r[440] : 
                      (N31)? piso_data_r[504] : 1'b0;
  assign data_o[55] = (N24)? piso_data_r[55] : 
                      (N26)? piso_data_r[119] : 
                      (N28)? piso_data_r[183] : 
                      (N30)? piso_data_r[247] : 
                      (N25)? piso_data_r[311] : 
                      (N27)? piso_data_r[375] : 
                      (N29)? piso_data_r[439] : 
                      (N31)? piso_data_r[503] : 1'b0;
  assign data_o[54] = (N24)? piso_data_r[54] : 
                      (N26)? piso_data_r[118] : 
                      (N28)? piso_data_r[182] : 
                      (N30)? piso_data_r[246] : 
                      (N25)? piso_data_r[310] : 
                      (N27)? piso_data_r[374] : 
                      (N29)? piso_data_r[438] : 
                      (N31)? piso_data_r[502] : 1'b0;
  assign data_o[53] = (N24)? piso_data_r[53] : 
                      (N26)? piso_data_r[117] : 
                      (N28)? piso_data_r[181] : 
                      (N30)? piso_data_r[245] : 
                      (N25)? piso_data_r[309] : 
                      (N27)? piso_data_r[373] : 
                      (N29)? piso_data_r[437] : 
                      (N31)? piso_data_r[501] : 1'b0;
  assign data_o[52] = (N24)? piso_data_r[52] : 
                      (N26)? piso_data_r[116] : 
                      (N28)? piso_data_r[180] : 
                      (N30)? piso_data_r[244] : 
                      (N25)? piso_data_r[308] : 
                      (N27)? piso_data_r[372] : 
                      (N29)? piso_data_r[436] : 
                      (N31)? piso_data_r[500] : 1'b0;
  assign data_o[51] = (N24)? piso_data_r[51] : 
                      (N26)? piso_data_r[115] : 
                      (N28)? piso_data_r[179] : 
                      (N30)? piso_data_r[243] : 
                      (N25)? piso_data_r[307] : 
                      (N27)? piso_data_r[371] : 
                      (N29)? piso_data_r[435] : 
                      (N31)? piso_data_r[499] : 1'b0;
  assign data_o[50] = (N24)? piso_data_r[50] : 
                      (N26)? piso_data_r[114] : 
                      (N28)? piso_data_r[178] : 
                      (N30)? piso_data_r[242] : 
                      (N25)? piso_data_r[306] : 
                      (N27)? piso_data_r[370] : 
                      (N29)? piso_data_r[434] : 
                      (N31)? piso_data_r[498] : 1'b0;
  assign data_o[49] = (N24)? piso_data_r[49] : 
                      (N26)? piso_data_r[113] : 
                      (N28)? piso_data_r[177] : 
                      (N30)? piso_data_r[241] : 
                      (N25)? piso_data_r[305] : 
                      (N27)? piso_data_r[369] : 
                      (N29)? piso_data_r[433] : 
                      (N31)? piso_data_r[497] : 1'b0;
  assign data_o[48] = (N24)? piso_data_r[48] : 
                      (N26)? piso_data_r[112] : 
                      (N28)? piso_data_r[176] : 
                      (N30)? piso_data_r[240] : 
                      (N25)? piso_data_r[304] : 
                      (N27)? piso_data_r[368] : 
                      (N29)? piso_data_r[432] : 
                      (N31)? piso_data_r[496] : 1'b0;
  assign data_o[47] = (N24)? piso_data_r[47] : 
                      (N26)? piso_data_r[111] : 
                      (N28)? piso_data_r[175] : 
                      (N30)? piso_data_r[239] : 
                      (N25)? piso_data_r[303] : 
                      (N27)? piso_data_r[367] : 
                      (N29)? piso_data_r[431] : 
                      (N31)? piso_data_r[495] : 1'b0;
  assign data_o[46] = (N24)? piso_data_r[46] : 
                      (N26)? piso_data_r[110] : 
                      (N28)? piso_data_r[174] : 
                      (N30)? piso_data_r[238] : 
                      (N25)? piso_data_r[302] : 
                      (N27)? piso_data_r[366] : 
                      (N29)? piso_data_r[430] : 
                      (N31)? piso_data_r[494] : 1'b0;
  assign data_o[45] = (N24)? piso_data_r[45] : 
                      (N26)? piso_data_r[109] : 
                      (N28)? piso_data_r[173] : 
                      (N30)? piso_data_r[237] : 
                      (N25)? piso_data_r[301] : 
                      (N27)? piso_data_r[365] : 
                      (N29)? piso_data_r[429] : 
                      (N31)? piso_data_r[493] : 1'b0;
  assign data_o[44] = (N24)? piso_data_r[44] : 
                      (N26)? piso_data_r[108] : 
                      (N28)? piso_data_r[172] : 
                      (N30)? piso_data_r[236] : 
                      (N25)? piso_data_r[300] : 
                      (N27)? piso_data_r[364] : 
                      (N29)? piso_data_r[428] : 
                      (N31)? piso_data_r[492] : 1'b0;
  assign data_o[43] = (N24)? piso_data_r[43] : 
                      (N26)? piso_data_r[107] : 
                      (N28)? piso_data_r[171] : 
                      (N30)? piso_data_r[235] : 
                      (N25)? piso_data_r[299] : 
                      (N27)? piso_data_r[363] : 
                      (N29)? piso_data_r[427] : 
                      (N31)? piso_data_r[491] : 1'b0;
  assign data_o[42] = (N24)? piso_data_r[42] : 
                      (N26)? piso_data_r[106] : 
                      (N28)? piso_data_r[170] : 
                      (N30)? piso_data_r[234] : 
                      (N25)? piso_data_r[298] : 
                      (N27)? piso_data_r[362] : 
                      (N29)? piso_data_r[426] : 
                      (N31)? piso_data_r[490] : 1'b0;
  assign data_o[41] = (N24)? piso_data_r[41] : 
                      (N26)? piso_data_r[105] : 
                      (N28)? piso_data_r[169] : 
                      (N30)? piso_data_r[233] : 
                      (N25)? piso_data_r[297] : 
                      (N27)? piso_data_r[361] : 
                      (N29)? piso_data_r[425] : 
                      (N31)? piso_data_r[489] : 1'b0;
  assign data_o[40] = (N24)? piso_data_r[40] : 
                      (N26)? piso_data_r[104] : 
                      (N28)? piso_data_r[168] : 
                      (N30)? piso_data_r[232] : 
                      (N25)? piso_data_r[296] : 
                      (N27)? piso_data_r[360] : 
                      (N29)? piso_data_r[424] : 
                      (N31)? piso_data_r[488] : 1'b0;
  assign data_o[39] = (N24)? piso_data_r[39] : 
                      (N26)? piso_data_r[103] : 
                      (N28)? piso_data_r[167] : 
                      (N30)? piso_data_r[231] : 
                      (N25)? piso_data_r[295] : 
                      (N27)? piso_data_r[359] : 
                      (N29)? piso_data_r[423] : 
                      (N31)? piso_data_r[487] : 1'b0;
  assign data_o[38] = (N24)? piso_data_r[38] : 
                      (N26)? piso_data_r[102] : 
                      (N28)? piso_data_r[166] : 
                      (N30)? piso_data_r[230] : 
                      (N25)? piso_data_r[294] : 
                      (N27)? piso_data_r[358] : 
                      (N29)? piso_data_r[422] : 
                      (N31)? piso_data_r[486] : 1'b0;
  assign data_o[37] = (N24)? piso_data_r[37] : 
                      (N26)? piso_data_r[101] : 
                      (N28)? piso_data_r[165] : 
                      (N30)? piso_data_r[229] : 
                      (N25)? piso_data_r[293] : 
                      (N27)? piso_data_r[357] : 
                      (N29)? piso_data_r[421] : 
                      (N31)? piso_data_r[485] : 1'b0;
  assign data_o[36] = (N24)? piso_data_r[36] : 
                      (N26)? piso_data_r[100] : 
                      (N28)? piso_data_r[164] : 
                      (N30)? piso_data_r[228] : 
                      (N25)? piso_data_r[292] : 
                      (N27)? piso_data_r[356] : 
                      (N29)? piso_data_r[420] : 
                      (N31)? piso_data_r[484] : 1'b0;
  assign data_o[35] = (N24)? piso_data_r[35] : 
                      (N26)? piso_data_r[99] : 
                      (N28)? piso_data_r[163] : 
                      (N30)? piso_data_r[227] : 
                      (N25)? piso_data_r[291] : 
                      (N27)? piso_data_r[355] : 
                      (N29)? piso_data_r[419] : 
                      (N31)? piso_data_r[483] : 1'b0;
  assign data_o[34] = (N24)? piso_data_r[34] : 
                      (N26)? piso_data_r[98] : 
                      (N28)? piso_data_r[162] : 
                      (N30)? piso_data_r[226] : 
                      (N25)? piso_data_r[290] : 
                      (N27)? piso_data_r[354] : 
                      (N29)? piso_data_r[418] : 
                      (N31)? piso_data_r[482] : 1'b0;
  assign data_o[33] = (N24)? piso_data_r[33] : 
                      (N26)? piso_data_r[97] : 
                      (N28)? piso_data_r[161] : 
                      (N30)? piso_data_r[225] : 
                      (N25)? piso_data_r[289] : 
                      (N27)? piso_data_r[353] : 
                      (N29)? piso_data_r[417] : 
                      (N31)? piso_data_r[481] : 1'b0;
  assign data_o[32] = (N24)? piso_data_r[32] : 
                      (N26)? piso_data_r[96] : 
                      (N28)? piso_data_r[160] : 
                      (N30)? piso_data_r[224] : 
                      (N25)? piso_data_r[288] : 
                      (N27)? piso_data_r[352] : 
                      (N29)? piso_data_r[416] : 
                      (N31)? piso_data_r[480] : 1'b0;
  assign data_o[31] = (N24)? piso_data_r[31] : 
                      (N26)? piso_data_r[95] : 
                      (N28)? piso_data_r[159] : 
                      (N30)? piso_data_r[223] : 
                      (N25)? piso_data_r[287] : 
                      (N27)? piso_data_r[351] : 
                      (N29)? piso_data_r[415] : 
                      (N31)? piso_data_r[479] : 1'b0;
  assign data_o[30] = (N24)? piso_data_r[30] : 
                      (N26)? piso_data_r[94] : 
                      (N28)? piso_data_r[158] : 
                      (N30)? piso_data_r[222] : 
                      (N25)? piso_data_r[286] : 
                      (N27)? piso_data_r[350] : 
                      (N29)? piso_data_r[414] : 
                      (N31)? piso_data_r[478] : 1'b0;
  assign data_o[29] = (N24)? piso_data_r[29] : 
                      (N26)? piso_data_r[93] : 
                      (N28)? piso_data_r[157] : 
                      (N30)? piso_data_r[221] : 
                      (N25)? piso_data_r[285] : 
                      (N27)? piso_data_r[349] : 
                      (N29)? piso_data_r[413] : 
                      (N31)? piso_data_r[477] : 1'b0;
  assign data_o[28] = (N24)? piso_data_r[28] : 
                      (N26)? piso_data_r[92] : 
                      (N28)? piso_data_r[156] : 
                      (N30)? piso_data_r[220] : 
                      (N25)? piso_data_r[284] : 
                      (N27)? piso_data_r[348] : 
                      (N29)? piso_data_r[412] : 
                      (N31)? piso_data_r[476] : 1'b0;
  assign data_o[27] = (N24)? piso_data_r[27] : 
                      (N26)? piso_data_r[91] : 
                      (N28)? piso_data_r[155] : 
                      (N30)? piso_data_r[219] : 
                      (N25)? piso_data_r[283] : 
                      (N27)? piso_data_r[347] : 
                      (N29)? piso_data_r[411] : 
                      (N31)? piso_data_r[475] : 1'b0;
  assign data_o[26] = (N24)? piso_data_r[26] : 
                      (N26)? piso_data_r[90] : 
                      (N28)? piso_data_r[154] : 
                      (N30)? piso_data_r[218] : 
                      (N25)? piso_data_r[282] : 
                      (N27)? piso_data_r[346] : 
                      (N29)? piso_data_r[410] : 
                      (N31)? piso_data_r[474] : 1'b0;
  assign data_o[25] = (N24)? piso_data_r[25] : 
                      (N26)? piso_data_r[89] : 
                      (N28)? piso_data_r[153] : 
                      (N30)? piso_data_r[217] : 
                      (N25)? piso_data_r[281] : 
                      (N27)? piso_data_r[345] : 
                      (N29)? piso_data_r[409] : 
                      (N31)? piso_data_r[473] : 1'b0;
  assign data_o[24] = (N24)? piso_data_r[24] : 
                      (N26)? piso_data_r[88] : 
                      (N28)? piso_data_r[152] : 
                      (N30)? piso_data_r[216] : 
                      (N25)? piso_data_r[280] : 
                      (N27)? piso_data_r[344] : 
                      (N29)? piso_data_r[408] : 
                      (N31)? piso_data_r[472] : 1'b0;
  assign data_o[23] = (N24)? piso_data_r[23] : 
                      (N26)? piso_data_r[87] : 
                      (N28)? piso_data_r[151] : 
                      (N30)? piso_data_r[215] : 
                      (N25)? piso_data_r[279] : 
                      (N27)? piso_data_r[343] : 
                      (N29)? piso_data_r[407] : 
                      (N31)? piso_data_r[471] : 1'b0;
  assign data_o[22] = (N24)? piso_data_r[22] : 
                      (N26)? piso_data_r[86] : 
                      (N28)? piso_data_r[150] : 
                      (N30)? piso_data_r[214] : 
                      (N25)? piso_data_r[278] : 
                      (N27)? piso_data_r[342] : 
                      (N29)? piso_data_r[406] : 
                      (N31)? piso_data_r[470] : 1'b0;
  assign data_o[21] = (N24)? piso_data_r[21] : 
                      (N26)? piso_data_r[85] : 
                      (N28)? piso_data_r[149] : 
                      (N30)? piso_data_r[213] : 
                      (N25)? piso_data_r[277] : 
                      (N27)? piso_data_r[341] : 
                      (N29)? piso_data_r[405] : 
                      (N31)? piso_data_r[469] : 1'b0;
  assign data_o[20] = (N24)? piso_data_r[20] : 
                      (N26)? piso_data_r[84] : 
                      (N28)? piso_data_r[148] : 
                      (N30)? piso_data_r[212] : 
                      (N25)? piso_data_r[276] : 
                      (N27)? piso_data_r[340] : 
                      (N29)? piso_data_r[404] : 
                      (N31)? piso_data_r[468] : 1'b0;
  assign data_o[19] = (N24)? piso_data_r[19] : 
                      (N26)? piso_data_r[83] : 
                      (N28)? piso_data_r[147] : 
                      (N30)? piso_data_r[211] : 
                      (N25)? piso_data_r[275] : 
                      (N27)? piso_data_r[339] : 
                      (N29)? piso_data_r[403] : 
                      (N31)? piso_data_r[467] : 1'b0;
  assign data_o[18] = (N24)? piso_data_r[18] : 
                      (N26)? piso_data_r[82] : 
                      (N28)? piso_data_r[146] : 
                      (N30)? piso_data_r[210] : 
                      (N25)? piso_data_r[274] : 
                      (N27)? piso_data_r[338] : 
                      (N29)? piso_data_r[402] : 
                      (N31)? piso_data_r[466] : 1'b0;
  assign data_o[17] = (N24)? piso_data_r[17] : 
                      (N26)? piso_data_r[81] : 
                      (N28)? piso_data_r[145] : 
                      (N30)? piso_data_r[209] : 
                      (N25)? piso_data_r[273] : 
                      (N27)? piso_data_r[337] : 
                      (N29)? piso_data_r[401] : 
                      (N31)? piso_data_r[465] : 1'b0;
  assign data_o[16] = (N24)? piso_data_r[16] : 
                      (N26)? piso_data_r[80] : 
                      (N28)? piso_data_r[144] : 
                      (N30)? piso_data_r[208] : 
                      (N25)? piso_data_r[272] : 
                      (N27)? piso_data_r[336] : 
                      (N29)? piso_data_r[400] : 
                      (N31)? piso_data_r[464] : 1'b0;
  assign data_o[15] = (N24)? piso_data_r[15] : 
                      (N26)? piso_data_r[79] : 
                      (N28)? piso_data_r[143] : 
                      (N30)? piso_data_r[207] : 
                      (N25)? piso_data_r[271] : 
                      (N27)? piso_data_r[335] : 
                      (N29)? piso_data_r[399] : 
                      (N31)? piso_data_r[463] : 1'b0;
  assign data_o[14] = (N24)? piso_data_r[14] : 
                      (N26)? piso_data_r[78] : 
                      (N28)? piso_data_r[142] : 
                      (N30)? piso_data_r[206] : 
                      (N25)? piso_data_r[270] : 
                      (N27)? piso_data_r[334] : 
                      (N29)? piso_data_r[398] : 
                      (N31)? piso_data_r[462] : 1'b0;
  assign data_o[13] = (N24)? piso_data_r[13] : 
                      (N26)? piso_data_r[77] : 
                      (N28)? piso_data_r[141] : 
                      (N30)? piso_data_r[205] : 
                      (N25)? piso_data_r[269] : 
                      (N27)? piso_data_r[333] : 
                      (N29)? piso_data_r[397] : 
                      (N31)? piso_data_r[461] : 1'b0;
  assign data_o[12] = (N24)? piso_data_r[12] : 
                      (N26)? piso_data_r[76] : 
                      (N28)? piso_data_r[140] : 
                      (N30)? piso_data_r[204] : 
                      (N25)? piso_data_r[268] : 
                      (N27)? piso_data_r[332] : 
                      (N29)? piso_data_r[396] : 
                      (N31)? piso_data_r[460] : 1'b0;
  assign data_o[11] = (N24)? piso_data_r[11] : 
                      (N26)? piso_data_r[75] : 
                      (N28)? piso_data_r[139] : 
                      (N30)? piso_data_r[203] : 
                      (N25)? piso_data_r[267] : 
                      (N27)? piso_data_r[331] : 
                      (N29)? piso_data_r[395] : 
                      (N31)? piso_data_r[459] : 1'b0;
  assign data_o[10] = (N24)? piso_data_r[10] : 
                      (N26)? piso_data_r[74] : 
                      (N28)? piso_data_r[138] : 
                      (N30)? piso_data_r[202] : 
                      (N25)? piso_data_r[266] : 
                      (N27)? piso_data_r[330] : 
                      (N29)? piso_data_r[394] : 
                      (N31)? piso_data_r[458] : 1'b0;
  assign data_o[9] = (N24)? piso_data_r[9] : 
                     (N26)? piso_data_r[73] : 
                     (N28)? piso_data_r[137] : 
                     (N30)? piso_data_r[201] : 
                     (N25)? piso_data_r[265] : 
                     (N27)? piso_data_r[329] : 
                     (N29)? piso_data_r[393] : 
                     (N31)? piso_data_r[457] : 1'b0;
  assign data_o[8] = (N24)? piso_data_r[8] : 
                     (N26)? piso_data_r[72] : 
                     (N28)? piso_data_r[136] : 
                     (N30)? piso_data_r[200] : 
                     (N25)? piso_data_r[264] : 
                     (N27)? piso_data_r[328] : 
                     (N29)? piso_data_r[392] : 
                     (N31)? piso_data_r[456] : 1'b0;
  assign data_o[7] = (N24)? piso_data_r[7] : 
                     (N26)? piso_data_r[71] : 
                     (N28)? piso_data_r[135] : 
                     (N30)? piso_data_r[199] : 
                     (N25)? piso_data_r[263] : 
                     (N27)? piso_data_r[327] : 
                     (N29)? piso_data_r[391] : 
                     (N31)? piso_data_r[455] : 1'b0;
  assign data_o[6] = (N24)? piso_data_r[6] : 
                     (N26)? piso_data_r[70] : 
                     (N28)? piso_data_r[134] : 
                     (N30)? piso_data_r[198] : 
                     (N25)? piso_data_r[262] : 
                     (N27)? piso_data_r[326] : 
                     (N29)? piso_data_r[390] : 
                     (N31)? piso_data_r[454] : 1'b0;
  assign data_o[5] = (N24)? piso_data_r[5] : 
                     (N26)? piso_data_r[69] : 
                     (N28)? piso_data_r[133] : 
                     (N30)? piso_data_r[197] : 
                     (N25)? piso_data_r[261] : 
                     (N27)? piso_data_r[325] : 
                     (N29)? piso_data_r[389] : 
                     (N31)? piso_data_r[453] : 1'b0;
  assign data_o[4] = (N24)? piso_data_r[4] : 
                     (N26)? piso_data_r[68] : 
                     (N28)? piso_data_r[132] : 
                     (N30)? piso_data_r[196] : 
                     (N25)? piso_data_r[260] : 
                     (N27)? piso_data_r[324] : 
                     (N29)? piso_data_r[388] : 
                     (N31)? piso_data_r[452] : 1'b0;
  assign data_o[3] = (N24)? piso_data_r[3] : 
                     (N26)? piso_data_r[67] : 
                     (N28)? piso_data_r[131] : 
                     (N30)? piso_data_r[195] : 
                     (N25)? piso_data_r[259] : 
                     (N27)? piso_data_r[323] : 
                     (N29)? piso_data_r[387] : 
                     (N31)? piso_data_r[451] : 1'b0;
  assign data_o[2] = (N24)? piso_data_r[2] : 
                     (N26)? piso_data_r[66] : 
                     (N28)? piso_data_r[130] : 
                     (N30)? piso_data_r[194] : 
                     (N25)? piso_data_r[258] : 
                     (N27)? piso_data_r[322] : 
                     (N29)? piso_data_r[386] : 
                     (N31)? piso_data_r[450] : 1'b0;
  assign data_o[1] = (N24)? piso_data_r[1] : 
                     (N26)? piso_data_r[65] : 
                     (N28)? piso_data_r[129] : 
                     (N30)? piso_data_r[193] : 
                     (N25)? piso_data_r[257] : 
                     (N27)? piso_data_r[321] : 
                     (N29)? piso_data_r[385] : 
                     (N31)? piso_data_r[449] : 1'b0;
  assign data_o[0] = (N24)? piso_data_r[0] : 
                     (N26)? piso_data_r[64] : 
                     (N28)? piso_data_r[128] : 
                     (N30)? piso_data_r[192] : 
                     (N25)? piso_data_r[256] : 
                     (N27)? piso_data_r[320] : 
                     (N29)? piso_data_r[384] : 
                     (N31)? piso_data_r[448] : 1'b0;
  assign N34 = ~valid_o;
  assign N35 = piso_shift_ctr_r[1] & piso_shift_ctr_r[2];
  assign N36 = piso_shift_ctr_r[0] & N35;
  assign { N16, N15, N14 } = piso_shift_ctr_r + 1'b1;
  assign piso_state_n[0] = (N0)? 1'b1 : 
                           (N5)? 1'b0 : 1'b0;
  assign N0 = N2;
  assign { N11, N10, N9 } = (N1)? { 1'b0, 1'b0, 1'b0 } : 
                            (N8)? { N16, N15, N14 } : 1'b0;
  assign N1 = N7;
  assign piso_done_tx_n = N37 & yumi_i;
  assign N37 = valid_o & N36;
  assign ready_o = N34 | piso_done_tx_n;
  assign N2 = ready_o & valid_i;
  assign N3 = piso_done_tx_n | N2;
  assign N4 = ~N2;
  assign N5 = piso_done_tx_n & N4;
  assign N6 = ready_o & valid_i;
  assign N7 = ready_o & valid_i;
  assign N8 = ~N7;
  assign N12 = N38 & N39;
  assign N38 = valid_o & yumi_i;
  assign N39 = ~piso_done_tx_n;
  assign N13 = ~N12;
  assign N17 = ~piso_shift_ctr_r[0];
  assign N18 = ~piso_shift_ctr_r[1];
  assign N19 = N17 & N18;
  assign N20 = N17 & piso_shift_ctr_r[1];
  assign N21 = piso_shift_ctr_r[0] & N18;
  assign N22 = piso_shift_ctr_r[0] & piso_shift_ctr_r[1];
  assign N23 = ~piso_shift_ctr_r[2];
  assign N24 = N19 & N23;
  assign N25 = N19 & piso_shift_ctr_r[2];
  assign N26 = N21 & N23;
  assign N27 = N21 & piso_shift_ctr_r[2];
  assign N28 = N20 & N23;
  assign N29 = N20 & piso_shift_ctr_r[2];
  assign N30 = N22 & N23;
  assign N31 = N22 & piso_shift_ctr_r[2];
  assign N32 = N13 & N8;
  assign N33 = ~N32;

endmodule