module xics_ics_16_3(clk, rst, \wb_in.adr , \wb_in.dat , \wb_in.sel , \wb_in.cyc , \wb_in.stb , \wb_in.we , int_level_in, \wb_out.dat , \wb_out.ack , \wb_out.stall , \icp_out.src , \icp_out.pri );
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire [2:0] _0010_;
  wire [2:0] _0011_;
  wire [2:0] _0012_;
  wire [2:0] _0013_;
  wire [2:0] _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire [2:0] _0025_;
  wire [2:0] _0026_;
  wire [2:0] _0027_;
  wire [2:0] _0028_;
  wire [2:0] _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  reg [15:0] _0034_;
  wire _0035_;
  wire [3:0] _0036_;
  wire _0037_;
  wire [7:0] _0038_;
  wire [31:0] _0039_;
  wire [31:0] _0040_;
  wire [31:0] _0041_;
  reg [32:0] _0042_;
  wire _0043_;
  wire [3:0] _0044_;
  wire _0045_;
  wire [2:0] _0046_;
  wire [47:0] _0047_;
  wire [47:0] _0048_;
  reg [47:0] _0049_;
  reg [11:0] _0050_;
  wire [7:0] _0051_;
  wire [7:0] _0052_;
  wire [7:0] _0053_;
  wire [7:0] _0054_;
  wire [7:0] _0055_;
  wire [7:0] _0056_;
  wire [7:0] _0057_;
  wire [7:0] _0058_;
  wire [7:0] _0059_;
  wire [7:0] _0060_;
  wire [7:0] _0061_;
  wire [7:0] _0062_;
  wire [7:0] _0063_;
  wire [7:0] _0064_;
  wire [7:0] _0065_;
  wire [7:0] _0066_;
  wire [7:0] _0067_;
  wire [7:0] _0068_;
  wire [7:0] _0069_;
  wire [7:0] _0070_;
  wire [7:0] _0071_;
  wire [7:0] _0072_;
  wire [7:0] _0073_;
  wire [7:0] _0074_;
  wire [7:0] _0075_;
  wire [7:0] _0076_;
  wire [7:0] _0077_;
  wire [7:0] _0078_;
  wire [7:0] _0079_;
  wire [7:0] _0080_;
  wire [7:0] _0081_;
  wire [6:0] _0082_;
  wire [6:0] _0083_;
  wire [6:0] _0084_;
  wire [6:0] _0085_;
  wire [6:0] _0086_;
  wire [6:0] _0087_;
  wire [6:0] _0088_;
  wire [6:0] _0089_;
  wire [6:0] _0090_;
  wire [6:0] _0091_;
  wire [6:0] _0092_;
  wire [6:0] _0093_;
  wire [6:0] _0094_;
  wire [6:0] _0095_;
  wire [6:0] _0096_;
  wire [6:0] _0097_;
  wire [7:0] _0098_;
  wire [7:0] _0099_;
  wire [7:0] _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire [15:0] _0464_;
  wire [15:0] _0465_;
  wire [15:0] _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire [7:0] _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire [2:0] _0794_;
  wire [2:0] _0795_;
  wire [2:0] _0796_;
  wire [2:0] _0797_;
  wire [2:0] _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire [2:0] _0832_;
  wire _0833_;
  wire [2:0] _0834_;
  wire _0835_;
  wire [2:0] _0836_;
  wire _0837_;
  wire [2:0] _0838_;
  wire _0839_;
  wire [2:0] _0840_;
  wire _0841_;
  wire [2:0] _0842_;
  wire _0843_;
  wire [2:0] _0844_;
  wire _0845_;
  wire [2:0] _0846_;
  wire _0847_;
  wire [2:0] _0848_;
  wire _0849_;
  wire [2:0] _0850_;
  wire _0851_;
  wire [2:0] _0852_;
  wire _0853_;
  wire [2:0] _0854_;
  wire _0855_;
  wire [2:0] _0856_;
  wire _0857_;
  wire [2:0] _0858_;
  wire _0859_;
  wire [2:0] _0860_;
  wire _0861_;
  wire [2:0] _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  input clk;
  wire clk;
  output [7:0] \icp_out.pri ;
  wire [7:0] \icp_out.pri ;
  output [3:0] \icp_out.src ;
  wire [3:0] \icp_out.src ;
  wire [11:0] icp_out_next;
  input [15:0] int_level_in;
  wire [15:0] int_level_in;
  wire [15:0] int_level_l;
  wire [3:0] reg_idx;
  wire reg_is_config;
  wire reg_is_debug;
  wire reg_is_xive;
  input rst;
  wire rst;
  input [29:0] \wb_in.adr ;
  wire [29:0] \wb_in.adr ;
  input \wb_in.cyc ;
  wire \wb_in.cyc ;
  input [31:0] \wb_in.dat ;
  wire [31:0] \wb_in.dat ;
  input [3:0] \wb_in.sel ;
  wire [3:0] \wb_in.sel ;
  input \wb_in.stb ;
  wire \wb_in.stb ;
  input \wb_in.we ;
  wire \wb_in.we ;
  output \wb_out.ack ;
  wire \wb_out.ack ;
  output [31:0] \wb_out.dat ;
  wire [31:0] \wb_out.dat ;
  output \wb_out.stall ;
  wire \wb_out.stall ;
  wire wb_valid;
  wire [47:0] xives;
  assign _0000_ = reg_idx[0] ? int_level_l[1] : int_level_l[0];
  assign _0001_ = reg_idx[0] ? int_level_l[5] : int_level_l[4];
  assign _0002_ = reg_idx[0] ? int_level_l[9] : int_level_l[8];
  assign _0003_ = reg_idx[0] ? int_level_l[13] : int_level_l[12];
  assign _0004_ = reg_idx[2] ? _0785_ : _0784_;
  assign _0005_ = reg_idx[0] ? int_level_l[1] : int_level_l[0];
  assign _0006_ = reg_idx[0] ? int_level_l[5] : int_level_l[4];
  assign _0007_ = reg_idx[0] ? int_level_l[9] : int_level_l[8];
  assign _0008_ = reg_idx[0] ? int_level_l[13] : int_level_l[12];
  assign _0009_ = reg_idx[2] ? _0790_ : _0789_;
  assign _0010_ = _0036_[0] ? xives[5:3] : xives[2:0];
  assign _0011_ = _0036_[0] ? xives[17:15] : xives[14:12];
  assign _0012_ = _0036_[0] ? xives[29:27] : xives[26:24];
  assign _0013_ = _0036_[0] ? xives[41:39] : xives[38:36];
  assign _0014_ = _0036_[2] ? _0795_ : _0794_;
  assign _0015_ = reg_idx[0] ? int_level_l[3] : int_level_l[2];
  assign _0016_ = reg_idx[0] ? int_level_l[7] : int_level_l[6];
  assign _0017_ = reg_idx[0] ? int_level_l[11] : int_level_l[10];
  assign _0018_ = reg_idx[0] ? int_level_l[15] : int_level_l[14];
  assign _0019_ = reg_idx[2] ? _0787_ : _0786_;
  assign _0020_ = reg_idx[0] ? int_level_l[3] : int_level_l[2];
  assign _0021_ = reg_idx[0] ? int_level_l[7] : int_level_l[6];
  assign _0022_ = reg_idx[0] ? int_level_l[11] : int_level_l[10];
  assign _0023_ = reg_idx[0] ? int_level_l[15] : int_level_l[14];
  assign _0024_ = reg_idx[2] ? _0792_ : _0791_;
  assign _0025_ = _0036_[0] ? xives[11:9] : xives[8:6];
  assign _0026_ = _0036_[0] ? xives[23:21] : xives[20:18];
  assign _0027_ = _0036_[0] ? xives[35:33] : xives[32:30];
  assign _0028_ = _0036_[0] ? xives[47:45] : xives[44:42];
  assign _0029_ = _0036_[2] ? _0797_ : _0796_;
  assign _0784_ = reg_idx[1] ? _0015_ : _0000_;
  assign _0785_ = reg_idx[1] ? _0016_ : _0001_;
  assign _0786_ = reg_idx[1] ? _0017_ : _0002_;
  assign _0787_ = reg_idx[1] ? _0018_ : _0003_;
  assign _0788_ = reg_idx[3] ? _0019_ : _0004_;
  assign _0789_ = reg_idx[1] ? _0020_ : _0005_;
  assign _0790_ = reg_idx[1] ? _0021_ : _0006_;
  assign _0791_ = reg_idx[1] ? _0022_ : _0007_;
  assign _0792_ = reg_idx[1] ? _0023_ : _0008_;
  assign _0793_ = reg_idx[3] ? _0024_ : _0009_;
  assign _0794_ = _0036_[1] ? _0025_ : _0010_;
  assign _0795_ = _0036_[1] ? _0026_ : _0011_;
  assign _0796_ = _0036_[1] ? _0027_ : _0012_;
  assign _0797_ = _0036_[1] ? _0028_ : _0013_;
  assign _0798_ = _0036_[3] ? _0029_ : _0014_;
  assign _0030_ = \wb_in.adr [9:0] == 10'h000;
  assign _0031_ = _0030_ ? 1'h1 : 1'h0;
  assign _0032_ = \wb_in.adr [9:0] == 10'h001;
  assign _0033_ = _0032_ ? 1'h1 : 1'h0;
  always @(posedge clk)
    _0034_ <= int_level_in;
  assign _0035_ = \wb_in.cyc  & \wb_in.stb ;
  assign _0036_ = 4'hf - reg_idx;
  assign _0037_ = _0798_ == 3'h7;
  assign _0038_ = _0037_ ? 8'hff : { 5'h00, _0798_ };
  assign _0039_ = reg_is_debug ? { 20'h00000, icp_out_next[3:0], icp_out_next[11:4] } : 32'd0;
  assign _0040_ = reg_is_config ? 32'd50331664 : _0039_;
  assign _0041_ = reg_is_xive ? { _0788_, 1'h0, _0793_, 21'h000000, _0038_ } : _0040_;
  always @(posedge clk)
    _0042_ <= { wb_valid, _0041_[7:0], _0041_[15:8], _0041_[23:16], _0041_[31:24] };
  assign _0043_ = wb_valid & \wb_in.we ;
  assign _0044_ = 4'hf - reg_idx;
  assign _0045_ = \wb_in.dat [31:24] >= 8'h07;
  assign _0046_ = _0045_ ? 3'h7 : \wb_in.dat [26:24];
  assign _0047_ = _0043_ ? { _0862_, _0860_, _0858_, _0856_, _0854_, _0852_, _0850_, _0848_, _0846_, _0844_, _0842_, _0840_, _0838_, _0836_, _0834_, _0832_ } : xives;
  assign _0048_ = rst ? 48'hffffffffffff : _0047_;
  always @(posedge clk)
    _0049_ <= _0048_;
  always @(posedge clk)
    _0050_ <= icp_out_next;
  assign _0051_ = 8'h00 | { _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_ };
  assign _0052_ = int_level_l[0] ? _0051_ : 8'h00;
  assign _0053_ = _0052_ | { _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_ };
  assign _0054_ = int_level_l[1] ? _0053_ : _0052_;
  assign _0055_ = _0054_ | { _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_ };
  assign _0056_ = int_level_l[2] ? _0055_ : _0054_;
  assign _0057_ = _0056_ | { _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_ };
  assign _0058_ = int_level_l[3] ? _0057_ : _0056_;
  assign _0059_ = _0058_ | { _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_ };
  assign _0060_ = int_level_l[4] ? _0059_ : _0058_;
  assign _0061_ = _0060_ | { _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_ };
  assign _0062_ = int_level_l[5] ? _0061_ : _0060_;
  assign _0063_ = _0062_ | { _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_ };
  assign _0064_ = int_level_l[6] ? _0063_ : _0062_;
  assign _0065_ = _0064_ | { _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_ };
  assign _0066_ = int_level_l[7] ? _0065_ : _0064_;
  assign _0067_ = _0066_ | { _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_ };
  assign _0068_ = int_level_l[8] ? _0067_ : _0066_;
  assign _0069_ = _0068_ | { _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_ };
  assign _0070_ = int_level_l[9] ? _0069_ : _0068_;
  assign _0071_ = _0070_ | { _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_ };
  assign _0072_ = int_level_l[10] ? _0071_ : _0070_;
  assign _0073_ = _0072_ | { _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_ };
  assign _0074_ = int_level_l[11] ? _0073_ : _0072_;
  assign _0075_ = _0074_ | { _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_ };
  assign _0076_ = int_level_l[12] ? _0075_ : _0074_;
  assign _0077_ = _0076_ | { _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_ };
  assign _0078_ = int_level_l[13] ? _0077_ : _0076_;
  assign _0079_ = _0078_ | { _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_ };
  assign _0080_ = int_level_l[14] ? _0079_ : _0078_;
  assign _0081_ = _0080_ | { _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_ };
  assign _0082_ = int_level_l[0] ? _0051_[6:0] : 7'h00;
  assign _0083_ = int_level_l[1] ? _0053_[6:0] : _0082_;
  assign _0084_ = int_level_l[2] ? _0055_[6:0] : _0083_;
  assign _0085_ = int_level_l[3] ? _0057_[6:0] : _0084_;
  assign _0086_ = int_level_l[4] ? _0059_[6:0] : _0085_;
  assign _0087_ = int_level_l[5] ? _0061_[6:0] : _0086_;
  assign _0088_ = int_level_l[6] ? _0063_[6:0] : _0087_;
  assign _0089_ = int_level_l[7] ? _0065_[6:0] : _0088_;
  assign _0090_ = int_level_l[8] ? _0067_[6:0] : _0089_;
  assign _0091_ = int_level_l[9] ? _0069_[6:0] : _0090_;
  assign _0092_ = int_level_l[10] ? _0071_[6:0] : _0091_;
  assign _0093_ = int_level_l[11] ? _0073_[6:0] : _0092_;
  assign _0094_ = int_level_l[12] ? _0075_[6:0] : _0093_;
  assign _0095_ = int_level_l[13] ? _0077_[6:0] : _0094_;
  assign _0096_ = int_level_l[14] ? _0079_[6:0] : _0095_;
  assign _0097_ = int_level_l[15] ? _0081_[6:0] : _0096_;
  assign _0098_ = - $signed({ 1'h1, _0097_ });
  assign _0099_ = _0098_ & { 1'h1, _0097_ };
  assign _0100_ = _0098_ | { 1'h1, _0097_ };
  assign _0101_ = ~ _0100_[0];
  assign _0102_ = _0100_[1] & _0101_;
  assign _0103_ = 1'h0 | _0102_;
  assign _0104_ = ~ _0100_[2];
  assign _0105_ = _0100_[3] & _0104_;
  assign _0106_ = _0103_ | _0105_;
  assign _0107_ = ~ _0100_[4];
  assign _0108_ = _0100_[5] & _0107_;
  assign _0109_ = _0106_ | _0108_;
  assign _0110_ = ~ _0100_[6];
  assign _0111_ = _0100_[7] & _0110_;
  assign _0112_ = _0109_ | _0111_;
  assign _0113_ = ~ _0100_[7];
  assign _0114_ = _0100_[7] & _0113_;
  assign _0115_ = _0112_ | _0114_;
  assign _0116_ = ~ _0100_[7];
  assign _0117_ = _0100_[7] & _0116_;
  assign _0118_ = _0115_ | _0117_;
  assign _0119_ = ~ _0100_[7];
  assign _0120_ = _0100_[7] & _0119_;
  assign _0121_ = _0118_ | _0120_;
  assign _0122_ = ~ _0100_[7];
  assign _0123_ = _0100_[7] & _0122_;
  assign _0124_ = _0121_ | _0123_;
  assign _0125_ = ~ _0100_[7];
  assign _0126_ = _0100_[7] & _0125_;
  assign _0127_ = _0124_ | _0126_;
  assign _0128_ = ~ _0100_[7];
  assign _0129_ = _0100_[7] & _0128_;
  assign _0130_ = _0127_ | _0129_;
  assign _0131_ = ~ _0100_[7];
  assign _0132_ = _0100_[7] & _0131_;
  assign _0133_ = _0130_ | _0132_;
  assign _0134_ = ~ _0100_[7];
  assign _0135_ = _0100_[7] & _0134_;
  assign _0136_ = _0133_ | _0135_;
  assign _0137_ = ~ _0100_[7];
  assign _0138_ = _0100_[7] & _0137_;
  assign _0139_ = _0136_ | _0138_;
  assign _0140_ = ~ _0100_[7];
  assign _0141_ = _0100_[7] & _0140_;
  assign _0142_ = _0139_ | _0141_;
  assign _0143_ = ~ _0100_[7];
  assign _0144_ = _0100_[7] & _0143_;
  assign _0145_ = _0142_ | _0144_;
  assign _0146_ = ~ _0100_[7];
  assign _0147_ = _0100_[7] & _0146_;
  assign _0148_ = _0145_ | _0147_;
  assign _0149_ = ~ _0100_[7];
  assign _0150_ = _0100_[7] & _0149_;
  assign _0151_ = _0148_ | _0150_;
  assign _0152_ = ~ _0100_[7];
  assign _0153_ = _0100_[7] & _0152_;
  assign _0154_ = _0151_ | _0153_;
  assign _0155_ = ~ _0100_[7];
  assign _0156_ = _0100_[7] & _0155_;
  assign _0157_ = _0154_ | _0156_;
  assign _0158_ = ~ _0100_[7];
  assign _0159_ = _0100_[7] & _0158_;
  assign _0160_ = _0157_ | _0159_;
  assign _0161_ = ~ _0100_[7];
  assign _0162_ = _0100_[7] & _0161_;
  assign _0163_ = _0160_ | _0162_;
  assign _0164_ = ~ _0100_[7];
  assign _0165_ = _0100_[7] & _0164_;
  assign _0166_ = _0163_ | _0165_;
  assign _0167_ = ~ _0100_[7];
  assign _0168_ = _0100_[7] & _0167_;
  assign _0169_ = _0166_ | _0168_;
  assign _0170_ = ~ _0100_[7];
  assign _0171_ = _0100_[7] & _0170_;
  assign _0172_ = _0169_ | _0171_;
  assign _0173_ = ~ _0100_[7];
  assign _0174_ = _0100_[7] & _0173_;
  assign _0175_ = _0172_ | _0174_;
  assign _0176_ = ~ _0100_[7];
  assign _0177_ = _0100_[7] & _0176_;
  assign _0178_ = _0175_ | _0177_;
  assign _0179_ = ~ _0100_[7];
  assign _0180_ = _0100_[7] & _0179_;
  assign _0181_ = _0178_ | _0180_;
  assign _0182_ = ~ _0100_[7];
  assign _0183_ = _0100_[7] & _0182_;
  assign _0184_ = _0181_ | _0183_;
  assign _0185_ = ~ _0100_[7];
  assign _0186_ = _0100_[7] & _0185_;
  assign _0187_ = _0184_ | _0186_;
  assign _0188_ = ~ _0100_[7];
  assign _0189_ = _0100_[7] & _0188_;
  assign _0190_ = _0187_ | _0189_;
  assign _0191_ = ~ _0100_[7];
  assign _0192_ = _0100_[7] & _0191_;
  assign _0193_ = _0190_ | _0192_;
  assign _0194_ = ~ _0100_[7];
  assign _0195_ = _0100_[7] & _0194_;
  assign _0196_ = _0193_ | _0195_;
  assign _0197_ = ~ _0100_[1];
  assign _0198_ = _0100_[3] & _0197_;
  assign _0199_ = 1'h0 | _0198_;
  assign _0200_ = ~ _0100_[5];
  assign _0201_ = _0100_[7] & _0200_;
  assign _0202_ = _0199_ | _0201_;
  assign _0203_ = ~ _0100_[7];
  assign _0204_ = _0100_[7] & _0203_;
  assign _0205_ = _0202_ | _0204_;
  assign _0206_ = ~ _0100_[7];
  assign _0207_ = _0100_[7] & _0206_;
  assign _0208_ = _0205_ | _0207_;
  assign _0209_ = ~ _0100_[7];
  assign _0210_ = _0100_[7] & _0209_;
  assign _0211_ = _0208_ | _0210_;
  assign _0212_ = ~ _0100_[7];
  assign _0213_ = _0100_[7] & _0212_;
  assign _0214_ = _0211_ | _0213_;
  assign _0215_ = ~ _0100_[7];
  assign _0216_ = _0100_[7] & _0215_;
  assign _0217_ = _0214_ | _0216_;
  assign _0218_ = ~ _0100_[7];
  assign _0219_ = _0100_[7] & _0218_;
  assign _0220_ = _0217_ | _0219_;
  assign _0221_ = ~ _0100_[7];
  assign _0222_ = _0100_[7] & _0221_;
  assign _0223_ = _0220_ | _0222_;
  assign _0224_ = ~ _0100_[7];
  assign _0225_ = _0100_[7] & _0224_;
  assign _0226_ = _0223_ | _0225_;
  assign _0227_ = ~ _0100_[7];
  assign _0228_ = _0100_[7] & _0227_;
  assign _0229_ = _0226_ | _0228_;
  assign _0230_ = ~ _0100_[7];
  assign _0231_ = _0100_[7] & _0230_;
  assign _0232_ = _0229_ | _0231_;
  assign _0233_ = ~ _0100_[7];
  assign _0234_ = _0100_[7] & _0233_;
  assign _0235_ = _0232_ | _0234_;
  assign _0236_ = ~ _0100_[7];
  assign _0237_ = _0100_[7] & _0236_;
  assign _0238_ = _0235_ | _0237_;
  assign _0239_ = ~ _0100_[7];
  assign _0240_ = _0100_[7] & _0239_;
  assign _0241_ = _0238_ | _0240_;
  assign _0242_ = ~ _0100_[7];
  assign _0243_ = _0100_[7] & _0242_;
  assign _0244_ = _0241_ | _0243_;
  assign _0245_ = ~ _0100_[3];
  assign _0246_ = _0100_[7] & _0245_;
  assign _0247_ = 1'h0 | _0246_;
  assign _0248_ = ~ _0100_[7];
  assign _0249_ = _0100_[7] & _0248_;
  assign _0250_ = _0247_ | _0249_;
  assign _0251_ = ~ _0100_[7];
  assign _0252_ = _0100_[7] & _0251_;
  assign _0253_ = _0250_ | _0252_;
  assign _0254_ = ~ _0100_[7];
  assign _0255_ = _0100_[7] & _0254_;
  assign _0256_ = _0253_ | _0255_;
  assign _0257_ = ~ _0100_[7];
  assign _0258_ = _0100_[7] & _0257_;
  assign _0259_ = _0256_ | _0258_;
  assign _0260_ = ~ _0100_[7];
  assign _0261_ = _0100_[7] & _0260_;
  assign _0262_ = _0259_ | _0261_;
  assign _0263_ = ~ _0100_[7];
  assign _0264_ = _0100_[7] & _0263_;
  assign _0265_ = _0262_ | _0264_;
  assign _0266_ = ~ _0100_[7];
  assign _0267_ = _0100_[7] & _0266_;
  assign _0268_ = _0265_ | _0267_;
  assign _0269_ = ~ _0100_[7];
  assign _0270_ = _0100_[7] & _0269_;
  assign _0271_ = 1'h0 | _0270_;
  assign _0272_ = ~ _0100_[7];
  assign _0273_ = _0100_[7] & _0272_;
  assign _0274_ = _0271_ | _0273_;
  assign _0275_ = ~ _0100_[7];
  assign _0276_ = _0100_[7] & _0275_;
  assign _0277_ = _0274_ | _0276_;
  assign _0278_ = ~ _0100_[7];
  assign _0279_ = _0100_[7] & _0278_;
  assign _0280_ = _0277_ | _0279_;
  assign _0281_ = ~ _0100_[7];
  assign _0282_ = _0100_[7] & _0281_;
  assign _0283_ = 1'h0 | _0282_;
  assign _0284_ = ~ _0100_[7];
  assign _0285_ = _0100_[7] & _0284_;
  assign _0286_ = _0283_ | _0285_;
  assign _0287_ = ~ _0100_[7];
  assign _0288_ = _0100_[7] & _0287_;
  assign _0289_ = 1'h0 | _0288_;
  assign _0290_ = | _0099_[1];
  assign _0291_ = 1'h0 | _0290_;
  assign _0292_ = | _0099_[3];
  assign _0293_ = _0291_ | _0292_;
  assign _0294_ = | _0099_[5];
  assign _0295_ = _0293_ | _0294_;
  assign _0296_ = | _0099_[7];
  assign _0297_ = _0295_ | _0296_;
  assign _0298_ = | 1'h0;
  assign _0299_ = _0297_ | _0298_;
  assign _0300_ = | 1'h0;
  assign _0301_ = _0299_ | _0300_;
  assign _0302_ = | 1'h0;
  assign _0303_ = _0301_ | _0302_;
  assign _0304_ = | 1'h0;
  assign _0305_ = _0303_ | _0304_;
  assign _0306_ = | 1'h0;
  assign _0307_ = _0305_ | _0306_;
  assign _0308_ = | 1'h0;
  assign _0309_ = _0307_ | _0308_;
  assign _0310_ = | 1'h0;
  assign _0311_ = _0309_ | _0310_;
  assign _0312_ = | 1'h0;
  assign _0313_ = _0311_ | _0312_;
  assign _0314_ = | 1'h0;
  assign _0315_ = _0313_ | _0314_;
  assign _0316_ = | 1'h0;
  assign _0317_ = _0315_ | _0316_;
  assign _0318_ = | 1'h0;
  assign _0319_ = _0317_ | _0318_;
  assign _0320_ = | 1'h0;
  assign _0321_ = _0319_ | _0320_;
  assign _0322_ = | 1'h0;
  assign _0323_ = _0321_ | _0322_;
  assign _0324_ = | 1'h0;
  assign _0325_ = _0323_ | _0324_;
  assign _0326_ = | 1'h0;
  assign _0327_ = _0325_ | _0326_;
  assign _0328_ = | 1'h0;
  assign _0329_ = _0327_ | _0328_;
  assign _0330_ = | 1'h0;
  assign _0331_ = _0329_ | _0330_;
  assign _0332_ = | 1'h0;
  assign _0333_ = _0331_ | _0332_;
  assign _0334_ = | 1'h0;
  assign _0335_ = _0333_ | _0334_;
  assign _0336_ = | 1'h0;
  assign _0337_ = _0335_ | _0336_;
  assign _0338_ = | 1'h0;
  assign _0339_ = _0337_ | _0338_;
  assign _0340_ = | 1'h0;
  assign _0341_ = _0339_ | _0340_;
  assign _0342_ = | 1'h0;
  assign _0343_ = _0341_ | _0342_;
  assign _0344_ = | 1'h0;
  assign _0345_ = _0343_ | _0344_;
  assign _0346_ = | 1'h0;
  assign _0347_ = _0345_ | _0346_;
  assign _0348_ = | 1'h0;
  assign _0349_ = _0347_ | _0348_;
  assign _0350_ = | 1'h0;
  assign _0351_ = _0349_ | _0350_;
  assign _0352_ = | 1'h0;
  assign _0353_ = _0351_ | _0352_;
  assign _0354_ = | _0099_[3:2];
  assign _0355_ = 1'h0 | _0354_;
  assign _0356_ = | _0099_[7:6];
  assign _0357_ = _0355_ | _0356_;
  assign _0358_ = | 2'h0;
  assign _0359_ = _0357_ | _0358_;
  assign _0360_ = | 2'h0;
  assign _0361_ = _0359_ | _0360_;
  assign _0362_ = | 2'h0;
  assign _0363_ = _0361_ | _0362_;
  assign _0364_ = | 2'h0;
  assign _0365_ = _0363_ | _0364_;
  assign _0366_ = | 2'h0;
  assign _0367_ = _0365_ | _0366_;
  assign _0368_ = | 2'h0;
  assign _0369_ = _0367_ | _0368_;
  assign _0370_ = | 2'h0;
  assign _0371_ = _0369_ | _0370_;
  assign _0372_ = | 2'h0;
  assign _0373_ = _0371_ | _0372_;
  assign _0374_ = | 2'h0;
  assign _0375_ = _0373_ | _0374_;
  assign _0376_ = | 2'h0;
  assign _0377_ = _0375_ | _0376_;
  assign _0378_ = | 2'h0;
  assign _0379_ = _0377_ | _0378_;
  assign _0380_ = | 2'h0;
  assign _0381_ = _0379_ | _0380_;
  assign _0382_ = | 2'h0;
  assign _0383_ = _0381_ | _0382_;
  assign _0384_ = | 2'h0;
  assign _0385_ = _0383_ | _0384_;
  assign _0386_ = | _0099_[7:4];
  assign _0387_ = 1'h0 | _0386_;
  assign _0388_ = | 4'h0;
  assign _0389_ = _0387_ | _0388_;
  assign _0390_ = | 4'h0;
  assign _0391_ = _0389_ | _0390_;
  assign _0392_ = | 4'h0;
  assign _0393_ = _0391_ | _0392_;
  assign _0394_ = | 4'h0;
  assign _0395_ = _0393_ | _0394_;
  assign _0396_ = | 4'h0;
  assign _0397_ = _0395_ | _0396_;
  assign _0398_ = | 4'h0;
  assign _0399_ = _0397_ | _0398_;
  assign _0400_ = | 4'h0;
  assign _0401_ = _0399_ | _0400_;
  assign _0402_ = | 8'h00;
  assign _0403_ = 1'h0 | _0402_;
  assign _0404_ = | 8'h00;
  assign _0405_ = _0403_ | _0404_;
  assign _0406_ = | 8'h00;
  assign _0407_ = _0405_ | _0406_;
  assign _0408_ = | 8'h00;
  assign _0409_ = _0407_ | _0408_;
  assign _0410_ = | 16'h0000;
  assign _0411_ = 1'h0 | _0410_;
  assign _0412_ = | 16'h0000;
  assign _0413_ = _0411_ | _0412_;
  assign _0414_ = | 32'd0;
  assign _0415_ = 1'h0 | _0414_;
  assign _0416_ = xives[47:45] == { _0268_, _0385_, _0353_ };
  assign _0417_ = int_level_l[0] & _0416_;
  assign _0418_ = _0417_ ? 1'h1 : 1'h0;
  assign _0419_ = xives[44:42] == { _0268_, _0385_, _0353_ };
  assign _0420_ = int_level_l[1] & _0419_;
  assign _0421_ = _0420_ ? 1'h1 : 1'h0;
  assign _0422_ = xives[41:39] == { _0268_, _0385_, _0353_ };
  assign _0423_ = int_level_l[2] & _0422_;
  assign _0424_ = _0423_ ? 1'h1 : 1'h0;
  assign _0425_ = xives[38:36] == { _0268_, _0385_, _0353_ };
  assign _0426_ = int_level_l[3] & _0425_;
  assign _0427_ = _0426_ ? 1'h1 : 1'h0;
  assign _0428_ = xives[35:33] == { _0268_, _0385_, _0353_ };
  assign _0429_ = int_level_l[4] & _0428_;
  assign _0430_ = _0429_ ? 1'h1 : 1'h0;
  assign _0431_ = xives[32:30] == { _0268_, _0385_, _0353_ };
  assign _0432_ = int_level_l[5] & _0431_;
  assign _0433_ = _0432_ ? 1'h1 : 1'h0;
  assign _0434_ = xives[29:27] == { _0268_, _0385_, _0353_ };
  assign _0435_ = int_level_l[6] & _0434_;
  assign _0436_ = _0435_ ? 1'h1 : 1'h0;
  assign _0437_ = xives[26:24] == { _0268_, _0385_, _0353_ };
  assign _0438_ = int_level_l[7] & _0437_;
  assign _0439_ = _0438_ ? 1'h1 : 1'h0;
  assign _0440_ = xives[23:21] == { _0268_, _0385_, _0353_ };
  assign _0441_ = int_level_l[8] & _0440_;
  assign _0442_ = _0441_ ? 1'h1 : 1'h0;
  assign _0443_ = xives[20:18] == { _0268_, _0385_, _0353_ };
  assign _0444_ = int_level_l[9] & _0443_;
  assign _0445_ = _0444_ ? 1'h1 : 1'h0;
  assign _0446_ = xives[17:15] == { _0268_, _0385_, _0353_ };
  assign _0447_ = int_level_l[10] & _0446_;
  assign _0448_ = _0447_ ? 1'h1 : 1'h0;
  assign _0449_ = xives[14:12] == { _0268_, _0385_, _0353_ };
  assign _0450_ = int_level_l[11] & _0449_;
  assign _0451_ = _0450_ ? 1'h1 : 1'h0;
  assign _0452_ = xives[11:9] == { _0268_, _0385_, _0353_ };
  assign _0453_ = int_level_l[12] & _0452_;
  assign _0454_ = _0453_ ? 1'h1 : 1'h0;
  assign _0455_ = xives[8:6] == { _0268_, _0385_, _0353_ };
  assign _0456_ = int_level_l[13] & _0455_;
  assign _0457_ = _0456_ ? 1'h1 : 1'h0;
  assign _0458_ = xives[5:3] == { _0268_, _0385_, _0353_ };
  assign _0459_ = int_level_l[14] & _0458_;
  assign _0460_ = _0459_ ? 1'h1 : 1'h0;
  assign _0461_ = xives[2:0] == { _0268_, _0385_, _0353_ };
  assign _0462_ = int_level_l[15] & _0461_;
  assign _0463_ = _0462_ ? 1'h1 : 1'h0;
  assign _0464_ = - $signed({ 1'h1, _0460_, _0457_, _0454_, _0451_, _0448_, _0445_, _0442_, _0439_, _0436_, _0433_, _0430_, _0427_, _0424_, _0421_, _0418_ });
  assign _0465_ = _0464_ & { 1'h1, _0460_, _0457_, _0454_, _0451_, _0448_, _0445_, _0442_, _0439_, _0436_, _0433_, _0430_, _0427_, _0424_, _0421_, _0418_ };
  assign _0466_ = _0464_ | { 1'h1, _0460_, _0457_, _0454_, _0451_, _0448_, _0445_, _0442_, _0439_, _0436_, _0433_, _0430_, _0427_, _0424_, _0421_, _0418_ };
  assign _0467_ = ~ _0466_[0];
  assign _0468_ = _0466_[1] & _0467_;
  assign _0469_ = 1'h0 | _0468_;
  assign _0470_ = ~ _0466_[2];
  assign _0471_ = _0466_[3] & _0470_;
  assign _0472_ = _0469_ | _0471_;
  assign _0473_ = ~ _0466_[4];
  assign _0474_ = _0466_[5] & _0473_;
  assign _0475_ = _0472_ | _0474_;
  assign _0476_ = ~ _0466_[6];
  assign _0477_ = _0466_[7] & _0476_;
  assign _0478_ = _0475_ | _0477_;
  assign _0479_ = ~ _0466_[8];
  assign _0480_ = _0466_[9] & _0479_;
  assign _0481_ = _0478_ | _0480_;
  assign _0482_ = ~ _0466_[10];
  assign _0483_ = _0466_[11] & _0482_;
  assign _0484_ = _0481_ | _0483_;
  assign _0485_ = ~ _0466_[12];
  assign _0486_ = _0466_[13] & _0485_;
  assign _0487_ = _0484_ | _0486_;
  assign _0488_ = ~ _0466_[14];
  assign _0489_ = _0466_[15] & _0488_;
  assign _0490_ = _0487_ | _0489_;
  assign _0491_ = ~ _0466_[15];
  assign _0492_ = _0466_[15] & _0491_;
  assign _0493_ = _0490_ | _0492_;
  assign _0494_ = ~ _0466_[15];
  assign _0495_ = _0466_[15] & _0494_;
  assign _0496_ = _0493_ | _0495_;
  assign _0497_ = ~ _0466_[15];
  assign _0498_ = _0466_[15] & _0497_;
  assign _0499_ = _0496_ | _0498_;
  assign _0500_ = ~ _0466_[15];
  assign _0501_ = _0466_[15] & _0500_;
  assign _0502_ = _0499_ | _0501_;
  assign _0503_ = ~ _0466_[15];
  assign _0504_ = _0466_[15] & _0503_;
  assign _0505_ = _0502_ | _0504_;
  assign _0506_ = ~ _0466_[15];
  assign _0507_ = _0466_[15] & _0506_;
  assign _0508_ = _0505_ | _0507_;
  assign _0509_ = ~ _0466_[15];
  assign _0510_ = _0466_[15] & _0509_;
  assign _0511_ = _0508_ | _0510_;
  assign _0512_ = ~ _0466_[15];
  assign _0513_ = _0466_[15] & _0512_;
  assign _0514_ = _0511_ | _0513_;
  assign _0515_ = ~ _0466_[15];
  assign _0516_ = _0466_[15] & _0515_;
  assign _0517_ = _0514_ | _0516_;
  assign _0518_ = ~ _0466_[15];
  assign _0519_ = _0466_[15] & _0518_;
  assign _0520_ = _0517_ | _0519_;
  assign _0521_ = ~ _0466_[15];
  assign _0522_ = _0466_[15] & _0521_;
  assign _0523_ = _0520_ | _0522_;
  assign _0524_ = ~ _0466_[15];
  assign _0525_ = _0466_[15] & _0524_;
  assign _0526_ = _0523_ | _0525_;
  assign _0527_ = ~ _0466_[15];
  assign _0528_ = _0466_[15] & _0527_;
  assign _0529_ = _0526_ | _0528_;
  assign _0530_ = ~ _0466_[15];
  assign _0531_ = _0466_[15] & _0530_;
  assign _0532_ = _0529_ | _0531_;
  assign _0533_ = ~ _0466_[15];
  assign _0534_ = _0466_[15] & _0533_;
  assign _0535_ = _0532_ | _0534_;
  assign _0536_ = ~ _0466_[15];
  assign _0537_ = _0466_[15] & _0536_;
  assign _0538_ = _0535_ | _0537_;
  assign _0539_ = ~ _0466_[15];
  assign _0540_ = _0466_[15] & _0539_;
  assign _0541_ = _0538_ | _0540_;
  assign _0542_ = ~ _0466_[15];
  assign _0543_ = _0466_[15] & _0542_;
  assign _0544_ = _0541_ | _0543_;
  assign _0545_ = ~ _0466_[15];
  assign _0546_ = _0466_[15] & _0545_;
  assign _0547_ = _0544_ | _0546_;
  assign _0548_ = ~ _0466_[15];
  assign _0549_ = _0466_[15] & _0548_;
  assign _0550_ = _0547_ | _0549_;
  assign _0551_ = ~ _0466_[15];
  assign _0552_ = _0466_[15] & _0551_;
  assign _0553_ = _0550_ | _0552_;
  assign _0554_ = ~ _0466_[15];
  assign _0555_ = _0466_[15] & _0554_;
  assign _0556_ = _0553_ | _0555_;
  assign _0557_ = ~ _0466_[15];
  assign _0558_ = _0466_[15] & _0557_;
  assign _0559_ = _0556_ | _0558_;
  assign _0560_ = ~ _0466_[15];
  assign _0561_ = _0466_[15] & _0560_;
  assign _0562_ = _0559_ | _0561_;
  assign _0563_ = ~ _0466_[1];
  assign _0564_ = _0466_[3] & _0563_;
  assign _0565_ = 1'h0 | _0564_;
  assign _0566_ = ~ _0466_[5];
  assign _0567_ = _0466_[7] & _0566_;
  assign _0568_ = _0565_ | _0567_;
  assign _0569_ = ~ _0466_[9];
  assign _0570_ = _0466_[11] & _0569_;
  assign _0571_ = _0568_ | _0570_;
  assign _0572_ = ~ _0466_[13];
  assign _0573_ = _0466_[15] & _0572_;
  assign _0574_ = _0571_ | _0573_;
  assign _0575_ = ~ _0466_[15];
  assign _0576_ = _0466_[15] & _0575_;
  assign _0577_ = _0574_ | _0576_;
  assign _0578_ = ~ _0466_[15];
  assign _0579_ = _0466_[15] & _0578_;
  assign _0580_ = _0577_ | _0579_;
  assign _0581_ = ~ _0466_[15];
  assign _0582_ = _0466_[15] & _0581_;
  assign _0583_ = _0580_ | _0582_;
  assign _0584_ = ~ _0466_[15];
  assign _0585_ = _0466_[15] & _0584_;
  assign _0586_ = _0583_ | _0585_;
  assign _0587_ = ~ _0466_[15];
  assign _0588_ = _0466_[15] & _0587_;
  assign _0589_ = _0586_ | _0588_;
  assign _0590_ = ~ _0466_[15];
  assign _0591_ = _0466_[15] & _0590_;
  assign _0592_ = _0589_ | _0591_;
  assign _0593_ = ~ _0466_[15];
  assign _0594_ = _0466_[15] & _0593_;
  assign _0595_ = _0592_ | _0594_;
  assign _0596_ = ~ _0466_[15];
  assign _0597_ = _0466_[15] & _0596_;
  assign _0598_ = _0595_ | _0597_;
  assign _0599_ = ~ _0466_[15];
  assign _0600_ = _0466_[15] & _0599_;
  assign _0601_ = _0598_ | _0600_;
  assign _0602_ = ~ _0466_[15];
  assign _0603_ = _0466_[15] & _0602_;
  assign _0604_ = _0601_ | _0603_;
  assign _0605_ = ~ _0466_[15];
  assign _0606_ = _0466_[15] & _0605_;
  assign _0607_ = _0604_ | _0606_;
  assign _0608_ = ~ _0466_[15];
  assign _0609_ = _0466_[15] & _0608_;
  assign _0610_ = _0607_ | _0609_;
  assign _0611_ = ~ _0466_[3];
  assign _0612_ = _0466_[7] & _0611_;
  assign _0613_ = 1'h0 | _0612_;
  assign _0614_ = ~ _0466_[11];
  assign _0615_ = _0466_[15] & _0614_;
  assign _0616_ = _0613_ | _0615_;
  assign _0617_ = ~ _0466_[15];
  assign _0618_ = _0466_[15] & _0617_;
  assign _0619_ = _0616_ | _0618_;
  assign _0620_ = ~ _0466_[15];
  assign _0621_ = _0466_[15] & _0620_;
  assign _0622_ = _0619_ | _0621_;
  assign _0623_ = ~ _0466_[15];
  assign _0624_ = _0466_[15] & _0623_;
  assign _0625_ = _0622_ | _0624_;
  assign _0626_ = ~ _0466_[15];
  assign _0627_ = _0466_[15] & _0626_;
  assign _0628_ = _0625_ | _0627_;
  assign _0629_ = ~ _0466_[15];
  assign _0630_ = _0466_[15] & _0629_;
  assign _0631_ = _0628_ | _0630_;
  assign _0632_ = ~ _0466_[15];
  assign _0633_ = _0466_[15] & _0632_;
  assign _0634_ = _0631_ | _0633_;
  assign _0635_ = ~ _0466_[7];
  assign _0636_ = _0466_[15] & _0635_;
  assign _0637_ = 1'h0 | _0636_;
  assign _0638_ = ~ _0466_[15];
  assign _0639_ = _0466_[15] & _0638_;
  assign _0640_ = _0637_ | _0639_;
  assign _0641_ = ~ _0466_[15];
  assign _0642_ = _0466_[15] & _0641_;
  assign _0643_ = _0640_ | _0642_;
  assign _0644_ = ~ _0466_[15];
  assign _0645_ = _0466_[15] & _0644_;
  assign _0646_ = _0643_ | _0645_;
  assign _0647_ = ~ _0466_[15];
  assign _0648_ = _0466_[15] & _0647_;
  assign _0649_ = 1'h0 | _0648_;
  assign _0650_ = ~ _0466_[15];
  assign _0651_ = _0466_[15] & _0650_;
  assign _0652_ = _0649_ | _0651_;
  assign _0653_ = ~ _0466_[15];
  assign _0654_ = _0466_[15] & _0653_;
  assign _0655_ = 1'h0 | _0654_;
  assign _0656_ = | _0465_[1];
  assign _0657_ = 1'h0 | _0656_;
  assign _0658_ = | _0465_[3];
  assign _0659_ = _0657_ | _0658_;
  assign _0660_ = | _0465_[5];
  assign _0661_ = _0659_ | _0660_;
  assign _0662_ = | _0465_[7];
  assign _0663_ = _0661_ | _0662_;
  assign _0664_ = | _0465_[9];
  assign _0665_ = _0663_ | _0664_;
  assign _0666_ = | _0465_[11];
  assign _0667_ = _0665_ | _0666_;
  assign _0668_ = | _0465_[13];
  assign _0669_ = _0667_ | _0668_;
  assign _0670_ = | _0465_[15];
  assign _0671_ = _0669_ | _0670_;
  assign _0672_ = | 1'h0;
  assign _0673_ = _0671_ | _0672_;
  assign _0674_ = | 1'h0;
  assign _0675_ = _0673_ | _0674_;
  assign _0676_ = | 1'h0;
  assign _0677_ = _0675_ | _0676_;
  assign _0678_ = | 1'h0;
  assign _0679_ = _0677_ | _0678_;
  assign _0680_ = | 1'h0;
  assign _0681_ = _0679_ | _0680_;
  assign _0682_ = | 1'h0;
  assign _0683_ = _0681_ | _0682_;
  assign _0684_ = | 1'h0;
  assign _0685_ = _0683_ | _0684_;
  assign _0686_ = | 1'h0;
  assign _0687_ = _0685_ | _0686_;
  assign _0688_ = | 1'h0;
  assign _0689_ = _0687_ | _0688_;
  assign _0690_ = | 1'h0;
  assign _0691_ = _0689_ | _0690_;
  assign _0692_ = | 1'h0;
  assign _0693_ = _0691_ | _0692_;
  assign _0694_ = | 1'h0;
  assign _0695_ = _0693_ | _0694_;
  assign _0696_ = | 1'h0;
  assign _0697_ = _0695_ | _0696_;
  assign _0698_ = | 1'h0;
  assign _0699_ = _0697_ | _0698_;
  assign _0700_ = | 1'h0;
  assign _0701_ = _0699_ | _0700_;
  assign _0702_ = | 1'h0;
  assign _0703_ = _0701_ | _0702_;
  assign _0704_ = | 1'h0;
  assign _0705_ = _0703_ | _0704_;
  assign _0706_ = | 1'h0;
  assign _0707_ = _0705_ | _0706_;
  assign _0708_ = | 1'h0;
  assign _0709_ = _0707_ | _0708_;
  assign _0710_ = | 1'h0;
  assign _0711_ = _0709_ | _0710_;
  assign _0712_ = | 1'h0;
  assign _0713_ = _0711_ | _0712_;
  assign _0714_ = | 1'h0;
  assign _0715_ = _0713_ | _0714_;
  assign _0716_ = | 1'h0;
  assign _0717_ = _0715_ | _0716_;
  assign _0718_ = | 1'h0;
  assign _0719_ = _0717_ | _0718_;
  assign _0720_ = | _0465_[3:2];
  assign _0721_ = 1'h0 | _0720_;
  assign _0722_ = | _0465_[7:6];
  assign _0723_ = _0721_ | _0722_;
  assign _0724_ = | _0465_[11:10];
  assign _0725_ = _0723_ | _0724_;
  assign _0726_ = | _0465_[15:14];
  assign _0727_ = _0725_ | _0726_;
  assign _0728_ = | 2'h0;
  assign _0729_ = _0727_ | _0728_;
  assign _0730_ = | 2'h0;
  assign _0731_ = _0729_ | _0730_;
  assign _0732_ = | 2'h0;
  assign _0733_ = _0731_ | _0732_;
  assign _0734_ = | 2'h0;
  assign _0735_ = _0733_ | _0734_;
  assign _0736_ = | 2'h0;
  assign _0737_ = _0735_ | _0736_;
  assign _0738_ = | 2'h0;
  assign _0739_ = _0737_ | _0738_;
  assign _0740_ = | 2'h0;
  assign _0741_ = _0739_ | _0740_;
  assign _0742_ = | 2'h0;
  assign _0743_ = _0741_ | _0742_;
  assign _0744_ = | 2'h0;
  assign _0745_ = _0743_ | _0744_;
  assign _0746_ = | 2'h0;
  assign _0747_ = _0745_ | _0746_;
  assign _0748_ = | 2'h0;
  assign _0749_ = _0747_ | _0748_;
  assign _0750_ = | 2'h0;
  assign _0751_ = _0749_ | _0750_;
  assign _0752_ = | _0465_[7:4];
  assign _0753_ = 1'h0 | _0752_;
  assign _0754_ = | _0465_[15:12];
  assign _0755_ = _0753_ | _0754_;
  assign _0756_ = | 4'h0;
  assign _0757_ = _0755_ | _0756_;
  assign _0758_ = | 4'h0;
  assign _0759_ = _0757_ | _0758_;
  assign _0760_ = | 4'h0;
  assign _0761_ = _0759_ | _0760_;
  assign _0762_ = | 4'h0;
  assign _0763_ = _0761_ | _0762_;
  assign _0764_ = | 4'h0;
  assign _0765_ = _0763_ | _0764_;
  assign _0766_ = | 4'h0;
  assign _0767_ = _0765_ | _0766_;
  assign _0768_ = | _0465_[15:8];
  assign _0769_ = 1'h0 | _0768_;
  assign _0770_ = | 8'h00;
  assign _0771_ = _0769_ | _0770_;
  assign _0772_ = | 8'h00;
  assign _0773_ = _0771_ | _0772_;
  assign _0774_ = | 8'h00;
  assign _0775_ = _0773_ | _0774_;
  assign _0776_ = | 16'h0000;
  assign _0777_ = 1'h0 | _0776_;
  assign _0778_ = | 16'h0000;
  assign _0779_ = _0777_ | _0778_;
  assign _0780_ = | 32'd0;
  assign _0781_ = 1'h0 | _0780_;
  assign _0782_ = { _0268_, _0385_, _0353_ } == 3'h7;
  assign _0783_ = _0782_ ? 8'hff : { 5'h00, _0268_, _0385_, _0353_ };
  assign _0799_ = ~ _0044_[3];
  assign _0800_ = ~ _0044_[2];
  assign _0801_ = _0799_ & _0800_;
  assign _0802_ = _0799_ & _0044_[2];
  assign _0803_ = _0044_[3] & _0800_;
  assign _0804_ = _0044_[3] & _0044_[2];
  assign _0805_ = ~ _0044_[1];
  assign _0806_ = _0801_ & _0805_;
  assign _0807_ = _0801_ & _0044_[1];
  assign _0808_ = _0802_ & _0805_;
  assign _0809_ = _0802_ & _0044_[1];
  assign _0810_ = _0803_ & _0805_;
  assign _0811_ = _0803_ & _0044_[1];
  assign _0812_ = _0804_ & _0805_;
  assign _0813_ = _0804_ & _0044_[1];
  assign _0814_ = ~ _0044_[0];
  assign _0815_ = _0806_ & _0814_;
  assign _0816_ = _0806_ & _0044_[0];
  assign _0817_ = _0807_ & _0814_;
  assign _0818_ = _0807_ & _0044_[0];
  assign _0819_ = _0808_ & _0814_;
  assign _0820_ = _0808_ & _0044_[0];
  assign _0821_ = _0809_ & _0814_;
  assign _0822_ = _0809_ & _0044_[0];
  assign _0823_ = _0810_ & _0814_;
  assign _0824_ = _0810_ & _0044_[0];
  assign _0825_ = _0811_ & _0814_;
  assign _0826_ = _0811_ & _0044_[0];
  assign _0827_ = _0812_ & _0814_;
  assign _0828_ = _0812_ & _0044_[0];
  assign _0829_ = _0813_ & _0814_;
  assign _0830_ = _0813_ & _0044_[0];
  assign _0831_ = _0815_ & reg_is_xive;
  assign _0832_ = _0831_ ? _0046_ : xives[2:0];
  assign _0833_ = _0816_ & reg_is_xive;
  assign _0834_ = _0833_ ? _0046_ : xives[5:3];
  assign _0835_ = _0817_ & reg_is_xive;
  assign _0836_ = _0835_ ? _0046_ : xives[8:6];
  assign _0837_ = _0818_ & reg_is_xive;
  assign _0838_ = _0837_ ? _0046_ : xives[11:9];
  assign _0839_ = _0819_ & reg_is_xive;
  assign _0840_ = _0839_ ? _0046_ : xives[14:12];
  assign _0841_ = _0820_ & reg_is_xive;
  assign _0842_ = _0841_ ? _0046_ : xives[17:15];
  assign _0843_ = _0821_ & reg_is_xive;
  assign _0844_ = _0843_ ? _0046_ : xives[20:18];
  assign _0845_ = _0822_ & reg_is_xive;
  assign _0846_ = _0845_ ? _0046_ : xives[23:21];
  assign _0847_ = _0823_ & reg_is_xive;
  assign _0848_ = _0847_ ? _0046_ : xives[26:24];
  assign _0849_ = _0824_ & reg_is_xive;
  assign _0850_ = _0849_ ? _0046_ : xives[29:27];
  assign _0851_ = _0825_ & reg_is_xive;
  assign _0852_ = _0851_ ? _0046_ : xives[32:30];
  assign _0853_ = _0826_ & reg_is_xive;
  assign _0854_ = _0853_ ? _0046_ : xives[35:33];
  assign _0855_ = _0827_ & reg_is_xive;
  assign _0856_ = _0855_ ? _0046_ : xives[38:36];
  assign _0857_ = _0828_ & reg_is_xive;
  assign _0858_ = _0857_ ? _0046_ : xives[41:39];
  assign _0859_ = _0829_ & reg_is_xive;
  assign _0860_ = _0859_ ? _0046_ : xives[44:42];
  assign _0861_ = _0830_ & reg_is_xive;
  assign _0862_ = _0861_ ? _0046_ : xives[47:45];
  assign _0863_ = ~ xives[47];
  assign _0864_ = ~ xives[46];
  assign _0865_ = _0863_ & _0864_;
  assign _0866_ = _0863_ & xives[46];
  assign _0867_ = xives[47] & _0864_;
  assign _0868_ = xives[47] & xives[46];
  assign _0869_ = ~ xives[45];
  assign _0870_ = _0865_ & _0869_;
  assign _0871_ = _0865_ & xives[45];
  assign _0872_ = _0866_ & _0869_;
  assign _0873_ = _0866_ & xives[45];
  assign _0874_ = _0867_ & _0869_;
  assign _0875_ = _0867_ & xives[45];
  assign _0876_ = _0868_ & _0869_;
  assign _0877_ = _0868_ & xives[45];
  assign _0878_ = _0870_ ? 1'h1 : 1'h0;
  assign _0879_ = _0871_ ? 1'h1 : 1'h0;
  assign _0880_ = _0872_ ? 1'h1 : 1'h0;
  assign _0881_ = _0873_ ? 1'h1 : 1'h0;
  assign _0882_ = _0874_ ? 1'h1 : 1'h0;
  assign _0883_ = _0875_ ? 1'h1 : 1'h0;
  assign _0884_ = _0876_ ? 1'h1 : 1'h0;
  assign _0885_ = _0877_ ? 1'h1 : 1'h0;
  assign _0886_ = ~ xives[44];
  assign _0887_ = ~ xives[43];
  assign _0888_ = _0886_ & _0887_;
  assign _0889_ = _0886_ & xives[43];
  assign _0890_ = xives[44] & _0887_;
  assign _0891_ = xives[44] & xives[43];
  assign _0892_ = ~ xives[42];
  assign _0893_ = _0888_ & _0892_;
  assign _0894_ = _0888_ & xives[42];
  assign _0895_ = _0889_ & _0892_;
  assign _0896_ = _0889_ & xives[42];
  assign _0897_ = _0890_ & _0892_;
  assign _0898_ = _0890_ & xives[42];
  assign _0899_ = _0891_ & _0892_;
  assign _0900_ = _0891_ & xives[42];
  assign _0901_ = _0893_ ? 1'h1 : 1'h0;
  assign _0902_ = _0894_ ? 1'h1 : 1'h0;
  assign _0903_ = _0895_ ? 1'h1 : 1'h0;
  assign _0904_ = _0896_ ? 1'h1 : 1'h0;
  assign _0905_ = _0897_ ? 1'h1 : 1'h0;
  assign _0906_ = _0898_ ? 1'h1 : 1'h0;
  assign _0907_ = _0899_ ? 1'h1 : 1'h0;
  assign _0908_ = _0900_ ? 1'h1 : 1'h0;
  assign _0909_ = ~ xives[41];
  assign _0910_ = ~ xives[40];
  assign _0911_ = _0909_ & _0910_;
  assign _0912_ = _0909_ & xives[40];
  assign _0913_ = xives[41] & _0910_;
  assign _0914_ = xives[41] & xives[40];
  assign _0915_ = ~ xives[39];
  assign _0916_ = _0911_ & _0915_;
  assign _0917_ = _0911_ & xives[39];
  assign _0918_ = _0912_ & _0915_;
  assign _0919_ = _0912_ & xives[39];
  assign _0920_ = _0913_ & _0915_;
  assign _0921_ = _0913_ & xives[39];
  assign _0922_ = _0914_ & _0915_;
  assign _0923_ = _0914_ & xives[39];
  assign _0924_ = _0916_ ? 1'h1 : 1'h0;
  assign _0925_ = _0917_ ? 1'h1 : 1'h0;
  assign _0926_ = _0918_ ? 1'h1 : 1'h0;
  assign _0927_ = _0919_ ? 1'h1 : 1'h0;
  assign _0928_ = _0920_ ? 1'h1 : 1'h0;
  assign _0929_ = _0921_ ? 1'h1 : 1'h0;
  assign _0930_ = _0922_ ? 1'h1 : 1'h0;
  assign _0931_ = _0923_ ? 1'h1 : 1'h0;
  assign _0932_ = ~ xives[38];
  assign _0933_ = ~ xives[37];
  assign _0934_ = _0932_ & _0933_;
  assign _0935_ = _0932_ & xives[37];
  assign _0936_ = xives[38] & _0933_;
  assign _0937_ = xives[38] & xives[37];
  assign _0938_ = ~ xives[36];
  assign _0939_ = _0934_ & _0938_;
  assign _0940_ = _0934_ & xives[36];
  assign _0941_ = _0935_ & _0938_;
  assign _0942_ = _0935_ & xives[36];
  assign _0943_ = _0936_ & _0938_;
  assign _0944_ = _0936_ & xives[36];
  assign _0945_ = _0937_ & _0938_;
  assign _0946_ = _0937_ & xives[36];
  assign _0947_ = _0939_ ? 1'h1 : 1'h0;
  assign _0948_ = _0940_ ? 1'h1 : 1'h0;
  assign _0949_ = _0941_ ? 1'h1 : 1'h0;
  assign _0950_ = _0942_ ? 1'h1 : 1'h0;
  assign _0951_ = _0943_ ? 1'h1 : 1'h0;
  assign _0952_ = _0944_ ? 1'h1 : 1'h0;
  assign _0953_ = _0945_ ? 1'h1 : 1'h0;
  assign _0954_ = _0946_ ? 1'h1 : 1'h0;
  assign _0955_ = ~ xives[35];
  assign _0956_ = ~ xives[34];
  assign _0957_ = _0955_ & _0956_;
  assign _0958_ = _0955_ & xives[34];
  assign _0959_ = xives[35] & _0956_;
  assign _0960_ = xives[35] & xives[34];
  assign _0961_ = ~ xives[33];
  assign _0962_ = _0957_ & _0961_;
  assign _0963_ = _0957_ & xives[33];
  assign _0964_ = _0958_ & _0961_;
  assign _0965_ = _0958_ & xives[33];
  assign _0966_ = _0959_ & _0961_;
  assign _0967_ = _0959_ & xives[33];
  assign _0968_ = _0960_ & _0961_;
  assign _0969_ = _0960_ & xives[33];
  assign _0970_ = _0962_ ? 1'h1 : 1'h0;
  assign _0971_ = _0963_ ? 1'h1 : 1'h0;
  assign _0972_ = _0964_ ? 1'h1 : 1'h0;
  assign _0973_ = _0965_ ? 1'h1 : 1'h0;
  assign _0974_ = _0966_ ? 1'h1 : 1'h0;
  assign _0975_ = _0967_ ? 1'h1 : 1'h0;
  assign _0976_ = _0968_ ? 1'h1 : 1'h0;
  assign _0977_ = _0969_ ? 1'h1 : 1'h0;
  assign _0978_ = ~ xives[32];
  assign _0979_ = ~ xives[31];
  assign _0980_ = _0978_ & _0979_;
  assign _0981_ = _0978_ & xives[31];
  assign _0982_ = xives[32] & _0979_;
  assign _0983_ = xives[32] & xives[31];
  assign _0984_ = ~ xives[30];
  assign _0985_ = _0980_ & _0984_;
  assign _0986_ = _0980_ & xives[30];
  assign _0987_ = _0981_ & _0984_;
  assign _0988_ = _0981_ & xives[30];
  assign _0989_ = _0982_ & _0984_;
  assign _0990_ = _0982_ & xives[30];
  assign _0991_ = _0983_ & _0984_;
  assign _0992_ = _0983_ & xives[30];
  assign _0993_ = _0985_ ? 1'h1 : 1'h0;
  assign _0994_ = _0986_ ? 1'h1 : 1'h0;
  assign _0995_ = _0987_ ? 1'h1 : 1'h0;
  assign _0996_ = _0988_ ? 1'h1 : 1'h0;
  assign _0997_ = _0989_ ? 1'h1 : 1'h0;
  assign _0998_ = _0990_ ? 1'h1 : 1'h0;
  assign _0999_ = _0991_ ? 1'h1 : 1'h0;
  assign _1000_ = _0992_ ? 1'h1 : 1'h0;
  assign _1001_ = ~ xives[29];
  assign _1002_ = ~ xives[28];
  assign _1003_ = _1001_ & _1002_;
  assign _1004_ = _1001_ & xives[28];
  assign _1005_ = xives[29] & _1002_;
  assign _1006_ = xives[29] & xives[28];
  assign _1007_ = ~ xives[27];
  assign _1008_ = _1003_ & _1007_;
  assign _1009_ = _1003_ & xives[27];
  assign _1010_ = _1004_ & _1007_;
  assign _1011_ = _1004_ & xives[27];
  assign _1012_ = _1005_ & _1007_;
  assign _1013_ = _1005_ & xives[27];
  assign _1014_ = _1006_ & _1007_;
  assign _1015_ = _1006_ & xives[27];
  assign _1016_ = _1008_ ? 1'h1 : 1'h0;
  assign _1017_ = _1009_ ? 1'h1 : 1'h0;
  assign _1018_ = _1010_ ? 1'h1 : 1'h0;
  assign _1019_ = _1011_ ? 1'h1 : 1'h0;
  assign _1020_ = _1012_ ? 1'h1 : 1'h0;
  assign _1021_ = _1013_ ? 1'h1 : 1'h0;
  assign _1022_ = _1014_ ? 1'h1 : 1'h0;
  assign _1023_ = _1015_ ? 1'h1 : 1'h0;
  assign _1024_ = ~ xives[26];
  assign _1025_ = ~ xives[25];
  assign _1026_ = _1024_ & _1025_;
  assign _1027_ = _1024_ & xives[25];
  assign _1028_ = xives[26] & _1025_;
  assign _1029_ = xives[26] & xives[25];
  assign _1030_ = ~ xives[24];
  assign _1031_ = _1026_ & _1030_;
  assign _1032_ = _1026_ & xives[24];
  assign _1033_ = _1027_ & _1030_;
  assign _1034_ = _1027_ & xives[24];
  assign _1035_ = _1028_ & _1030_;
  assign _1036_ = _1028_ & xives[24];
  assign _1037_ = _1029_ & _1030_;
  assign _1038_ = _1029_ & xives[24];
  assign _1039_ = _1031_ ? 1'h1 : 1'h0;
  assign _1040_ = _1032_ ? 1'h1 : 1'h0;
  assign _1041_ = _1033_ ? 1'h1 : 1'h0;
  assign _1042_ = _1034_ ? 1'h1 : 1'h0;
  assign _1043_ = _1035_ ? 1'h1 : 1'h0;
  assign _1044_ = _1036_ ? 1'h1 : 1'h0;
  assign _1045_ = _1037_ ? 1'h1 : 1'h0;
  assign _1046_ = _1038_ ? 1'h1 : 1'h0;
  assign _1047_ = ~ xives[23];
  assign _1048_ = ~ xives[22];
  assign _1049_ = _1047_ & _1048_;
  assign _1050_ = _1047_ & xives[22];
  assign _1051_ = xives[23] & _1048_;
  assign _1052_ = xives[23] & xives[22];
  assign _1053_ = ~ xives[21];
  assign _1054_ = _1049_ & _1053_;
  assign _1055_ = _1049_ & xives[21];
  assign _1056_ = _1050_ & _1053_;
  assign _1057_ = _1050_ & xives[21];
  assign _1058_ = _1051_ & _1053_;
  assign _1059_ = _1051_ & xives[21];
  assign _1060_ = _1052_ & _1053_;
  assign _1061_ = _1052_ & xives[21];
  assign _1062_ = _1054_ ? 1'h1 : 1'h0;
  assign _1063_ = _1055_ ? 1'h1 : 1'h0;
  assign _1064_ = _1056_ ? 1'h1 : 1'h0;
  assign _1065_ = _1057_ ? 1'h1 : 1'h0;
  assign _1066_ = _1058_ ? 1'h1 : 1'h0;
  assign _1067_ = _1059_ ? 1'h1 : 1'h0;
  assign _1068_ = _1060_ ? 1'h1 : 1'h0;
  assign _1069_ = _1061_ ? 1'h1 : 1'h0;
  assign _1070_ = ~ xives[20];
  assign _1071_ = ~ xives[19];
  assign _1072_ = _1070_ & _1071_;
  assign _1073_ = _1070_ & xives[19];
  assign _1074_ = xives[20] & _1071_;
  assign _1075_ = xives[20] & xives[19];
  assign _1076_ = ~ xives[18];
  assign _1077_ = _1072_ & _1076_;
  assign _1078_ = _1072_ & xives[18];
  assign _1079_ = _1073_ & _1076_;
  assign _1080_ = _1073_ & xives[18];
  assign _1081_ = _1074_ & _1076_;
  assign _1082_ = _1074_ & xives[18];
  assign _1083_ = _1075_ & _1076_;
  assign _1084_ = _1075_ & xives[18];
  assign _1085_ = _1077_ ? 1'h1 : 1'h0;
  assign _1086_ = _1078_ ? 1'h1 : 1'h0;
  assign _1087_ = _1079_ ? 1'h1 : 1'h0;
  assign _1088_ = _1080_ ? 1'h1 : 1'h0;
  assign _1089_ = _1081_ ? 1'h1 : 1'h0;
  assign _1090_ = _1082_ ? 1'h1 : 1'h0;
  assign _1091_ = _1083_ ? 1'h1 : 1'h0;
  assign _1092_ = _1084_ ? 1'h1 : 1'h0;
  assign _1093_ = ~ xives[17];
  assign _1094_ = ~ xives[16];
  assign _1095_ = _1093_ & _1094_;
  assign _1096_ = _1093_ & xives[16];
  assign _1097_ = xives[17] & _1094_;
  assign _1098_ = xives[17] & xives[16];
  assign _1099_ = ~ xives[15];
  assign _1100_ = _1095_ & _1099_;
  assign _1101_ = _1095_ & xives[15];
  assign _1102_ = _1096_ & _1099_;
  assign _1103_ = _1096_ & xives[15];
  assign _1104_ = _1097_ & _1099_;
  assign _1105_ = _1097_ & xives[15];
  assign _1106_ = _1098_ & _1099_;
  assign _1107_ = _1098_ & xives[15];
  assign _1108_ = _1100_ ? 1'h1 : 1'h0;
  assign _1109_ = _1101_ ? 1'h1 : 1'h0;
  assign _1110_ = _1102_ ? 1'h1 : 1'h0;
  assign _1111_ = _1103_ ? 1'h1 : 1'h0;
  assign _1112_ = _1104_ ? 1'h1 : 1'h0;
  assign _1113_ = _1105_ ? 1'h1 : 1'h0;
  assign _1114_ = _1106_ ? 1'h1 : 1'h0;
  assign _1115_ = _1107_ ? 1'h1 : 1'h0;
  assign _1116_ = ~ xives[14];
  assign _1117_ = ~ xives[13];
  assign _1118_ = _1116_ & _1117_;
  assign _1119_ = _1116_ & xives[13];
  assign _1120_ = xives[14] & _1117_;
  assign _1121_ = xives[14] & xives[13];
  assign _1122_ = ~ xives[12];
  assign _1123_ = _1118_ & _1122_;
  assign _1124_ = _1118_ & xives[12];
  assign _1125_ = _1119_ & _1122_;
  assign _1126_ = _1119_ & xives[12];
  assign _1127_ = _1120_ & _1122_;
  assign _1128_ = _1120_ & xives[12];
  assign _1129_ = _1121_ & _1122_;
  assign _1130_ = _1121_ & xives[12];
  assign _1131_ = _1123_ ? 1'h1 : 1'h0;
  assign _1132_ = _1124_ ? 1'h1 : 1'h0;
  assign _1133_ = _1125_ ? 1'h1 : 1'h0;
  assign _1134_ = _1126_ ? 1'h1 : 1'h0;
  assign _1135_ = _1127_ ? 1'h1 : 1'h0;
  assign _1136_ = _1128_ ? 1'h1 : 1'h0;
  assign _1137_ = _1129_ ? 1'h1 : 1'h0;
  assign _1138_ = _1130_ ? 1'h1 : 1'h0;
  assign _1139_ = ~ xives[11];
  assign _1140_ = ~ xives[10];
  assign _1141_ = _1139_ & _1140_;
  assign _1142_ = _1139_ & xives[10];
  assign _1143_ = xives[11] & _1140_;
  assign _1144_ = xives[11] & xives[10];
  assign _1145_ = ~ xives[9];
  assign _1146_ = _1141_ & _1145_;
  assign _1147_ = _1141_ & xives[9];
  assign _1148_ = _1142_ & _1145_;
  assign _1149_ = _1142_ & xives[9];
  assign _1150_ = _1143_ & _1145_;
  assign _1151_ = _1143_ & xives[9];
  assign _1152_ = _1144_ & _1145_;
  assign _1153_ = _1144_ & xives[9];
  assign _1154_ = _1146_ ? 1'h1 : 1'h0;
  assign _1155_ = _1147_ ? 1'h1 : 1'h0;
  assign _1156_ = _1148_ ? 1'h1 : 1'h0;
  assign _1157_ = _1149_ ? 1'h1 : 1'h0;
  assign _1158_ = _1150_ ? 1'h1 : 1'h0;
  assign _1159_ = _1151_ ? 1'h1 : 1'h0;
  assign _1160_ = _1152_ ? 1'h1 : 1'h0;
  assign _1161_ = _1153_ ? 1'h1 : 1'h0;
  assign _1162_ = ~ xives[8];
  assign _1163_ = ~ xives[7];
  assign _1164_ = _1162_ & _1163_;
  assign _1165_ = _1162_ & xives[7];
  assign _1166_ = xives[8] & _1163_;
  assign _1167_ = xives[8] & xives[7];
  assign _1168_ = ~ xives[6];
  assign _1169_ = _1164_ & _1168_;
  assign _1170_ = _1164_ & xives[6];
  assign _1171_ = _1165_ & _1168_;
  assign _1172_ = _1165_ & xives[6];
  assign _1173_ = _1166_ & _1168_;
  assign _1174_ = _1166_ & xives[6];
  assign _1175_ = _1167_ & _1168_;
  assign _1176_ = _1167_ & xives[6];
  assign _1177_ = _1169_ ? 1'h1 : 1'h0;
  assign _1178_ = _1170_ ? 1'h1 : 1'h0;
  assign _1179_ = _1171_ ? 1'h1 : 1'h0;
  assign _1180_ = _1172_ ? 1'h1 : 1'h0;
  assign _1181_ = _1173_ ? 1'h1 : 1'h0;
  assign _1182_ = _1174_ ? 1'h1 : 1'h0;
  assign _1183_ = _1175_ ? 1'h1 : 1'h0;
  assign _1184_ = _1176_ ? 1'h1 : 1'h0;
  assign _1185_ = ~ xives[5];
  assign _1186_ = ~ xives[4];
  assign _1187_ = _1185_ & _1186_;
  assign _1188_ = _1185_ & xives[4];
  assign _1189_ = xives[5] & _1186_;
  assign _1190_ = xives[5] & xives[4];
  assign _1191_ = ~ xives[3];
  assign _1192_ = _1187_ & _1191_;
  assign _1193_ = _1187_ & xives[3];
  assign _1194_ = _1188_ & _1191_;
  assign _1195_ = _1188_ & xives[3];
  assign _1196_ = _1189_ & _1191_;
  assign _1197_ = _1189_ & xives[3];
  assign _1198_ = _1190_ & _1191_;
  assign _1199_ = _1190_ & xives[3];
  assign _1200_ = _1192_ ? 1'h1 : 1'h0;
  assign _1201_ = _1193_ ? 1'h1 : 1'h0;
  assign _1202_ = _1194_ ? 1'h1 : 1'h0;
  assign _1203_ = _1195_ ? 1'h1 : 1'h0;
  assign _1204_ = _1196_ ? 1'h1 : 1'h0;
  assign _1205_ = _1197_ ? 1'h1 : 1'h0;
  assign _1206_ = _1198_ ? 1'h1 : 1'h0;
  assign _1207_ = _1199_ ? 1'h1 : 1'h0;
  assign _1208_ = ~ xives[2];
  assign _1209_ = ~ xives[1];
  assign _1210_ = _1208_ & _1209_;
  assign _1211_ = _1208_ & xives[1];
  assign _1212_ = xives[2] & _1209_;
  assign _1213_ = xives[2] & xives[1];
  assign _1214_ = ~ xives[0];
  assign _1215_ = _1210_ & _1214_;
  assign _1216_ = _1210_ & xives[0];
  assign _1217_ = _1211_ & _1214_;
  assign _1218_ = _1211_ & xives[0];
  assign _1219_ = _1212_ & _1214_;
  assign _1220_ = _1212_ & xives[0];
  assign _1221_ = _1213_ & _1214_;
  assign _1222_ = _1213_ & xives[0];
  assign _1223_ = _1215_ ? 1'h1 : 1'h0;
  assign _1224_ = _1216_ ? 1'h1 : 1'h0;
  assign _1225_ = _1217_ ? 1'h1 : 1'h0;
  assign _1226_ = _1218_ ? 1'h1 : 1'h0;
  assign _1227_ = _1219_ ? 1'h1 : 1'h0;
  assign _1228_ = _1220_ ? 1'h1 : 1'h0;
  assign _1229_ = _1221_ ? 1'h1 : 1'h0;
  assign _1230_ = _1222_ ? 1'h1 : 1'h0;
  assign xives = _0049_;
  assign wb_valid = _0035_;
  assign reg_idx = \wb_in.adr [3:0];
  assign icp_out_next = { _0783_, _0646_, _0634_, _0751_, _0719_ };
  assign int_level_l = _0034_;
  assign reg_is_xive = \wb_in.adr [9];
  assign reg_is_config = _0031_;
  assign reg_is_debug = _0033_;
  assign \wb_out.dat  = _0042_[31:0];
  assign \wb_out.ack  = _0042_[32];
  assign \wb_out.stall  = 1'h0;
  assign \icp_out.src  = _0050_[3:0];
  assign \icp_out.pri  = _0050_[11:4];
endmodule