module bsg_mux_width_p39_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [77:0] data_i;
  input [0:0] sel_i;
  output [38:0] data_o;
  wire [38:0] data_o;
  wire N0,N1;
  assign data_o[38] = (N1)? data_i[38] : 
                      (N0)? data_i[77] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[37] = (N1)? data_i[37] : 
                      (N0)? data_i[76] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] : 
                      (N0)? data_i[75] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] : 
                      (N0)? data_i[74] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] : 
                      (N0)? data_i[73] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] : 
                      (N0)? data_i[72] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] : 
                      (N0)? data_i[71] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[70] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[69] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[68] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[67] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[66] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[65] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[64] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[63] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[62] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[61] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[60] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[59] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[58] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[57] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[56] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[55] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[54] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[53] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[52] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[51] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[50] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[49] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[48] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[47] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[46] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[45] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[44] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[43] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[42] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[41] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[40] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[39] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule