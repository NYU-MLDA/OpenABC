module AMOALU
(
  io_addr,
  io_cmd,
  io_typ,
  io_lhs,
  io_rhs,
  io_out
);

  input [5:0] io_addr;
  input [4:0] io_cmd;
  input [2:0] io_typ;
  input [63:0] io_lhs;
  input [63:0] io_rhs;
  output [63:0] io_out;
  wire [63:0] io_out,T49,T1,T2,out,adder_out,T50,T111,T51,T109,T52,T107,T53,T54,T116,T113,
  mask;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,wmask_63,wmask_48,wmask_47,wmask_40,
  wmask_39,wmask_32,wmask_31,wmask_24,wmask_23,wmask_16,wmask_15,wmask_8,wmask_7,
  wmask_0,N33,N34,T16,T28,T69,N35,T55_63_,T55_62_,T55_61_,T55_60_,T55_59_,T55_58_,
  T55_57_,T55_56_,T55_55_,T55_54_,T55_53_,T55_52_,T55_51_,T55_50_,T55_49_,T55_48_,
  T55_47_,T55_46_,T55_45_,T55_44_,T55_43_,T55_42_,T55_41_,T55_40_,T55_39_,T55_38_,
  T55_37_,T55_36_,T55_35_,T55_34_,T55_33_,T55_32_,T55_31_,T55_30_,T55_29_,T55_28_,
  T55_27_,T55_26_,T55_25_,T55_24_,T55_23_,T55_22_,T55_21_,T55_20_,T55_19_,T55_18_,
  T55_17_,T55_16_,less,N36,min,max,T106,N37,lt,T74,sgned,N38,cmp_lhs,cmp_rhs,T80,N39,
  word,T81,T84,T86,T91,N40,T92,N41,T104,T96,lt_hi,T97,eq_hi,lt_lo,N42,N43,N44,N45,
  N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,
  N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,
  N86,N87,N88,N89,N90;
  wire [56:55] wmask;
  wire [0:0] T119;
  wire [7:1] T8;
  wire [3:0] T10,T29;
  wire [1:1] T12,T21;
  wire [1:0] T23;
  wire [3:3] T27;
  wire [63:32] T56,rhs;
  assign T28 = { 1'b1, 1'b1 } <= io_typ[1:0];
  assign lt_lo = io_lhs[31:0] < io_rhs[31:0];
  assign eq_hi = io_lhs[63:32] == rhs;
  assign lt_hi = io_lhs[63:32] < rhs;
  assign N0 = cmp_lhs ^ cmp_rhs;
  assign T106 = ~N0;
  assign N42 = ~io_cmd[3];
  assign N43 = N42 | io_cmd[4];
  assign N44 = io_cmd[2] | N43;
  assign N45 = io_cmd[1] | N44;
  assign N46 = io_cmd[0] | N45;
  assign N47 = ~N46;
  assign N48 = ~io_cmd[1];
  assign N49 = ~io_cmd[0];
  assign N50 = N48 | N44;
  assign N51 = N49 | N50;
  assign N52 = ~N51;
  assign N53 = io_cmd[0] | N50;
  assign N54 = ~N53;
  assign N55 = ~io_addr[0];
  assign N56 = N49 | N45;
  assign N57 = ~N56;
  assign N58 = io_typ[0] | io_typ[1];
  assign N59 = ~N58;
  assign N60 = ~io_typ[0];
  assign N61 = N60 | io_typ[1];
  assign N62 = ~N61;
  assign N63 = ~io_cmd[2];
  assign N64 = N63 | N43;
  assign N65 = io_cmd[1] | N64;
  assign N66 = io_cmd[0] | N65;
  assign N67 = ~N66;
  assign N68 = N48 | N64;
  assign N69 = io_cmd[0] | N68;
  assign N70 = ~N69;
  assign N71 = N49 | N65;
  assign N72 = ~N71;
  assign N73 = N49 | N68;
  assign N74 = ~N73;
  assign N75 = ~io_typ[1];
  assign N76 = io_typ[0] | N75;
  assign N77 = ~N76;
  assign N78 = ~io_typ[2];
  assign N79 = io_typ[1] | N78;
  assign N80 = io_typ[0] | N79;
  assign N81 = ~N80;
  assign N82 = io_typ[1] | io_typ[2];
  assign N83 = io_typ[0] | N82;
  assign N84 = ~N83;
  assign N85 = N75 | io_typ[2];
  assign N86 = io_typ[0] | N85;
  assign N87 = ~N86;
  assign N88 = N75 | N78;
  assign N89 = io_typ[0] | N88;
  assign N90 = ~N89;
  assign adder_out = T116 + T113;
  assign { wmask_7, wmask_0 } = 1'b0 - T119[0];
  assign { wmask_15, wmask_8 } = 1'b0 - T8[1];
  assign { wmask_23, wmask_16 } = 1'b0 - T8[2];
  assign { wmask_31, wmask_24 } = 1'b0 - T8[3];
  assign { wmask_39, wmask_32 } = 1'b0 - T8[4];
  assign { wmask_47, wmask_40 } = 1'b0 - T8[5];
  assign { wmask[55:55], wmask_48 } = 1'b0 - T8[6];
  assign { wmask_63, wmask[56:56] } = 1'b0 - T8[7];
  assign { T8[3:1], T119[0:0] } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N2)? T10 : 1'b0;
  assign N1 = io_addr[2];
  assign N2 = N33;
  assign T10[1:0] = (N3)? { 1'b0, 1'b0 } : 
                    (N4)? { T12[1:1], N55 } : 1'b0;
  assign N3 = io_addr[1];
  assign N4 = N34;
  assign T23 = (N3)? { T12[1:1], N55 } : 
               (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign T29 = (N1)? T10 : 
               (N2)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign out = (N5)? adder_out : 
               (N6)? T50 : 1'b0;
  assign N5 = N47;
  assign N6 = N46;
  assign T50 = (N7)? T111 : 
               (N8)? T51 : 1'b0;
  assign N7 = N52;
  assign N8 = N51;
  assign T51 = (N9)? T109 : 
               (N10)? T52 : 1'b0;
  assign N9 = N54;
  assign N10 = N53;
  assign T52 = (N11)? T107 : 
               (N12)? T53 : 1'b0;
  assign N11 = N57;
  assign N12 = N56;
  assign T53 = (N13)? io_lhs : 
               (N14)? T54 : 1'b0;
  assign N13 = T69;
  assign N14 = N35;
  assign T54 = (N15)? { io_rhs[7:0], io_rhs[7:0], io_rhs[7:0], io_rhs[7:0], io_rhs[7:0], io_rhs[7:0], io_rhs[7:0], io_rhs[7:0] } : 
               (N16)? { T55_63_, T55_62_, T55_61_, T55_60_, T55_59_, T55_58_, T55_57_, T55_56_, T55_55_, T55_54_, T55_53_, T55_52_, T55_51_, T55_50_, T55_49_, T55_48_, T55_47_, T55_46_, T55_45_, T55_44_, T55_43_, T55_42_, T55_41_, T55_40_, T55_39_, T55_38_, T55_37_, T55_36_, T55_35_, T55_34_, T55_33_, T55_32_, T55_31_, T55_30_, T55_29_, T55_28_, T55_27_, T55_26_, T55_25_, T55_24_, T55_23_, T55_22_, T55_21_, T55_20_, T55_19_, T55_18_, T55_17_, T55_16_, io_rhs[15:0] } : 1'b0;
  assign N15 = N59;
  assign N16 = N58;
  assign { T55_63_, T55_62_, T55_61_, T55_60_, T55_59_, T55_58_, T55_57_, T55_56_, T55_55_, T55_54_, T55_53_, T55_52_, T55_51_, T55_50_, T55_49_, T55_48_, T55_47_, T55_46_, T55_45_, T55_44_, T55_43_, T55_42_, T55_41_, T55_40_, T55_39_, T55_38_, T55_37_, T55_36_, T55_35_, T55_34_, T55_33_, T55_32_, T55_31_, T55_30_, T55_29_, T55_28_, T55_27_, T55_26_, T55_25_, T55_24_, T55_23_, T55_22_, T55_21_, T55_20_, T55_19_, T55_18_, T55_17_, T55_16_ } = (N17)? { io_rhs[15:0], io_rhs[15:0], io_rhs[15:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N18)? { T56, io_rhs[31:16] } : 1'b0;
  assign N17 = N62;
  assign N18 = N61;
  assign T56 = (N19)? io_rhs[31:0] : 
               (N20)? io_rhs[63:32] : 1'b0;
  assign N19 = N77;
  assign N20 = N76;
  assign T69 = (N21)? min : 
               (N22)? max : 1'b0;
  assign N21 = less;
  assign N22 = N36;
  assign less = (N23)? lt : 
                (N24)? T74 : 1'b0;
  assign N23 = T106;
  assign N24 = N37;
  assign T74 = (N25)? cmp_lhs : 
               (N26)? cmp_rhs : 1'b0;
  assign N25 = sgned;
  assign N26 = N38;
  assign cmp_rhs = (N27)? io_rhs[31] : 
                   (N28)? rhs[63] : 1'b0;
  assign N27 = T80;
  assign N28 = N39;
  assign rhs = (N19)? io_rhs[31:0] : 
               (N20)? io_rhs[63:32] : 1'b0;
  assign cmp_lhs = (N29)? io_lhs[31] : 
                   (N30)? io_lhs[63] : 1'b0;
  assign N29 = T91;
  assign N30 = N40;
  assign lt = (N31)? T104 : 
              (N32)? T96 : 1'b0;
  assign N31 = word;
  assign N32 = N41;
  assign T104 = (N1)? lt_hi : 
                (N2)? lt_lo : 1'b0;
  assign io_out[63] = T49[63] | T1[63];
  assign io_out[62] = T49[62] | T1[62];
  assign io_out[61] = T49[61] | T1[61];
  assign io_out[60] = T49[60] | T1[60];
  assign io_out[59] = T49[59] | T1[59];
  assign io_out[58] = T49[58] | T1[58];
  assign io_out[57] = T49[57] | T1[57];
  assign io_out[56] = T49[56] | T1[56];
  assign io_out[55] = T49[55] | T1[55];
  assign io_out[54] = T49[54] | T1[54];
  assign io_out[53] = T49[53] | T1[53];
  assign io_out[52] = T49[52] | T1[52];
  assign io_out[51] = T49[51] | T1[51];
  assign io_out[50] = T49[50] | T1[50];
  assign io_out[49] = T49[49] | T1[49];
  assign io_out[48] = T49[48] | T1[48];
  assign io_out[47] = T49[47] | T1[47];
  assign io_out[46] = T49[46] | T1[46];
  assign io_out[45] = T49[45] | T1[45];
  assign io_out[44] = T49[44] | T1[44];
  assign io_out[43] = T49[43] | T1[43];
  assign io_out[42] = T49[42] | T1[42];
  assign io_out[41] = T49[41] | T1[41];
  assign io_out[40] = T49[40] | T1[40];
  assign io_out[39] = T49[39] | T1[39];
  assign io_out[38] = T49[38] | T1[38];
  assign io_out[37] = T49[37] | T1[37];
  assign io_out[36] = T49[36] | T1[36];
  assign io_out[35] = T49[35] | T1[35];
  assign io_out[34] = T49[34] | T1[34];
  assign io_out[33] = T49[33] | T1[33];
  assign io_out[32] = T49[32] | T1[32];
  assign io_out[31] = T49[31] | T1[31];
  assign io_out[30] = T49[30] | T1[30];
  assign io_out[29] = T49[29] | T1[29];
  assign io_out[28] = T49[28] | T1[28];
  assign io_out[27] = T49[27] | T1[27];
  assign io_out[26] = T49[26] | T1[26];
  assign io_out[25] = T49[25] | T1[25];
  assign io_out[24] = T49[24] | T1[24];
  assign io_out[23] = T49[23] | T1[23];
  assign io_out[22] = T49[22] | T1[22];
  assign io_out[21] = T49[21] | T1[21];
  assign io_out[20] = T49[20] | T1[20];
  assign io_out[19] = T49[19] | T1[19];
  assign io_out[18] = T49[18] | T1[18];
  assign io_out[17] = T49[17] | T1[17];
  assign io_out[16] = T49[16] | T1[16];
  assign io_out[15] = T49[15] | T1[15];
  assign io_out[14] = T49[14] | T1[14];
  assign io_out[13] = T49[13] | T1[13];
  assign io_out[12] = T49[12] | T1[12];
  assign io_out[11] = T49[11] | T1[11];
  assign io_out[10] = T49[10] | T1[10];
  assign io_out[9] = T49[9] | T1[9];
  assign io_out[8] = T49[8] | T1[8];
  assign io_out[7] = T49[7] | T1[7];
  assign io_out[6] = T49[6] | T1[6];
  assign io_out[5] = T49[5] | T1[5];
  assign io_out[4] = T49[4] | T1[4];
  assign io_out[3] = T49[3] | T1[3];
  assign io_out[2] = T49[2] | T1[2];
  assign io_out[1] = T49[1] | T1[1];
  assign io_out[0] = T49[0] | T1[0];
  assign T1[63] = T2[63] & io_lhs[63];
  assign T1[62] = T2[62] & io_lhs[62];
  assign T1[61] = T2[61] & io_lhs[61];
  assign T1[60] = T2[60] & io_lhs[60];
  assign T1[59] = T2[59] & io_lhs[59];
  assign T1[58] = T2[58] & io_lhs[58];
  assign T1[57] = T2[57] & io_lhs[57];
  assign T1[56] = T2[56] & io_lhs[56];
  assign T1[55] = T2[55] & io_lhs[55];
  assign T1[54] = T2[54] & io_lhs[54];
  assign T1[53] = T2[53] & io_lhs[53];
  assign T1[52] = T2[52] & io_lhs[52];
  assign T1[51] = T2[51] & io_lhs[51];
  assign T1[50] = T2[50] & io_lhs[50];
  assign T1[49] = T2[49] & io_lhs[49];
  assign T1[48] = T2[48] & io_lhs[48];
  assign T1[47] = T2[47] & io_lhs[47];
  assign T1[46] = T2[46] & io_lhs[46];
  assign T1[45] = T2[45] & io_lhs[45];
  assign T1[44] = T2[44] & io_lhs[44];
  assign T1[43] = T2[43] & io_lhs[43];
  assign T1[42] = T2[42] & io_lhs[42];
  assign T1[41] = T2[41] & io_lhs[41];
  assign T1[40] = T2[40] & io_lhs[40];
  assign T1[39] = T2[39] & io_lhs[39];
  assign T1[38] = T2[38] & io_lhs[38];
  assign T1[37] = T2[37] & io_lhs[37];
  assign T1[36] = T2[36] & io_lhs[36];
  assign T1[35] = T2[35] & io_lhs[35];
  assign T1[34] = T2[34] & io_lhs[34];
  assign T1[33] = T2[33] & io_lhs[33];
  assign T1[32] = T2[32] & io_lhs[32];
  assign T1[31] = T2[31] & io_lhs[31];
  assign T1[30] = T2[30] & io_lhs[30];
  assign T1[29] = T2[29] & io_lhs[29];
  assign T1[28] = T2[28] & io_lhs[28];
  assign T1[27] = T2[27] & io_lhs[27];
  assign T1[26] = T2[26] & io_lhs[26];
  assign T1[25] = T2[25] & io_lhs[25];
  assign T1[24] = T2[24] & io_lhs[24];
  assign T1[23] = T2[23] & io_lhs[23];
  assign T1[22] = T2[22] & io_lhs[22];
  assign T1[21] = T2[21] & io_lhs[21];
  assign T1[20] = T2[20] & io_lhs[20];
  assign T1[19] = T2[19] & io_lhs[19];
  assign T1[18] = T2[18] & io_lhs[18];
  assign T1[17] = T2[17] & io_lhs[17];
  assign T1[16] = T2[16] & io_lhs[16];
  assign T1[15] = T2[15] & io_lhs[15];
  assign T1[14] = T2[14] & io_lhs[14];
  assign T1[13] = T2[13] & io_lhs[13];
  assign T1[12] = T2[12] & io_lhs[12];
  assign T1[11] = T2[11] & io_lhs[11];
  assign T1[10] = T2[10] & io_lhs[10];
  assign T1[9] = T2[9] & io_lhs[9];
  assign T1[8] = T2[8] & io_lhs[8];
  assign T1[7] = T2[7] & io_lhs[7];
  assign T1[6] = T2[6] & io_lhs[6];
  assign T1[5] = T2[5] & io_lhs[5];
  assign T1[4] = T2[4] & io_lhs[4];
  assign T1[3] = T2[3] & io_lhs[3];
  assign T1[2] = T2[2] & io_lhs[2];
  assign T1[1] = T2[1] & io_lhs[1];
  assign T1[0] = T2[0] & io_lhs[0];
  assign T2[63] = ~wmask_63;
  assign T2[62] = ~wmask_63;
  assign T2[61] = ~wmask_63;
  assign T2[60] = ~wmask_63;
  assign T2[59] = ~wmask_63;
  assign T2[58] = ~wmask_63;
  assign T2[57] = ~wmask_63;
  assign T2[56] = ~wmask[56];
  assign T2[55] = ~wmask[55];
  assign T2[54] = ~wmask[55];
  assign T2[53] = ~wmask[55];
  assign T2[52] = ~wmask[55];
  assign T2[51] = ~wmask[55];
  assign T2[50] = ~wmask[55];
  assign T2[49] = ~wmask[55];
  assign T2[48] = ~wmask_48;
  assign T2[47] = ~wmask_47;
  assign T2[46] = ~wmask_47;
  assign T2[45] = ~wmask_47;
  assign T2[44] = ~wmask_47;
  assign T2[43] = ~wmask_47;
  assign T2[42] = ~wmask_47;
  assign T2[41] = ~wmask_47;
  assign T2[40] = ~wmask_40;
  assign T2[39] = ~wmask_39;
  assign T2[38] = ~wmask_39;
  assign T2[37] = ~wmask_39;
  assign T2[36] = ~wmask_39;
  assign T2[35] = ~wmask_39;
  assign T2[34] = ~wmask_39;
  assign T2[33] = ~wmask_39;
  assign T2[32] = ~wmask_32;
  assign T2[31] = ~wmask_31;
  assign T2[30] = ~wmask_31;
  assign T2[29] = ~wmask_31;
  assign T2[28] = ~wmask_31;
  assign T2[27] = ~wmask_31;
  assign T2[26] = ~wmask_31;
  assign T2[25] = ~wmask_31;
  assign T2[24] = ~wmask_24;
  assign T2[23] = ~wmask_23;
  assign T2[22] = ~wmask_23;
  assign T2[21] = ~wmask_23;
  assign T2[20] = ~wmask_23;
  assign T2[19] = ~wmask_23;
  assign T2[18] = ~wmask_23;
  assign T2[17] = ~wmask_23;
  assign T2[16] = ~wmask_16;
  assign T2[15] = ~wmask_15;
  assign T2[14] = ~wmask_15;
  assign T2[13] = ~wmask_15;
  assign T2[12] = ~wmask_15;
  assign T2[11] = ~wmask_15;
  assign T2[10] = ~wmask_15;
  assign T2[9] = ~wmask_15;
  assign T2[8] = ~wmask_8;
  assign T2[7] = ~wmask_7;
  assign T2[6] = ~wmask_7;
  assign T2[5] = ~wmask_7;
  assign T2[4] = ~wmask_7;
  assign T2[3] = ~wmask_7;
  assign T2[2] = ~wmask_7;
  assign T2[1] = ~wmask_7;
  assign T2[0] = ~wmask_0;
  assign N33 = ~io_addr[2];
  assign N34 = ~io_addr[1];
  assign T12[1] = io_addr[0] | T16;
  assign T16 = io_typ[1] | io_typ[0];
  assign T10[3] = T23[1] | T21[1];
  assign T10[2] = T23[0] | T21[1];
  assign T21[1] = io_typ[1];
  assign T8[7] = T29[3] | T27[3];
  assign T8[6] = T29[2] | T27[3];
  assign T8[5] = T29[1] | T27[3];
  assign T8[4] = T29[0] | T27[3];
  assign T27[3] = T28;
  assign T49[63] = wmask_63 & out[63];
  assign T49[62] = wmask_63 & out[62];
  assign T49[61] = wmask_63 & out[61];
  assign T49[60] = wmask_63 & out[60];
  assign T49[59] = wmask_63 & out[59];
  assign T49[58] = wmask_63 & out[58];
  assign T49[57] = wmask_63 & out[57];
  assign T49[56] = wmask[56] & out[56];
  assign T49[55] = wmask[55] & out[55];
  assign T49[54] = wmask[55] & out[54];
  assign T49[53] = wmask[55] & out[53];
  assign T49[52] = wmask[55] & out[52];
  assign T49[51] = wmask[55] & out[51];
  assign T49[50] = wmask[55] & out[50];
  assign T49[49] = wmask[55] & out[49];
  assign T49[48] = wmask_48 & out[48];
  assign T49[47] = wmask_47 & out[47];
  assign T49[46] = wmask_47 & out[46];
  assign T49[45] = wmask_47 & out[45];
  assign T49[44] = wmask_47 & out[44];
  assign T49[43] = wmask_47 & out[43];
  assign T49[42] = wmask_47 & out[42];
  assign T49[41] = wmask_47 & out[41];
  assign T49[40] = wmask_40 & out[40];
  assign T49[39] = wmask_39 & out[39];
  assign T49[38] = wmask_39 & out[38];
  assign T49[37] = wmask_39 & out[37];
  assign T49[36] = wmask_39 & out[36];
  assign T49[35] = wmask_39 & out[35];
  assign T49[34] = wmask_39 & out[34];
  assign T49[33] = wmask_39 & out[33];
  assign T49[32] = wmask_32 & out[32];
  assign T49[31] = wmask_31 & out[31];
  assign T49[30] = wmask_31 & out[30];
  assign T49[29] = wmask_31 & out[29];
  assign T49[28] = wmask_31 & out[28];
  assign T49[27] = wmask_31 & out[27];
  assign T49[26] = wmask_31 & out[26];
  assign T49[25] = wmask_31 & out[25];
  assign T49[24] = wmask_24 & out[24];
  assign T49[23] = wmask_23 & out[23];
  assign T49[22] = wmask_23 & out[22];
  assign T49[21] = wmask_23 & out[21];
  assign T49[20] = wmask_23 & out[20];
  assign T49[19] = wmask_23 & out[19];
  assign T49[18] = wmask_23 & out[18];
  assign T49[17] = wmask_23 & out[17];
  assign T49[16] = wmask_16 & out[16];
  assign T49[15] = wmask_15 & out[15];
  assign T49[14] = wmask_15 & out[14];
  assign T49[13] = wmask_15 & out[13];
  assign T49[12] = wmask_15 & out[12];
  assign T49[11] = wmask_15 & out[11];
  assign T49[10] = wmask_15 & out[10];
  assign T49[9] = wmask_15 & out[9];
  assign T49[8] = wmask_8 & out[8];
  assign T49[7] = wmask_7 & out[7];
  assign T49[6] = wmask_7 & out[6];
  assign T49[5] = wmask_7 & out[5];
  assign T49[4] = wmask_7 & out[4];
  assign T49[3] = wmask_7 & out[3];
  assign T49[2] = wmask_7 & out[2];
  assign T49[1] = wmask_7 & out[1];
  assign T49[0] = wmask_0 & out[0];
  assign N35 = ~T69;
  assign N36 = ~less;
  assign max = N72 | N74;
  assign min = N67 | N70;
  assign N37 = ~T106;
  assign N38 = ~sgned;
  assign N39 = ~T80;
  assign T80 = word & T81;
  assign T81 = ~io_addr[2];
  assign word = T84 | N81;
  assign T84 = T86 | N84;
  assign T86 = N87 | N90;
  assign N40 = ~T91;
  assign T91 = word & T92;
  assign T92 = ~io_addr[2];
  assign sgned = N67 | N72;
  assign N41 = ~word;
  assign T96 = lt_hi | T97;
  assign T97 = eq_hi & lt_lo;
  assign T107[63] = io_lhs[63] ^ rhs[63];
  assign T107[62] = io_lhs[62] ^ rhs[62];
  assign T107[61] = io_lhs[61] ^ rhs[61];
  assign T107[60] = io_lhs[60] ^ rhs[60];
  assign T107[59] = io_lhs[59] ^ rhs[59];
  assign T107[58] = io_lhs[58] ^ rhs[58];
  assign T107[57] = io_lhs[57] ^ rhs[57];
  assign T107[56] = io_lhs[56] ^ rhs[56];
  assign T107[55] = io_lhs[55] ^ rhs[55];
  assign T107[54] = io_lhs[54] ^ rhs[54];
  assign T107[53] = io_lhs[53] ^ rhs[53];
  assign T107[52] = io_lhs[52] ^ rhs[52];
  assign T107[51] = io_lhs[51] ^ rhs[51];
  assign T107[50] = io_lhs[50] ^ rhs[50];
  assign T107[49] = io_lhs[49] ^ rhs[49];
  assign T107[48] = io_lhs[48] ^ rhs[48];
  assign T107[47] = io_lhs[47] ^ rhs[47];
  assign T107[46] = io_lhs[46] ^ rhs[46];
  assign T107[45] = io_lhs[45] ^ rhs[45];
  assign T107[44] = io_lhs[44] ^ rhs[44];
  assign T107[43] = io_lhs[43] ^ rhs[43];
  assign T107[42] = io_lhs[42] ^ rhs[42];
  assign T107[41] = io_lhs[41] ^ rhs[41];
  assign T107[40] = io_lhs[40] ^ rhs[40];
  assign T107[39] = io_lhs[39] ^ rhs[39];
  assign T107[38] = io_lhs[38] ^ rhs[38];
  assign T107[37] = io_lhs[37] ^ rhs[37];
  assign T107[36] = io_lhs[36] ^ rhs[36];
  assign T107[35] = io_lhs[35] ^ rhs[35];
  assign T107[34] = io_lhs[34] ^ rhs[34];
  assign T107[33] = io_lhs[33] ^ rhs[33];
  assign T107[32] = io_lhs[32] ^ rhs[32];
  assign T107[31] = io_lhs[31] ^ io_rhs[31];
  assign T107[30] = io_lhs[30] ^ io_rhs[30];
  assign T107[29] = io_lhs[29] ^ io_rhs[29];
  assign T107[28] = io_lhs[28] ^ io_rhs[28];
  assign T107[27] = io_lhs[27] ^ io_rhs[27];
  assign T107[26] = io_lhs[26] ^ io_rhs[26];
  assign T107[25] = io_lhs[25] ^ io_rhs[25];
  assign T107[24] = io_lhs[24] ^ io_rhs[24];
  assign T107[23] = io_lhs[23] ^ io_rhs[23];
  assign T107[22] = io_lhs[22] ^ io_rhs[22];
  assign T107[21] = io_lhs[21] ^ io_rhs[21];
  assign T107[20] = io_lhs[20] ^ io_rhs[20];
  assign T107[19] = io_lhs[19] ^ io_rhs[19];
  assign T107[18] = io_lhs[18] ^ io_rhs[18];
  assign T107[17] = io_lhs[17] ^ io_rhs[17];
  assign T107[16] = io_lhs[16] ^ io_rhs[16];
  assign T107[15] = io_lhs[15] ^ io_rhs[15];
  assign T107[14] = io_lhs[14] ^ io_rhs[14];
  assign T107[13] = io_lhs[13] ^ io_rhs[13];
  assign T107[12] = io_lhs[12] ^ io_rhs[12];
  assign T107[11] = io_lhs[11] ^ io_rhs[11];
  assign T107[10] = io_lhs[10] ^ io_rhs[10];
  assign T107[9] = io_lhs[9] ^ io_rhs[9];
  assign T107[8] = io_lhs[8] ^ io_rhs[8];
  assign T107[7] = io_lhs[7] ^ io_rhs[7];
  assign T107[6] = io_lhs[6] ^ io_rhs[6];
  assign T107[5] = io_lhs[5] ^ io_rhs[5];
  assign T107[4] = io_lhs[4] ^ io_rhs[4];
  assign T107[3] = io_lhs[3] ^ io_rhs[3];
  assign T107[2] = io_lhs[2] ^ io_rhs[2];
  assign T107[1] = io_lhs[1] ^ io_rhs[1];
  assign T107[0] = io_lhs[0] ^ io_rhs[0];
  assign T109[63] = io_lhs[63] | rhs[63];
  assign T109[62] = io_lhs[62] | rhs[62];
  assign T109[61] = io_lhs[61] | rhs[61];
  assign T109[60] = io_lhs[60] | rhs[60];
  assign T109[59] = io_lhs[59] | rhs[59];
  assign T109[58] = io_lhs[58] | rhs[58];
  assign T109[57] = io_lhs[57] | rhs[57];
  assign T109[56] = io_lhs[56] | rhs[56];
  assign T109[55] = io_lhs[55] | rhs[55];
  assign T109[54] = io_lhs[54] | rhs[54];
  assign T109[53] = io_lhs[53] | rhs[53];
  assign T109[52] = io_lhs[52] | rhs[52];
  assign T109[51] = io_lhs[51] | rhs[51];
  assign T109[50] = io_lhs[50] | rhs[50];
  assign T109[49] = io_lhs[49] | rhs[49];
  assign T109[48] = io_lhs[48] | rhs[48];
  assign T109[47] = io_lhs[47] | rhs[47];
  assign T109[46] = io_lhs[46] | rhs[46];
  assign T109[45] = io_lhs[45] | rhs[45];
  assign T109[44] = io_lhs[44] | rhs[44];
  assign T109[43] = io_lhs[43] | rhs[43];
  assign T109[42] = io_lhs[42] | rhs[42];
  assign T109[41] = io_lhs[41] | rhs[41];
  assign T109[40] = io_lhs[40] | rhs[40];
  assign T109[39] = io_lhs[39] | rhs[39];
  assign T109[38] = io_lhs[38] | rhs[38];
  assign T109[37] = io_lhs[37] | rhs[37];
  assign T109[36] = io_lhs[36] | rhs[36];
  assign T109[35] = io_lhs[35] | rhs[35];
  assign T109[34] = io_lhs[34] | rhs[34];
  assign T109[33] = io_lhs[33] | rhs[33];
  assign T109[32] = io_lhs[32] | rhs[32];
  assign T109[31] = io_lhs[31] | io_rhs[31];
  assign T109[30] = io_lhs[30] | io_rhs[30];
  assign T109[29] = io_lhs[29] | io_rhs[29];
  assign T109[28] = io_lhs[28] | io_rhs[28];
  assign T109[27] = io_lhs[27] | io_rhs[27];
  assign T109[26] = io_lhs[26] | io_rhs[26];
  assign T109[25] = io_lhs[25] | io_rhs[25];
  assign T109[24] = io_lhs[24] | io_rhs[24];
  assign T109[23] = io_lhs[23] | io_rhs[23];
  assign T109[22] = io_lhs[22] | io_rhs[22];
  assign T109[21] = io_lhs[21] | io_rhs[21];
  assign T109[20] = io_lhs[20] | io_rhs[20];
  assign T109[19] = io_lhs[19] | io_rhs[19];
  assign T109[18] = io_lhs[18] | io_rhs[18];
  assign T109[17] = io_lhs[17] | io_rhs[17];
  assign T109[16] = io_lhs[16] | io_rhs[16];
  assign T109[15] = io_lhs[15] | io_rhs[15];
  assign T109[14] = io_lhs[14] | io_rhs[14];
  assign T109[13] = io_lhs[13] | io_rhs[13];
  assign T109[12] = io_lhs[12] | io_rhs[12];
  assign T109[11] = io_lhs[11] | io_rhs[11];
  assign T109[10] = io_lhs[10] | io_rhs[10];
  assign T109[9] = io_lhs[9] | io_rhs[9];
  assign T109[8] = io_lhs[8] | io_rhs[8];
  assign T109[7] = io_lhs[7] | io_rhs[7];
  assign T109[6] = io_lhs[6] | io_rhs[6];
  assign T109[5] = io_lhs[5] | io_rhs[5];
  assign T109[4] = io_lhs[4] | io_rhs[4];
  assign T109[3] = io_lhs[3] | io_rhs[3];
  assign T109[2] = io_lhs[2] | io_rhs[2];
  assign T109[1] = io_lhs[1] | io_rhs[1];
  assign T109[0] = io_lhs[0] | io_rhs[0];
  assign T111[63] = io_lhs[63] & rhs[63];
  assign T111[62] = io_lhs[62] & rhs[62];
  assign T111[61] = io_lhs[61] & rhs[61];
  assign T111[60] = io_lhs[60] & rhs[60];
  assign T111[59] = io_lhs[59] & rhs[59];
  assign T111[58] = io_lhs[58] & rhs[58];
  assign T111[57] = io_lhs[57] & rhs[57];
  assign T111[56] = io_lhs[56] & rhs[56];
  assign T111[55] = io_lhs[55] & rhs[55];
  assign T111[54] = io_lhs[54] & rhs[54];
  assign T111[53] = io_lhs[53] & rhs[53];
  assign T111[52] = io_lhs[52] & rhs[52];
  assign T111[51] = io_lhs[51] & rhs[51];
  assign T111[50] = io_lhs[50] & rhs[50];
  assign T111[49] = io_lhs[49] & rhs[49];
  assign T111[48] = io_lhs[48] & rhs[48];
  assign T111[47] = io_lhs[47] & rhs[47];
  assign T111[46] = io_lhs[46] & rhs[46];
  assign T111[45] = io_lhs[45] & rhs[45];
  assign T111[44] = io_lhs[44] & rhs[44];
  assign T111[43] = io_lhs[43] & rhs[43];
  assign T111[42] = io_lhs[42] & rhs[42];
  assign T111[41] = io_lhs[41] & rhs[41];
  assign T111[40] = io_lhs[40] & rhs[40];
  assign T111[39] = io_lhs[39] & rhs[39];
  assign T111[38] = io_lhs[38] & rhs[38];
  assign T111[37] = io_lhs[37] & rhs[37];
  assign T111[36] = io_lhs[36] & rhs[36];
  assign T111[35] = io_lhs[35] & rhs[35];
  assign T111[34] = io_lhs[34] & rhs[34];
  assign T111[33] = io_lhs[33] & rhs[33];
  assign T111[32] = io_lhs[32] & rhs[32];
  assign T111[31] = io_lhs[31] & io_rhs[31];
  assign T111[30] = io_lhs[30] & io_rhs[30];
  assign T111[29] = io_lhs[29] & io_rhs[29];
  assign T111[28] = io_lhs[28] & io_rhs[28];
  assign T111[27] = io_lhs[27] & io_rhs[27];
  assign T111[26] = io_lhs[26] & io_rhs[26];
  assign T111[25] = io_lhs[25] & io_rhs[25];
  assign T111[24] = io_lhs[24] & io_rhs[24];
  assign T111[23] = io_lhs[23] & io_rhs[23];
  assign T111[22] = io_lhs[22] & io_rhs[22];
  assign T111[21] = io_lhs[21] & io_rhs[21];
  assign T111[20] = io_lhs[20] & io_rhs[20];
  assign T111[19] = io_lhs[19] & io_rhs[19];
  assign T111[18] = io_lhs[18] & io_rhs[18];
  assign T111[17] = io_lhs[17] & io_rhs[17];
  assign T111[16] = io_lhs[16] & io_rhs[16];
  assign T111[15] = io_lhs[15] & io_rhs[15];
  assign T111[14] = io_lhs[14] & io_rhs[14];
  assign T111[13] = io_lhs[13] & io_rhs[13];
  assign T111[12] = io_lhs[12] & io_rhs[12];
  assign T111[11] = io_lhs[11] & io_rhs[11];
  assign T111[10] = io_lhs[10] & io_rhs[10];
  assign T111[9] = io_lhs[9] & io_rhs[9];
  assign T111[8] = io_lhs[8] & io_rhs[8];
  assign T111[7] = io_lhs[7] & io_rhs[7];
  assign T111[6] = io_lhs[6] & io_rhs[6];
  assign T111[5] = io_lhs[5] & io_rhs[5];
  assign T111[4] = io_lhs[4] & io_rhs[4];
  assign T111[3] = io_lhs[3] & io_rhs[3];
  assign T111[2] = io_lhs[2] & io_rhs[2];
  assign T111[1] = io_lhs[1] & io_rhs[1];
  assign T111[0] = io_lhs[0] & io_rhs[0];
  assign T113[63] = rhs[63] & mask[63];
  assign T113[62] = rhs[62] & mask[62];
  assign T113[61] = rhs[61] & mask[61];
  assign T113[60] = rhs[60] & mask[60];
  assign T113[59] = rhs[59] & mask[59];
  assign T113[58] = rhs[58] & mask[58];
  assign T113[57] = rhs[57] & mask[57];
  assign T113[56] = rhs[56] & mask[56];
  assign T113[55] = rhs[55] & mask[55];
  assign T113[54] = rhs[54] & mask[54];
  assign T113[53] = rhs[53] & mask[53];
  assign T113[52] = rhs[52] & mask[52];
  assign T113[51] = rhs[51] & mask[51];
  assign T113[50] = rhs[50] & mask[50];
  assign T113[49] = rhs[49] & mask[49];
  assign T113[48] = rhs[48] & mask[48];
  assign T113[47] = rhs[47] & mask[47];
  assign T113[46] = rhs[46] & mask[46];
  assign T113[45] = rhs[45] & mask[45];
  assign T113[44] = rhs[44] & mask[44];
  assign T113[43] = rhs[43] & mask[43];
  assign T113[42] = rhs[42] & mask[42];
  assign T113[41] = rhs[41] & mask[41];
  assign T113[40] = rhs[40] & mask[40];
  assign T113[39] = rhs[39] & mask[39];
  assign T113[38] = rhs[38] & mask[38];
  assign T113[37] = rhs[37] & mask[37];
  assign T113[36] = rhs[36] & mask[36];
  assign T113[35] = rhs[35] & mask[35];
  assign T113[34] = rhs[34] & mask[34];
  assign T113[33] = rhs[33] & mask[33];
  assign T113[32] = rhs[32] & mask[32];
  assign T113[31] = io_rhs[31] & mask[31];
  assign T113[30] = io_rhs[30] & mask[30];
  assign T113[29] = io_rhs[29] & mask[29];
  assign T113[28] = io_rhs[28] & mask[28];
  assign T113[27] = io_rhs[27] & mask[27];
  assign T113[26] = io_rhs[26] & mask[26];
  assign T113[25] = io_rhs[25] & mask[25];
  assign T113[24] = io_rhs[24] & mask[24];
  assign T113[23] = io_rhs[23] & mask[23];
  assign T113[22] = io_rhs[22] & mask[22];
  assign T113[21] = io_rhs[21] & mask[21];
  assign T113[20] = io_rhs[20] & mask[20];
  assign T113[19] = io_rhs[19] & mask[19];
  assign T113[18] = io_rhs[18] & mask[18];
  assign T113[17] = io_rhs[17] & mask[17];
  assign T113[16] = io_rhs[16] & mask[16];
  assign T113[15] = io_rhs[15] & mask[15];
  assign T113[14] = io_rhs[14] & mask[14];
  assign T113[13] = io_rhs[13] & mask[13];
  assign T113[12] = io_rhs[12] & mask[12];
  assign T113[11] = io_rhs[11] & mask[11];
  assign T113[10] = io_rhs[10] & mask[10];
  assign T113[9] = io_rhs[9] & mask[9];
  assign T113[8] = io_rhs[8] & mask[8];
  assign T113[7] = io_rhs[7] & mask[7];
  assign T113[6] = io_rhs[6] & mask[6];
  assign T113[5] = io_rhs[5] & mask[5];
  assign T113[4] = io_rhs[4] & mask[4];
  assign T113[3] = io_rhs[3] & mask[3];
  assign T113[2] = io_rhs[2] & mask[2];
  assign T113[1] = io_rhs[1] & mask[1];
  assign T113[0] = io_rhs[0] & mask[0];
  assign mask[63] = ~1'b0;
  assign mask[62] = ~1'b0;
  assign mask[61] = ~1'b0;
  assign mask[60] = ~1'b0;
  assign mask[59] = ~1'b0;
  assign mask[58] = ~1'b0;
  assign mask[57] = ~1'b0;
  assign mask[56] = ~1'b0;
  assign mask[55] = ~1'b0;
  assign mask[54] = ~1'b0;
  assign mask[53] = ~1'b0;
  assign mask[52] = ~1'b0;
  assign mask[51] = ~1'b0;
  assign mask[50] = ~1'b0;
  assign mask[49] = ~1'b0;
  assign mask[48] = ~1'b0;
  assign mask[47] = ~1'b0;
  assign mask[46] = ~1'b0;
  assign mask[45] = ~1'b0;
  assign mask[44] = ~1'b0;
  assign mask[43] = ~1'b0;
  assign mask[42] = ~1'b0;
  assign mask[41] = ~1'b0;
  assign mask[40] = ~1'b0;
  assign mask[39] = ~1'b0;
  assign mask[38] = ~1'b0;
  assign mask[37] = ~1'b0;
  assign mask[36] = ~1'b0;
  assign mask[35] = ~1'b0;
  assign mask[34] = ~1'b0;
  assign mask[33] = ~1'b0;
  assign mask[32] = ~1'b0;
  assign mask[31] = ~io_addr[2];
  assign mask[30] = ~1'b0;
  assign mask[29] = ~1'b0;
  assign mask[28] = ~1'b0;
  assign mask[27] = ~1'b0;
  assign mask[26] = ~1'b0;
  assign mask[25] = ~1'b0;
  assign mask[24] = ~1'b0;
  assign mask[23] = ~1'b0;
  assign mask[22] = ~1'b0;
  assign mask[21] = ~1'b0;
  assign mask[20] = ~1'b0;
  assign mask[19] = ~1'b0;
  assign mask[18] = ~1'b0;
  assign mask[17] = ~1'b0;
  assign mask[16] = ~1'b0;
  assign mask[15] = ~1'b0;
  assign mask[14] = ~1'b0;
  assign mask[13] = ~1'b0;
  assign mask[12] = ~1'b0;
  assign mask[11] = ~1'b0;
  assign mask[10] = ~1'b0;
  assign mask[9] = ~1'b0;
  assign mask[8] = ~1'b0;
  assign mask[7] = ~1'b0;
  assign mask[6] = ~1'b0;
  assign mask[5] = ~1'b0;
  assign mask[4] = ~1'b0;
  assign mask[3] = ~1'b0;
  assign mask[2] = ~1'b0;
  assign mask[1] = ~1'b0;
  assign mask[0] = ~1'b0;
  assign T116[63] = io_lhs[63] & mask[63];
  assign T116[62] = io_lhs[62] & mask[62];
  assign T116[61] = io_lhs[61] & mask[61];
  assign T116[60] = io_lhs[60] & mask[60];
  assign T116[59] = io_lhs[59] & mask[59];
  assign T116[58] = io_lhs[58] & mask[58];
  assign T116[57] = io_lhs[57] & mask[57];
  assign T116[56] = io_lhs[56] & mask[56];
  assign T116[55] = io_lhs[55] & mask[55];
  assign T116[54] = io_lhs[54] & mask[54];
  assign T116[53] = io_lhs[53] & mask[53];
  assign T116[52] = io_lhs[52] & mask[52];
  assign T116[51] = io_lhs[51] & mask[51];
  assign T116[50] = io_lhs[50] & mask[50];
  assign T116[49] = io_lhs[49] & mask[49];
  assign T116[48] = io_lhs[48] & mask[48];
  assign T116[47] = io_lhs[47] & mask[47];
  assign T116[46] = io_lhs[46] & mask[46];
  assign T116[45] = io_lhs[45] & mask[45];
  assign T116[44] = io_lhs[44] & mask[44];
  assign T116[43] = io_lhs[43] & mask[43];
  assign T116[42] = io_lhs[42] & mask[42];
  assign T116[41] = io_lhs[41] & mask[41];
  assign T116[40] = io_lhs[40] & mask[40];
  assign T116[39] = io_lhs[39] & mask[39];
  assign T116[38] = io_lhs[38] & mask[38];
  assign T116[37] = io_lhs[37] & mask[37];
  assign T116[36] = io_lhs[36] & mask[36];
  assign T116[35] = io_lhs[35] & mask[35];
  assign T116[34] = io_lhs[34] & mask[34];
  assign T116[33] = io_lhs[33] & mask[33];
  assign T116[32] = io_lhs[32] & mask[32];
  assign T116[31] = io_lhs[31] & mask[31];
  assign T116[30] = io_lhs[30] & mask[30];
  assign T116[29] = io_lhs[29] & mask[29];
  assign T116[28] = io_lhs[28] & mask[28];
  assign T116[27] = io_lhs[27] & mask[27];
  assign T116[26] = io_lhs[26] & mask[26];
  assign T116[25] = io_lhs[25] & mask[25];
  assign T116[24] = io_lhs[24] & mask[24];
  assign T116[23] = io_lhs[23] & mask[23];
  assign T116[22] = io_lhs[22] & mask[22];
  assign T116[21] = io_lhs[21] & mask[21];
  assign T116[20] = io_lhs[20] & mask[20];
  assign T116[19] = io_lhs[19] & mask[19];
  assign T116[18] = io_lhs[18] & mask[18];
  assign T116[17] = io_lhs[17] & mask[17];
  assign T116[16] = io_lhs[16] & mask[16];
  assign T116[15] = io_lhs[15] & mask[15];
  assign T116[14] = io_lhs[14] & mask[14];
  assign T116[13] = io_lhs[13] & mask[13];
  assign T116[12] = io_lhs[12] & mask[12];
  assign T116[11] = io_lhs[11] & mask[11];
  assign T116[10] = io_lhs[10] & mask[10];
  assign T116[9] = io_lhs[9] & mask[9];
  assign T116[8] = io_lhs[8] & mask[8];
  assign T116[7] = io_lhs[7] & mask[7];
  assign T116[6] = io_lhs[6] & mask[6];
  assign T116[5] = io_lhs[5] & mask[5];
  assign T116[4] = io_lhs[4] & mask[4];
  assign T116[3] = io_lhs[3] & mask[3];
  assign T116[2] = io_lhs[2] & mask[2];
  assign T116[1] = io_lhs[1] & mask[1];
  assign T116[0] = io_lhs[0] & mask[0];

endmodule