module cache_ctrl_0000000080000000
(
  clk_i,
  rst_ni,
  flush_i,
  bypass_i,
  busy_o,
  req_port_i,
  req_port_o,
  req_o,
  addr_o,
  gnt_i,
  data_o,
  be_o,
  tag_o,
  data_i,
  we_o,
  hit_way_i,
  miss_req_o,
  miss_gnt_i,
  active_serving_i,
  critical_word_i,
  critical_word_valid_i,
  bypass_gnt_i,
  bypass_valid_i,
  bypass_data_i,
  mshr_addr_o,
  mshr_addr_matches_i,
  mshr_index_matches_i
);

  input [133:0] req_port_i;
  output [65:0] req_port_o;
  output [7:0] req_o;
  output [11:0] addr_o;
  output [173:0] data_o;
  output [29:0] be_o;
  output [43:0] tag_o;
  input [1391:0] data_i;
  input [7:0] hit_way_i;
  output [140:0] miss_req_o;
  input [63:0] critical_word_i;
  input [63:0] bypass_data_i;
  output [55:0] mshr_addr_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input bypass_i;
  input gnt_i;
  input miss_gnt_i;
  input active_serving_i;
  input critical_word_valid_i;
  input bypass_gnt_i;
  input bypass_valid_i;
  input mshr_addr_matches_i;
  input mshr_index_matches_i;
  output busy_o;
  output we_o;
  wire [65:0] req_port_o;
  wire [7:0] req_o,hit_way_d;
  wire [11:0] addr_o;
  wire [173:0] data_o;
  wire [29:0] be_o;
  wire [43:0] tag_o;
  wire [140:0] miss_req_o;
  wire [55:0] mshr_addr_o;
  wire busy_o,we_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,
  N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,
  N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,
  N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,
  N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,
  N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
  N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,
  N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,
  N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,
  N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,
  N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,
  N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
  N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,
  N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,
  N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,
  N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,
  N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,
  N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,
  N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,
  N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,
  N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,
  N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
  N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,
  N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,
  N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,
  N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,
  N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,
  N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
  N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,
  N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,
  N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,
  N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,
  N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,
  N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,
  N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,
  N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,
  N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,
  N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,
  N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,
  N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,
  N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,
  N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,
  N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,
  N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,
  N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,
  N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,
  N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,
  N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,
  N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,
  N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,
  N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,
  N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,
  N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,
  N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,
  N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,
  N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,
  N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,
  N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,
  N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,
  N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,
  N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,
  N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,
  N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,
  N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,
  N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
  N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,
  N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,
  N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,
  N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,
  N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
  N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,
  N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,
  N1556,N1557,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,
  N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,
  N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,
  N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,
  N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,
  N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,
  N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,
  N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,
  N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,
  N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,
  N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,
  N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,
  N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,
  N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,
  N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,
  N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,
  N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,
  N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,
  N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,
  N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,
  N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,
  N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
  N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,
  N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,
  N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,
  N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,
  N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,
  N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,
  N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,
  N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,
  N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,
  N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,
  N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,
  N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,
  N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,
  N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,
  N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,
  N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,
  N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,
  N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,
  N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,
  N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,
  N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,
  N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,
  N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,
  N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,
  N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,
  N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,
  N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248;
  wire [127:0] cl_i;
  wire [3:0] state_d;
  wire [131:0] mem_req_d;
  reg [7:0] hit_way_q;
  reg [3:0] state_q;
  reg mem_req_q_index__11_,mem_req_q_index__10_,mem_req_q_index__9_,
  mem_req_q_index__8_,mem_req_q_index__7_,mem_req_q_index__6_,mem_req_q_index__5_,
  mem_req_q_index__4_,N1558,mem_req_q_index__2_,mem_req_q_index__1_,mem_req_q_index__0_,
  mem_req_q_tag__43_,mem_req_q_tag__42_,mem_req_q_tag__41_,mem_req_q_tag__40_,
  mem_req_q_tag__39_,mem_req_q_tag__38_,mem_req_q_tag__37_,mem_req_q_tag__36_,mem_req_q_tag__35_,
  mem_req_q_tag__34_,mem_req_q_tag__33_,mem_req_q_tag__32_,mem_req_q_tag__31_,
  mem_req_q_tag__30_,mem_req_q_tag__29_,mem_req_q_tag__28_,mem_req_q_tag__27_,
  mem_req_q_tag__26_,mem_req_q_tag__25_,mem_req_q_tag__24_,mem_req_q_tag__23_,
  mem_req_q_tag__22_,mem_req_q_tag__21_,mem_req_q_tag__20_,mem_req_q_tag__19_,
  mem_req_q_tag__18_,mem_req_q_tag__17_,mem_req_q_tag__16_,mem_req_q_tag__15_,mem_req_q_tag__14_,
  mem_req_q_tag__13_,mem_req_q_tag__12_,mem_req_q_tag__11_,mem_req_q_tag__10_,
  mem_req_q_tag__9_,mem_req_q_tag__8_,mem_req_q_tag__7_,mem_req_q_tag__6_,
  mem_req_q_tag__5_,mem_req_q_tag__4_,mem_req_q_tag__3_,mem_req_q_tag__2_,mem_req_q_tag__1_,
  mem_req_q_tag__0_,mem_req_q_be__7_,mem_req_q_be__6_,mem_req_q_be__5_,
  mem_req_q_be__4_,mem_req_q_be__3_,mem_req_q_be__2_,mem_req_q_be__1_,mem_req_q_be__0_,
  mem_req_q_size__1_,mem_req_q_size__0_,mem_req_q_we_,mem_req_q_wdata__63_,
  mem_req_q_wdata__62_,mem_req_q_wdata__61_,mem_req_q_wdata__60_,mem_req_q_wdata__59_,
  mem_req_q_wdata__58_,mem_req_q_wdata__57_,mem_req_q_wdata__56_,mem_req_q_wdata__55_,
  mem_req_q_wdata__54_,mem_req_q_wdata__53_,mem_req_q_wdata__52_,mem_req_q_wdata__51_,
  mem_req_q_wdata__50_,mem_req_q_wdata__49_,mem_req_q_wdata__48_,mem_req_q_wdata__47_,
  mem_req_q_wdata__46_,mem_req_q_wdata__45_,mem_req_q_wdata__44_,
  mem_req_q_wdata__43_,mem_req_q_wdata__42_,mem_req_q_wdata__41_,mem_req_q_wdata__40_,
  mem_req_q_wdata__39_,mem_req_q_wdata__38_,mem_req_q_wdata__37_,mem_req_q_wdata__36_,
  mem_req_q_wdata__35_,mem_req_q_wdata__34_,mem_req_q_wdata__33_,mem_req_q_wdata__32_,
  mem_req_q_wdata__31_,mem_req_q_wdata__30_,mem_req_q_wdata__29_,mem_req_q_wdata__28_,
  mem_req_q_wdata__27_,mem_req_q_wdata__26_,mem_req_q_wdata__25_,
  mem_req_q_wdata__24_,mem_req_q_wdata__23_,mem_req_q_wdata__22_,mem_req_q_wdata__21_,
  mem_req_q_wdata__20_,mem_req_q_wdata__19_,mem_req_q_wdata__18_,mem_req_q_wdata__17_,
  mem_req_q_wdata__16_,mem_req_q_wdata__15_,mem_req_q_wdata__14_,mem_req_q_wdata__13_,
  mem_req_q_wdata__12_,mem_req_q_wdata__11_,mem_req_q_wdata__10_,mem_req_q_wdata__9_,
  mem_req_q_wdata__8_,mem_req_q_wdata__7_,mem_req_q_wdata__6_,mem_req_q_wdata__5_,
  mem_req_q_wdata__4_,mem_req_q_wdata__3_,mem_req_q_wdata__2_,mem_req_q_wdata__1_,
  mem_req_q_wdata__0_,mem_req_q_bypass_;
  assign data_o[130] = 1'b0;
  assign data_o[131] = 1'b0;
  assign data_o[132] = 1'b0;
  assign data_o[133] = 1'b0;
  assign data_o[134] = 1'b0;
  assign data_o[135] = 1'b0;
  assign data_o[136] = 1'b0;
  assign data_o[137] = 1'b0;
  assign data_o[138] = 1'b0;
  assign data_o[139] = 1'b0;
  assign data_o[140] = 1'b0;
  assign data_o[141] = 1'b0;
  assign data_o[142] = 1'b0;
  assign data_o[143] = 1'b0;
  assign data_o[144] = 1'b0;
  assign data_o[145] = 1'b0;
  assign data_o[146] = 1'b0;
  assign data_o[147] = 1'b0;
  assign data_o[148] = 1'b0;
  assign data_o[149] = 1'b0;
  assign data_o[150] = 1'b0;
  assign data_o[151] = 1'b0;
  assign data_o[152] = 1'b0;
  assign data_o[153] = 1'b0;
  assign data_o[154] = 1'b0;
  assign data_o[155] = 1'b0;
  assign data_o[156] = 1'b0;
  assign data_o[157] = 1'b0;
  assign data_o[158] = 1'b0;
  assign data_o[159] = 1'b0;
  assign data_o[160] = 1'b0;
  assign data_o[161] = 1'b0;
  assign data_o[162] = 1'b0;
  assign data_o[163] = 1'b0;
  assign data_o[164] = 1'b0;
  assign data_o[165] = 1'b0;
  assign data_o[166] = 1'b0;
  assign data_o[167] = 1'b0;
  assign data_o[168] = 1'b0;
  assign data_o[169] = 1'b0;
  assign data_o[170] = 1'b0;
  assign data_o[171] = 1'b0;
  assign data_o[172] = 1'b0;
  assign data_o[173] = 1'b0;
  assign miss_req_o[132] = 1'b0;
  assign miss_req_o[133] = 1'b0;
  assign miss_req_o[134] = 1'b0;
  assign miss_req_o[135] = 1'b0;
  assign miss_req_o[136] = 1'b0;
  assign miss_req_o[137] = 1'b0;
  assign miss_req_o[138] = 1'b0;
  assign miss_req_o[139] = 1'b0;
  assign be_o[24] = 1'b0;
  assign be_o[25] = 1'b0;
  assign be_o[26] = 1'b0;
  assign be_o[27] = 1'b0;
  assign be_o[28] = 1'b0;
  assign be_o[29] = 1'b0;
  assign N953 = N951 & N2205;
  assign N954 = N2206 & N952;
  assign N955 = N953 & N954;
  assign N956 = state_q[3] | state_q[2];
  assign N957 = state_q[1] | N952;
  assign N958 = N956 | N957;
  assign N959 = state_q[3] | N2205;
  assign N960 = N2206 | state_q[0];
  assign N961 = N959 | N960;
  assign N963 = state_q[3] | state_q[2];
  assign N964 = N2206 | N952;
  assign N965 = N963 | N964;
  assign N967 = state_q[3] | N2205;
  assign N968 = N2206 | N952;
  assign N969 = N967 | N968;
  assign N971 = state_q[3] | state_q[2];
  assign N972 = N2206 | state_q[0];
  assign N973 = N971 | N972;
  assign N975 = state_q[3] | N2205;
  assign N976 = state_q[1] | N952;
  assign N977 = N975 | N976;
  assign N979 = N951 | state_q[2];
  assign N980 = state_q[1] | state_q[0];
  assign N981 = N979 | N980;
  assign N983 = state_q[3] | N2205;
  assign N984 = state_q[1] | state_q[0];
  assign N985 = N983 | N984;

  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[7] <= 1'b0;
    end else if(N2054) begin
      hit_way_q[7] <= hit_way_d[7];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[6] <= 1'b0;
    end else if(N2067) begin
      hit_way_q[6] <= hit_way_d[6];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[5] <= 1'b0;
    end else if(N2067) begin
      hit_way_q[5] <= hit_way_d[5];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[4] <= 1'b0;
    end else if(N2067) begin
      hit_way_q[4] <= hit_way_d[4];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[3] <= 1'b0;
    end else if(N2067) begin
      hit_way_q[3] <= hit_way_d[3];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[2] <= 1'b0;
    end else if(N2067) begin
      hit_way_q[2] <= hit_way_d[2];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[1] <= 1'b0;
    end else if(N2067) begin
      hit_way_q[1] <= hit_way_d[1];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      hit_way_q[0] <= 1'b0;
    end else if(N2067) begin
      hit_way_q[0] <= hit_way_d[0];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      state_q[3] <= 1'b0;
    end else if(N2100) begin
      state_q[3] <= state_d[3];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      state_q[2] <= 1'b0;
    end else if(N2100) begin
      state_q[2] <= state_d[2];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      state_q[1] <= 1'b0;
    end else if(N2100) begin
      state_q[1] <= state_d[1];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      state_q[0] <= 1'b0;
    end else if(N2100) begin
      state_q[0] <= state_d[0];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__11_ <= 1'b0;
    end else if(N2116) begin
      mem_req_q_index__11_ <= mem_req_d[131];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__10_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__10_ <= mem_req_d[130];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__9_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__9_ <= mem_req_d[129];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__8_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__8_ <= mem_req_d[128];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__7_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__7_ <= mem_req_d[127];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__6_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__6_ <= mem_req_d[126];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__5_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__5_ <= mem_req_d[125];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__4_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__4_ <= mem_req_d[124];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      N1558 <= 1'b0;
    end else if(N2131) begin
      N1558 <= mem_req_d[123];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__2_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__2_ <= mem_req_d[122];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__1_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__1_ <= mem_req_d[121];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_index__0_ <= 1'b0;
    end else if(N2131) begin
      mem_req_q_index__0_ <= mem_req_d[120];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__43_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__43_ <= mem_req_d[119];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__42_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__42_ <= mem_req_d[118];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__41_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__41_ <= mem_req_d[117];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__40_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__40_ <= mem_req_d[116];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__39_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__39_ <= mem_req_d[115];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__38_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__38_ <= mem_req_d[114];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__37_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__37_ <= mem_req_d[113];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__36_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__36_ <= mem_req_d[112];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__35_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__35_ <= mem_req_d[111];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__34_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__34_ <= mem_req_d[110];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__33_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__33_ <= mem_req_d[109];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__32_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__32_ <= mem_req_d[108];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__31_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__31_ <= mem_req_d[107];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__30_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__30_ <= mem_req_d[106];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__29_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__29_ <= mem_req_d[105];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__28_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__28_ <= mem_req_d[104];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__27_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__27_ <= mem_req_d[103];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__26_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__26_ <= mem_req_d[102];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__25_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__25_ <= mem_req_d[101];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__24_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__24_ <= mem_req_d[100];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__23_ <= 1'b0;
    end else if(N2141) begin
      mem_req_q_tag__23_ <= mem_req_d[99];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__22_ <= 1'b0;
    end else if(N2150) begin
      mem_req_q_tag__22_ <= mem_req_d[98];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__21_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__21_ <= mem_req_d[97];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__20_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__20_ <= mem_req_d[96];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__19_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__19_ <= mem_req_d[95];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__18_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__18_ <= mem_req_d[94];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__17_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__17_ <= mem_req_d[93];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__16_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__16_ <= mem_req_d[92];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__15_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__15_ <= mem_req_d[91];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__14_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__14_ <= mem_req_d[90];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__13_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__13_ <= mem_req_d[89];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__12_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__12_ <= mem_req_d[88];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__11_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__11_ <= mem_req_d[87];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__10_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__10_ <= mem_req_d[86];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__9_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__9_ <= mem_req_d[85];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__8_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__8_ <= mem_req_d[84];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__7_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__7_ <= mem_req_d[83];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__6_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__6_ <= mem_req_d[82];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__5_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__5_ <= mem_req_d[81];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__4_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__4_ <= mem_req_d[80];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__3_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__3_ <= mem_req_d[79];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__2_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__2_ <= mem_req_d[78];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__1_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__1_ <= mem_req_d[77];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_tag__0_ <= 1'b0;
    end else if(N2154) begin
      mem_req_q_tag__0_ <= mem_req_d[76];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__7_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__7_ <= mem_req_d[75];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__6_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__6_ <= mem_req_d[74];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__5_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__5_ <= mem_req_d[73];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__4_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__4_ <= mem_req_d[72];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__3_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__3_ <= mem_req_d[71];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__2_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__2_ <= mem_req_d[70];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__1_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__1_ <= mem_req_d[69];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_be__0_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_be__0_ <= mem_req_d[68];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_size__1_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_size__1_ <= mem_req_d[67];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_size__0_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_size__0_ <= mem_req_d[66];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_we_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_we_ <= mem_req_d[65];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__63_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__63_ <= mem_req_d[64];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__62_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__62_ <= mem_req_d[63];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__61_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__61_ <= mem_req_d[62];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__60_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__60_ <= mem_req_d[61];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__59_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__59_ <= mem_req_d[60];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__58_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__58_ <= mem_req_d[59];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__57_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__57_ <= mem_req_d[58];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__56_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__56_ <= mem_req_d[57];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__55_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__55_ <= mem_req_d[56];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__54_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__54_ <= mem_req_d[55];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__53_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__53_ <= mem_req_d[54];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__52_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__52_ <= mem_req_d[53];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__51_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__51_ <= mem_req_d[52];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__50_ <= 1'b0;
    end else if(N2163) begin
      mem_req_q_wdata__50_ <= mem_req_d[51];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__49_ <= 1'b0;
    end else if(N2174) begin
      mem_req_q_wdata__49_ <= mem_req_d[50];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__48_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__48_ <= mem_req_d[49];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__47_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__47_ <= mem_req_d[48];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__46_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__46_ <= mem_req_d[47];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__45_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__45_ <= mem_req_d[46];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__44_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__44_ <= mem_req_d[45];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__43_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__43_ <= mem_req_d[44];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__42_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__42_ <= mem_req_d[43];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__41_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__41_ <= mem_req_d[42];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__40_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__40_ <= mem_req_d[41];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__39_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__39_ <= mem_req_d[40];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__38_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__38_ <= mem_req_d[39];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__37_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__37_ <= mem_req_d[38];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__36_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__36_ <= mem_req_d[37];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__35_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__35_ <= mem_req_d[36];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__34_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__34_ <= mem_req_d[35];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__33_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__33_ <= mem_req_d[34];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__32_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__32_ <= mem_req_d[33];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__31_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__31_ <= mem_req_d[32];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__30_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__30_ <= mem_req_d[31];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__29_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__29_ <= mem_req_d[30];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__28_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__28_ <= mem_req_d[29];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__27_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__27_ <= mem_req_d[28];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__26_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__26_ <= mem_req_d[27];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__25_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__25_ <= mem_req_d[26];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__24_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__24_ <= mem_req_d[25];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__23_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__23_ <= mem_req_d[24];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__22_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__22_ <= mem_req_d[23];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__21_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__21_ <= mem_req_d[22];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__20_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__20_ <= mem_req_d[21];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__19_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__19_ <= mem_req_d[20];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__18_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__18_ <= mem_req_d[19];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__17_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__17_ <= mem_req_d[18];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__16_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__16_ <= mem_req_d[17];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__15_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__15_ <= mem_req_d[16];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__14_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__14_ <= mem_req_d[15];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__13_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__13_ <= mem_req_d[14];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__12_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__12_ <= mem_req_d[13];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__11_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__11_ <= mem_req_d[12];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__10_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__10_ <= mem_req_d[11];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__9_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__9_ <= mem_req_d[10];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__8_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__8_ <= mem_req_d[9];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__7_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__7_ <= mem_req_d[8];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__6_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__6_ <= mem_req_d[7];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__5_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__5_ <= mem_req_d[6];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__4_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__4_ <= mem_req_d[5];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__3_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__3_ <= mem_req_d[4];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__2_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__2_ <= mem_req_d[3];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__1_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__1_ <= mem_req_d[2];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_wdata__0_ <= 1'b0;
    end else if(N2186) begin
      mem_req_q_wdata__0_ <= mem_req_d[1];
    end 
  end


  always @(posedge clk_i or posedge N2038) begin
    if(N2038) begin
      mem_req_q_bypass_ <= 1'b0;
    end else if(N2201) begin
      mem_req_q_bypass_ <= mem_req_d[0];
    end 
  end

  assign N2202 = state_q[2] | state_q[3];
  assign N2203 = state_q[1] | N2202;
  assign busy_o = state_q[0] | N2203;
  assign N2205 = ~state_q[2];
  assign N2206 = ~state_q[1];
  assign N2207 = N2205 | state_q[3];
  assign N2208 = N2206 | N2207;
  assign N2209 = state_q[0] | N2208;
  assign N2210 = N2205 | state_q[3];
  assign N2211 = N2206 | N2210;
  assign N2212 = state_q[0] | N2211;
  assign N2213 = ~N2212;
  assign N1557 = ~N1558;
  assign { N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 } = (N0)? data_i[129:2] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N42)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = hit_way_i[0];
  assign { N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172 } = (N1)? data_i[303:176] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N171)? { N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43 } : 1'b0;
  assign N1 = hit_way_i[1];
  assign { N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301 } = (N2)? data_i[477:350] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N300)? { N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172 } : 1'b0;
  assign N2 = hit_way_i[2];
  assign { N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430 } = (N3)? data_i[651:524] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N429)? { N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301 } : 1'b0;
  assign N3 = hit_way_i[3];
  assign { N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559 } = (N4)? data_i[825:698] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N558)? { N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430 } : 1'b0;
  assign N4 = hit_way_i[4];
  assign { N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688 } = (N5)? data_i[999:872] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N687)? { N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559 } : 1'b0;
  assign N5 = hit_way_i[5];
  assign { N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817 } = (N6)? data_i[1173:1046] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N816)? { N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688 } : 1'b0;
  assign N6 = hit_way_i[6];
  assign cl_i = (N7)? data_i[1347:1220] : 
                (N945)? { N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817 } : 1'b0;
  assign N7 = hit_way_i[7];
  assign N990 = ~req_port_i[12];
  assign { N994, N993, N992 } = (N8)? { req_port_i[12:12], N990, req_port_i[12:12] } : 
                                (N2035)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign N8 = bypass_i;
  assign N995 = (N8)? N990 : 
                (N2035)? N991 : 
                (N989)? 1'b0 : 1'b0;
  assign N996 = (N8)? 1'b1 : 
                (N2035)? 1'b0 : 1'b0;
  assign N997 = (N9)? N995 : 
                (N987)? 1'b0 : 1'b0;
  assign N9 = N947;
  assign { N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000 } = (N10)? { mem_req_q_tag__43_, mem_req_q_tag__42_, mem_req_q_tag__41_, mem_req_q_tag__40_, mem_req_q_tag__39_, mem_req_q_tag__38_, mem_req_q_tag__37_, mem_req_q_tag__36_, mem_req_q_tag__35_, mem_req_q_tag__34_, mem_req_q_tag__33_, mem_req_q_tag__32_, mem_req_q_tag__31_, mem_req_q_tag__30_, mem_req_q_tag__29_, mem_req_q_tag__28_, mem_req_q_tag__27_, mem_req_q_tag__26_, mem_req_q_tag__25_, mem_req_q_tag__24_, mem_req_q_tag__23_, mem_req_q_tag__22_, mem_req_q_tag__21_, mem_req_q_tag__20_, mem_req_q_tag__19_, mem_req_q_tag__18_, mem_req_q_tag__17_, mem_req_q_tag__16_, mem_req_q_tag__15_, mem_req_q_tag__14_, mem_req_q_tag__13_, mem_req_q_tag__12_, mem_req_q_tag__11_, mem_req_q_tag__10_, mem_req_q_tag__9_, mem_req_q_tag__8_, mem_req_q_tag__7_, mem_req_q_tag__6_, mem_req_q_tag__5_, mem_req_q_tag__4_, mem_req_q_tag__3_, mem_req_q_tag__2_, mem_req_q_tag__1_, mem_req_q_tag__0_ } : 
                                                                                                                                                                                                                                                                                                                                  (N999)? req_port_i[121:78] : 1'b0;
  assign N10 = N998;
  assign N1048 = (N11)? gnt_i : 
                 (N1047)? 1'b0 : 1'b0;
  assign N11 = N1046;
  assign { N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049 } = (N11)? { req_port_i[121:78], 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                         (N1047)? { mem_req_q_tag__43_, mem_req_q_tag__42_, mem_req_q_tag__41_, mem_req_q_tag__40_, mem_req_q_tag__39_, mem_req_q_tag__38_, mem_req_q_tag__37_, mem_req_q_tag__36_, mem_req_q_tag__35_, mem_req_q_tag__34_, mem_req_q_tag__33_, mem_req_q_tag__32_, mem_req_q_tag__31_, mem_req_q_tag__30_, mem_req_q_tag__29_, mem_req_q_tag__28_, mem_req_q_tag__27_, mem_req_q_tag__26_, mem_req_q_tag__25_, mem_req_q_tag__24_, mem_req_q_tag__23_, mem_req_q_tag__22_, mem_req_q_tag__21_, mem_req_q_tag__20_, mem_req_q_tag__19_, mem_req_q_tag__18_, mem_req_q_tag__17_, mem_req_q_tag__16_, mem_req_q_tag__15_, mem_req_q_tag__14_, mem_req_q_tag__13_, mem_req_q_tag__12_, mem_req_q_tag__11_, mem_req_q_tag__10_, mem_req_q_tag__9_, mem_req_q_tag__8_, mem_req_q_tag__7_, mem_req_q_tag__6_, mem_req_q_tag__5_, mem_req_q_tag__4_, mem_req_q_tag__3_, mem_req_q_tag__2_, mem_req_q_tag__1_, mem_req_q_tag__0_, mem_req_q_bypass_ } : 1'b0;
  assign N1094 = (N11)? gnt_i : 
                 (N1047)? 1'b0 : 1'b0;
  assign { N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095 } = (N12)? cl_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? cl_i[127:64] : 1'b0;
  assign N12 = N1557;
  assign N13 = N1558;
  assign N1159 = (N14)? N1048 : 
                 (N15)? 1'b1 : 1'b0;
  assign N14 = N948;
  assign N15 = mem_req_q_we_;
  assign { N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160 } = (N16)? { N1094, N948, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N1045)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N1044;
  assign N1228 = ~N1044;
  assign { N1227, N1226 } = (N16)? { mem_req_q_we_, N1159 } : 
                            (N1045)? { 1'b0, 1'b1 } : 1'b0;
  assign { N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229 } = (N16)? { N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049 } : 
                                                                                                                                                                                                                                                                                                                                         (N1045)? { req_port_i[121:78], mem_req_q_bypass_ } : 1'b0;
  assign { N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277 } = (N17)? req_port_i[121:78] : 
                                                                                                                                                                                                                                                                                                                                  (N1276)? { N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230 } : 1'b0;
  assign N17 = N2209;
  assign { N1323, N1322, N1321 } = (N18)? { 1'b1, 1'b1, 1'b1 } : 
                                   (N1275)? { N1228, N1227, N1226 } : 1'b0;
  assign N18 = N1274;
  assign { N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324 } = (N18)? { N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277 } : 
                                                                                                                                                                                                                                                                                                                                  (N1275)? { N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230 } : 1'b0;
  assign { N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369 } = (N19)? { req_port_i[121:78], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                         (N20)? { N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1229 } : 1'b0;
  assign N19 = N1368;
  assign N20 = N2247;
  assign { N1416, N1415, N1414 } = (N19)? { 1'b1, 1'b0, 1'b1 } : 
                                   (N20)? { N1323, N1322, N1321 } : 1'b0;
  assign { N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417 } = (N21)? { N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = N949;
  assign N22 = req_port_i[1];
  assign { N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483 } = (N21)? { N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                      (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541 } = (N13)? { mem_req_q_be__7_, mem_req_q_be__6_, mem_req_q_be__5_, mem_req_q_be__4_, mem_req_q_be__3_, mem_req_q_be__2_, mem_req_q_be__1_, mem_req_q_be__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                              (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_req_q_be__7_, mem_req_q_be__6_, mem_req_q_be__5_, mem_req_q_be__4_, mem_req_q_be__3_, mem_req_q_be__2_, mem_req_q_be__1_, mem_req_q_be__0_ } : 
                                                                                                                              (N1540)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561 } = (N13)? { mem_req_q_wdata__63_, mem_req_q_wdata__62_, mem_req_q_wdata__61_, mem_req_q_wdata__60_, mem_req_q_wdata__59_, mem_req_q_wdata__58_, mem_req_q_wdata__57_, mem_req_q_wdata__56_, mem_req_q_wdata__55_, mem_req_q_wdata__54_, mem_req_q_wdata__53_, mem_req_q_wdata__52_, mem_req_q_wdata__51_, mem_req_q_wdata__50_, mem_req_q_wdata__49_, mem_req_q_wdata__48_, mem_req_q_wdata__47_, mem_req_q_wdata__46_, mem_req_q_wdata__45_, mem_req_q_wdata__44_, mem_req_q_wdata__43_, mem_req_q_wdata__42_, mem_req_q_wdata__41_, mem_req_q_wdata__40_, mem_req_q_wdata__39_, mem_req_q_wdata__38_, mem_req_q_wdata__37_, mem_req_q_wdata__36_, mem_req_q_wdata__35_, mem_req_q_wdata__34_, mem_req_q_wdata__33_, mem_req_q_wdata__32_, mem_req_q_wdata__31_, mem_req_q_wdata__30_, mem_req_q_wdata__29_, mem_req_q_wdata__28_, mem_req_q_wdata__27_, mem_req_q_wdata__26_, mem_req_q_wdata__25_, mem_req_q_wdata__24_, mem_req_q_wdata__23_, mem_req_q_wdata__22_, mem_req_q_wdata__21_, mem_req_q_wdata__20_, mem_req_q_wdata__19_, mem_req_q_wdata__18_, mem_req_q_wdata__17_, mem_req_q_wdata__16_, mem_req_q_wdata__15_, mem_req_q_wdata__14_, mem_req_q_wdata__13_, mem_req_q_wdata__12_, mem_req_q_wdata__11_, mem_req_q_wdata__10_, mem_req_q_wdata__9_, mem_req_q_wdata__8_, mem_req_q_wdata__7_, mem_req_q_wdata__6_, mem_req_q_wdata__5_, mem_req_q_wdata__4_, mem_req_q_wdata__3_, mem_req_q_wdata__2_, mem_req_q_wdata__1_, mem_req_q_wdata__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_req_q_wdata__63_, mem_req_q_wdata__62_, mem_req_q_wdata__61_, mem_req_q_wdata__60_, mem_req_q_wdata__59_, mem_req_q_wdata__58_, mem_req_q_wdata__57_, mem_req_q_wdata__56_, mem_req_q_wdata__55_, mem_req_q_wdata__54_, mem_req_q_wdata__53_, mem_req_q_wdata__52_, mem_req_q_wdata__51_, mem_req_q_wdata__50_, mem_req_q_wdata__49_, mem_req_q_wdata__48_, mem_req_q_wdata__47_, mem_req_q_wdata__46_, mem_req_q_wdata__45_, mem_req_q_wdata__44_, mem_req_q_wdata__43_, mem_req_q_wdata__42_, mem_req_q_wdata__41_, mem_req_q_wdata__40_, mem_req_q_wdata__39_, mem_req_q_wdata__38_, mem_req_q_wdata__37_, mem_req_q_wdata__36_, mem_req_q_wdata__35_, mem_req_q_wdata__34_, mem_req_q_wdata__33_, mem_req_q_wdata__32_, mem_req_q_wdata__31_, mem_req_q_wdata__30_, mem_req_q_wdata__29_, mem_req_q_wdata__28_, mem_req_q_wdata__27_, mem_req_q_wdata__26_, mem_req_q_wdata__25_, mem_req_q_wdata__24_, mem_req_q_wdata__23_, mem_req_q_wdata__22_, mem_req_q_wdata__21_, mem_req_q_wdata__20_, mem_req_q_wdata__19_, mem_req_q_wdata__18_, mem_req_q_wdata__17_, mem_req_q_wdata__16_, mem_req_q_wdata__15_, mem_req_q_wdata__14_, mem_req_q_wdata__13_, mem_req_q_wdata__12_, mem_req_q_wdata__11_, mem_req_q_wdata__10_, mem_req_q_wdata__9_, mem_req_q_wdata__8_, mem_req_q_wdata__7_, mem_req_q_wdata__6_, mem_req_q_wdata__5_, mem_req_q_wdata__4_, mem_req_q_wdata__3_, mem_req_q_wdata__2_, mem_req_q_wdata__1_, mem_req_q_wdata__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1560)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689 } = (N23)? hit_way_q : 
                                                                      (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = N950;
  assign N24 = mshr_index_matches_i;
  assign { N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697 } = (N23)? { mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_ } : 
                                                                                                  (N24)? req_port_i[133:122] : 1'b0;
  assign { N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709 } = (N23)? { N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, hit_way_q } : 
                                                                                                                                                                                      (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733 } = (N23)? { N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1861 = (N23)? gnt_i : 
                 (N24)? 1'b0 : 1'b0;
  assign { N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862 } = (N23)? { mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_ } : 
                                                                                                  (N24)? req_port_i[133:122] : 1'b0;
  assign N1875 = (N25)? mem_req_q_we_ : 
                 (N26)? 1'b0 : 1'b0;
  assign N25 = bypass_gnt_i;
  assign N26 = N1874;
  assign { N1880, N1879 } = (N27)? { 1'b1, 1'b0 } : 
                            (N2037)? { 1'b0, 1'b0 } : 
                            (N1878)? { 1'b0, 1'b1 } : 1'b0;
  assign N27 = N1876;
  assign N1881 = (N27)? N1875 : 
                 (N2037)? 1'b1 : 
                 (N1878)? N1875 : 1'b0;
  assign { N1885, N1884 } = (N28)? { 1'b0, 1'b1 } : 
                            (N1883)? { N1880, N1879 } : 1'b0;
  assign N28 = N1882;
  assign N1889 = (N29)? gnt_i : 
                 (N1887)? 1'b0 : 1'b0;
  assign N29 = req_port_i[13];
  assign { N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890 } = (N30)? { N1889, critical_word_i } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N31)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = critical_word_valid_i;
  assign N31 = N1886;
  assign { N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956 } = (N32)? bypass_data_i : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N33)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = bypass_valid_i;
  assign N33 = N1955;
  assign { N2031, N2030, N2029, N2028 } = (N34)? { 1'b0, N994, N993, N992 } : 
                                          (N35)? { 1'b0, N1416, N1415, N1414 } : 
                                          (N36)? { 1'b0, mshr_index_matches_i, mshr_index_matches_i, mshr_index_matches_i } : 
                                          (N37)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                          (N38)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                          (N39)? { N1885, N1884, N1882, N1882 } : 
                                          (N40)? { 1'b0, 1'b0, 1'b0, N1889 } : 
                                          (N41)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N2027)? state_q : 1'b0;
  assign N34 = N955;
  assign N35 = N962;
  assign N36 = N966;
  assign N37 = N970;
  assign N38 = N974;
  assign N39 = N978;
  assign N40 = N982;
  assign N41 = N986;
  assign req_o = (N34)? { N947, N947, N947, N947, N947, N947, N947, N947 } : 
                 (N35)? { N947, N947, N947, N947, N947, N947, N947, N947 } : 
                 (N36)? { N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689 } : 
                 (N37)? { N950, N950, N950, N950, N950, N950, N950, N950 } : 
                 (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N40)? { req_port_i[13:13], req_port_i[13:13], req_port_i[13:13], req_port_i[13:13], req_port_i[13:13], req_port_i[13:13], req_port_i[13:13], req_port_i[13:13] } : 
                 (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N2027)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { mem_req_d[131:120], mem_req_d[75:0] } = (N34)? { req_port_i[133:122], req_port_i[11:2], req_port_i[12:12], req_port_i[77:14], N996 } : 
                                                   (N35)? { req_port_i[133:122], req_port_i[11:2], req_port_i[12:12], req_port_i[77:14], N1369 } : 
                                                   (N40)? { req_port_i[133:122], req_port_i[11:2], req_port_i[12:12], req_port_i[77:14], 1'b0 } : 
                                                   (N2027)? { mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_, mem_req_q_be__7_, mem_req_q_be__6_, mem_req_q_be__5_, mem_req_q_be__4_, mem_req_q_be__3_, mem_req_q_be__2_, mem_req_q_be__1_, mem_req_q_be__0_, mem_req_q_size__1_, mem_req_q_size__0_, mem_req_q_we_, mem_req_q_wdata__63_, mem_req_q_wdata__62_, mem_req_q_wdata__61_, mem_req_q_wdata__60_, mem_req_q_wdata__59_, mem_req_q_wdata__58_, mem_req_q_wdata__57_, mem_req_q_wdata__56_, mem_req_q_wdata__55_, mem_req_q_wdata__54_, mem_req_q_wdata__53_, mem_req_q_wdata__52_, mem_req_q_wdata__51_, mem_req_q_wdata__50_, mem_req_q_wdata__49_, mem_req_q_wdata__48_, mem_req_q_wdata__47_, mem_req_q_wdata__46_, mem_req_q_wdata__45_, mem_req_q_wdata__44_, mem_req_q_wdata__43_, mem_req_q_wdata__42_, mem_req_q_wdata__41_, mem_req_q_wdata__40_, mem_req_q_wdata__39_, mem_req_q_wdata__38_, mem_req_q_wdata__37_, mem_req_q_wdata__36_, mem_req_q_wdata__35_, mem_req_q_wdata__34_, mem_req_q_wdata__33_, mem_req_q_wdata__32_, mem_req_q_wdata__31_, mem_req_q_wdata__30_, mem_req_q_wdata__29_, mem_req_q_wdata__28_, mem_req_q_wdata__27_, mem_req_q_wdata__26_, mem_req_q_wdata__25_, mem_req_q_wdata__24_, mem_req_q_wdata__23_, mem_req_q_wdata__22_, mem_req_q_wdata__21_, mem_req_q_wdata__20_, mem_req_q_wdata__19_, mem_req_q_wdata__18_, mem_req_q_wdata__17_, mem_req_q_wdata__16_, mem_req_q_wdata__15_, mem_req_q_wdata__14_, mem_req_q_wdata__13_, mem_req_q_wdata__12_, mem_req_q_wdata__11_, mem_req_q_wdata__10_, mem_req_q_wdata__9_, mem_req_q_wdata__8_, mem_req_q_wdata__7_, mem_req_q_wdata__6_, mem_req_q_wdata__5_, mem_req_q_wdata__4_, mem_req_q_wdata__3_, mem_req_q_wdata__2_, mem_req_q_wdata__1_, mem_req_q_wdata__0_, mem_req_q_bypass_ } : 1'b0;
  assign mem_req_d[119:76] = (N34)? req_port_i[121:78] : 
                             (N35)? { N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370 } : 
                             (N38)? req_port_i[121:78] : 
                             (N40)? req_port_i[121:78] : 
                             (N2027)? { mem_req_q_tag__43_, mem_req_q_tag__42_, mem_req_q_tag__41_, mem_req_q_tag__40_, mem_req_q_tag__39_, mem_req_q_tag__38_, mem_req_q_tag__37_, mem_req_q_tag__36_, mem_req_q_tag__35_, mem_req_q_tag__34_, mem_req_q_tag__33_, mem_req_q_tag__32_, mem_req_q_tag__31_, mem_req_q_tag__30_, mem_req_q_tag__29_, mem_req_q_tag__28_, mem_req_q_tag__27_, mem_req_q_tag__26_, mem_req_q_tag__25_, mem_req_q_tag__24_, mem_req_q_tag__23_, mem_req_q_tag__22_, mem_req_q_tag__21_, mem_req_q_tag__20_, mem_req_q_tag__19_, mem_req_q_tag__18_, mem_req_q_tag__17_, mem_req_q_tag__16_, mem_req_q_tag__15_, mem_req_q_tag__14_, mem_req_q_tag__13_, mem_req_q_tag__12_, mem_req_q_tag__11_, mem_req_q_tag__10_, mem_req_q_tag__9_, mem_req_q_tag__8_, mem_req_q_tag__7_, mem_req_q_tag__6_, mem_req_q_tag__5_, mem_req_q_tag__4_, mem_req_q_tag__3_, mem_req_q_tag__2_, mem_req_q_tag__1_, mem_req_q_tag__0_ } : 1'b0;
  assign { req_port_o[65:65], N2032, req_port_o[63:0] } = (N34)? { N997, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                          (N35)? { N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417 } : 
                                                          (N36)? { N1861, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                          (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                          (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                          (N39)? { N1881, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                          (N40)? { N1954, critical_word_valid_i, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890 } : 
                                                          (N41)? { 1'b0, bypass_valid_i, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956 } : 
                                                          (N2027)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_o = (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N35)? { N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000 } : 
                 (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N2027)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign mshr_addr_o = (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N35)? { N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483 } : 
                       (N36)? { mem_req_q_tag__43_, mem_req_q_tag__42_, mem_req_q_tag__41_, mem_req_q_tag__40_, mem_req_q_tag__39_, mem_req_q_tag__38_, mem_req_q_tag__37_, mem_req_q_tag__36_, mem_req_q_tag__35_, mem_req_q_tag__34_, mem_req_q_tag__33_, mem_req_q_tag__32_, mem_req_q_tag__31_, mem_req_q_tag__30_, mem_req_q_tag__29_, mem_req_q_tag__28_, mem_req_q_tag__27_, mem_req_q_tag__26_, mem_req_q_tag__25_, mem_req_q_tag__24_, mem_req_q_tag__23_, mem_req_q_tag__22_, mem_req_q_tag__21_, mem_req_q_tag__20_, mem_req_q_tag__19_, mem_req_q_tag__18_, mem_req_q_tag__17_, mem_req_q_tag__16_, mem_req_q_tag__15_, mem_req_q_tag__14_, mem_req_q_tag__13_, mem_req_q_tag__12_, mem_req_q_tag__11_, mem_req_q_tag__10_, mem_req_q_tag__9_, mem_req_q_tag__8_, mem_req_q_tag__7_, mem_req_q_tag__6_, mem_req_q_tag__5_, mem_req_q_tag__4_, mem_req_q_tag__3_, mem_req_q_tag__2_, mem_req_q_tag__1_, mem_req_q_tag__0_, mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_ } : 
                       (N37)? { mem_req_q_tag__43_, mem_req_q_tag__42_, mem_req_q_tag__41_, mem_req_q_tag__40_, mem_req_q_tag__39_, mem_req_q_tag__38_, mem_req_q_tag__37_, mem_req_q_tag__36_, mem_req_q_tag__35_, mem_req_q_tag__34_, mem_req_q_tag__33_, mem_req_q_tag__32_, mem_req_q_tag__31_, mem_req_q_tag__30_, mem_req_q_tag__29_, mem_req_q_tag__28_, mem_req_q_tag__27_, mem_req_q_tag__26_, mem_req_q_tag__25_, mem_req_q_tag__24_, mem_req_q_tag__23_, mem_req_q_tag__22_, mem_req_q_tag__21_, mem_req_q_tag__20_, mem_req_q_tag__19_, mem_req_q_tag__18_, mem_req_q_tag__17_, mem_req_q_tag__16_, mem_req_q_tag__15_, mem_req_q_tag__14_, mem_req_q_tag__13_, mem_req_q_tag__12_, mem_req_q_tag__11_, mem_req_q_tag__10_, mem_req_q_tag__9_, mem_req_q_tag__8_, mem_req_q_tag__7_, mem_req_q_tag__6_, mem_req_q_tag__5_, mem_req_q_tag__4_, mem_req_q_tag__3_, mem_req_q_tag__2_, mem_req_q_tag__1_, mem_req_q_tag__0_, mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_ } : 
                       (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N39)? { mem_req_q_tag__43_, mem_req_q_tag__42_, mem_req_q_tag__41_, mem_req_q_tag__40_, mem_req_q_tag__39_, mem_req_q_tag__38_, mem_req_q_tag__37_, mem_req_q_tag__36_, mem_req_q_tag__35_, mem_req_q_tag__34_, mem_req_q_tag__33_, mem_req_q_tag__32_, mem_req_q_tag__31_, mem_req_q_tag__30_, mem_req_q_tag__29_, mem_req_q_tag__28_, mem_req_q_tag__27_, mem_req_q_tag__26_, mem_req_q_tag__25_, mem_req_q_tag__24_, mem_req_q_tag__23_, mem_req_q_tag__22_, mem_req_q_tag__21_, mem_req_q_tag__20_, mem_req_q_tag__19_, mem_req_q_tag__18_, mem_req_q_tag__17_, mem_req_q_tag__16_, mem_req_q_tag__15_, mem_req_q_tag__14_, mem_req_q_tag__13_, mem_req_q_tag__12_, mem_req_q_tag__11_, mem_req_q_tag__10_, mem_req_q_tag__9_, mem_req_q_tag__8_, mem_req_q_tag__7_, mem_req_q_tag__6_, mem_req_q_tag__5_, mem_req_q_tag__4_, mem_req_q_tag__3_, mem_req_q_tag__2_, mem_req_q_tag__1_, mem_req_q_tag__0_, mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_ } : 
                       (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N2027)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign hit_way_d = (N35)? hit_way_i : 
                     (N2027)? hit_way_q : 1'b0;
  assign addr_o = (N34)? req_port_i[133:122] : 
                  (N35)? req_port_i[133:122] : 
                  (N36)? { N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697 } : 
                  (N37)? { N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862 } : 
                  (N38)? req_port_i[133:122] : 
                  (N39)? req_port_i[133:122] : 
                  (N40)? req_port_i[133:122] : 
                  (N41)? req_port_i[133:122] : 
                  (N2027)? req_port_i[133:122] : 1'b0;
  assign we_o = (N34)? 1'b0 : 
                (N35)? 1'b0 : 
                (N36)? N950 : 
                (N37)? 1'b0 : 
                (N38)? 1'b0 : 
                (N39)? 1'b0 : 
                (N40)? 1'b0 : 
                (N41)? 1'b0 : 
                (N2027)? 1'b0 : 1'b0;
  assign be_o[23:0] = (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N36)? { N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709 } : 
                      (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                      (N2027)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_o[129:0] = (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N36)? { N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N950, N950 } : 
                         (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N39)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N2027)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { miss_req_o[140:140], miss_req_o[131:0] } = (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N39)? { 1'b1, mem_req_q_tag__43_, mem_req_q_tag__42_, mem_req_q_tag__41_, mem_req_q_tag__40_, mem_req_q_tag__39_, mem_req_q_tag__38_, mem_req_q_tag__37_, mem_req_q_tag__36_, mem_req_q_tag__35_, mem_req_q_tag__34_, mem_req_q_tag__33_, mem_req_q_tag__32_, mem_req_q_tag__31_, mem_req_q_tag__30_, mem_req_q_tag__29_, mem_req_q_tag__28_, mem_req_q_tag__27_, mem_req_q_tag__26_, mem_req_q_tag__25_, mem_req_q_tag__24_, mem_req_q_tag__23_, mem_req_q_tag__22_, mem_req_q_tag__21_, mem_req_q_tag__20_, mem_req_q_tag__19_, mem_req_q_tag__18_, mem_req_q_tag__17_, mem_req_q_tag__16_, mem_req_q_tag__15_, mem_req_q_tag__14_, mem_req_q_tag__13_, mem_req_q_tag__12_, mem_req_q_tag__11_, mem_req_q_tag__10_, mem_req_q_tag__9_, mem_req_q_tag__8_, mem_req_q_tag__7_, mem_req_q_tag__6_, mem_req_q_tag__5_, mem_req_q_tag__4_, mem_req_q_tag__3_, mem_req_q_tag__2_, mem_req_q_tag__1_, mem_req_q_tag__0_, mem_req_q_index__11_, mem_req_q_index__10_, mem_req_q_index__9_, mem_req_q_index__8_, mem_req_q_index__7_, mem_req_q_index__6_, mem_req_q_index__5_, mem_req_q_index__4_, N1558, mem_req_q_index__2_, mem_req_q_index__1_, mem_req_q_index__0_, mem_req_q_be__7_, mem_req_q_be__6_, mem_req_q_be__5_, mem_req_q_be__4_, mem_req_q_be__3_, mem_req_q_be__2_, mem_req_q_be__1_, mem_req_q_be__0_, mem_req_q_size__1_, mem_req_q_size__0_, mem_req_q_we_, mem_req_q_wdata__63_, mem_req_q_wdata__62_, mem_req_q_wdata__61_, mem_req_q_wdata__60_, mem_req_q_wdata__59_, mem_req_q_wdata__58_, mem_req_q_wdata__57_, mem_req_q_wdata__56_, mem_req_q_wdata__55_, mem_req_q_wdata__54_, mem_req_q_wdata__53_, mem_req_q_wdata__52_, mem_req_q_wdata__51_, mem_req_q_wdata__50_, mem_req_q_wdata__49_, mem_req_q_wdata__48_, mem_req_q_wdata__47_, mem_req_q_wdata__46_, mem_req_q_wdata__45_, mem_req_q_wdata__44_, mem_req_q_wdata__43_, mem_req_q_wdata__42_, mem_req_q_wdata__41_, mem_req_q_wdata__40_, mem_req_q_wdata__39_, mem_req_q_wdata__38_, mem_req_q_wdata__37_, mem_req_q_wdata__36_, mem_req_q_wdata__35_, mem_req_q_wdata__34_, mem_req_q_wdata__33_, mem_req_q_wdata__32_, mem_req_q_wdata__31_, mem_req_q_wdata__30_, mem_req_q_wdata__29_, mem_req_q_wdata__28_, mem_req_q_wdata__27_, mem_req_q_wdata__26_, mem_req_q_wdata__25_, mem_req_q_wdata__24_, mem_req_q_wdata__23_, mem_req_q_wdata__22_, mem_req_q_wdata__21_, mem_req_q_wdata__20_, mem_req_q_wdata__19_, mem_req_q_wdata__18_, mem_req_q_wdata__17_, mem_req_q_wdata__16_, mem_req_q_wdata__15_, mem_req_q_wdata__14_, mem_req_q_wdata__13_, mem_req_q_wdata__12_, mem_req_q_wdata__11_, mem_req_q_wdata__10_, mem_req_q_wdata__9_, mem_req_q_wdata__8_, mem_req_q_wdata__7_, mem_req_q_wdata__6_, mem_req_q_wdata__5_, mem_req_q_wdata__4_, mem_req_q_wdata__3_, mem_req_q_wdata__2_, mem_req_q_wdata__1_, mem_req_q_wdata__0_, mem_req_q_bypass_ } : 
                                                      (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N2027)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign state_d = (N22)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                   (N2033)? { N2031, N2030, N2029, N2028 } : 1'b0;
  assign req_port_o[64] = (N22)? 1'b1 : 
                          (N2033)? N2032 : 1'b0;
  assign N42 = ~hit_way_i[0];
  assign N171 = ~hit_way_i[1];
  assign N300 = ~hit_way_i[2];
  assign N429 = ~hit_way_i[3];
  assign N558 = ~hit_way_i[4];
  assign N687 = ~hit_way_i[5];
  assign N816 = ~hit_way_i[6];
  assign N945 = ~hit_way_i[7];
  assign N946 = ~flush_i;
  assign N947 = req_port_i[13] & N946;
  assign N948 = ~mem_req_q_we_;
  assign N949 = ~req_port_i[1];
  assign N950 = ~mshr_index_matches_i;
  assign N951 = ~state_q[3];
  assign N952 = ~state_q[0];
  assign N962 = N2214 | N2215;
  assign N2214 = ~N958;
  assign N2215 = ~N961;
  assign N966 = ~N965;
  assign N970 = ~N969;
  assign N974 = ~N973;
  assign N978 = ~N977;
  assign N982 = ~N981;
  assign N986 = ~N985;
  assign N987 = ~N947;
  assign N988 = gnt_i | bypass_i;
  assign N989 = ~N988;
  assign N991 = ~req_port_i[12];
  assign N998 = N2213 | mem_req_q_we_;
  assign N999 = ~N998;
  assign N1044 = N2221 | hit_way_i[0];
  assign N2221 = N2220 | hit_way_i[1];
  assign N2220 = N2219 | hit_way_i[2];
  assign N2219 = N2218 | hit_way_i[3];
  assign N2218 = N2217 | hit_way_i[4];
  assign N2217 = N2216 | hit_way_i[5];
  assign N2216 = hit_way_i[7] | hit_way_i[6];
  assign N1045 = ~N1044;
  assign N1046 = N2222 & N946;
  assign N2222 = req_port_i[13] & N948;
  assign N1047 = ~N1046;
  assign N1274 = N2223 | mshr_addr_matches_i;
  assign N2223 = mshr_index_matches_i & mem_req_q_we_;
  assign N1275 = ~N1274;
  assign N1276 = ~N2209;
  assign N1368 = ~N2247;
  assign N2247 = N2246 | N1019;
  assign N2246 = N2245 | N1020;
  assign N2245 = N2244 | N1021;
  assign N2244 = N2243 | N1022;
  assign N2243 = N2242 | N1023;
  assign N2242 = N2241 | N1024;
  assign N2241 = N2240 | N1025;
  assign N2240 = N2239 | N1026;
  assign N2239 = N2238 | N1027;
  assign N2238 = N2237 | N1028;
  assign N2237 = N2236 | N1029;
  assign N2236 = N2235 | N1030;
  assign N2235 = N2234 | N1031;
  assign N2234 = N2233 | N1032;
  assign N2233 = N2232 | N1033;
  assign N2232 = N2231 | N1034;
  assign N2231 = N2230 | N1035;
  assign N2230 = N2229 | N1036;
  assign N2229 = N2228 | N1037;
  assign N2228 = N2227 | N1038;
  assign N2227 = N2226 | N1039;
  assign N2226 = N2225 | N1040;
  assign N2225 = N2224 | N1041;
  assign N2224 = N1043 | N1042;
  assign N1539 = N1557 | N1558;
  assign N1540 = ~N1539;
  assign N1559 = N1557 | N1558;
  assign N1560 = ~N1559;
  assign N1874 = ~bypass_gnt_i;
  assign N1876 = miss_gnt_i & N948;
  assign N1877 = miss_gnt_i | N1876;
  assign N1878 = ~N1877;
  assign N1882 = mshr_addr_matches_i & N2248;
  assign N2248 = ~active_serving_i;
  assign N1883 = ~N1882;
  assign N1886 = ~critical_word_valid_i;
  assign N1887 = ~req_port_i[13];
  assign N1888 = ~gnt_i;
  assign N1955 = ~bypass_valid_i;
  assign N2020 = N962 | N955;
  assign N2021 = N966 | N2020;
  assign N2022 = N970 | N2021;
  assign N2023 = N974 | N2022;
  assign N2024 = N978 | N2023;
  assign N2025 = N982 | N2024;
  assign N2026 = N986 | N2025;
  assign N2027 = ~N2026;
  assign N2033 = ~req_port_i[1];
  assign N2034 = ~bypass_i;
  assign N2035 = gnt_i & N2034;
  assign N2036 = ~N1876;
  assign N2037 = miss_gnt_i & N2036;
  assign N2038 = ~rst_ni;
  assign N2039 = N949 & N962;
  assign N2040 = N1044 & N2039;
  assign N2041 = N948 & N2040;
  assign N2042 = N955 | N2041;
  assign N2043 = N949 & N962;
  assign N2044 = N1045 & N2043;
  assign N2045 = N2042 | N2044;
  assign N2046 = req_port_i[1] & N962;
  assign N2047 = N2045 | N2046;
  assign N2048 = N2047 | N966;
  assign N2049 = N2048 | N970;
  assign N2050 = N2049 | N974;
  assign N2051 = N2050 | N978;
  assign N2052 = N2051 | N982;
  assign N2053 = N2052 | N986;
  assign N2054 = ~N2053;
  assign N2055 = N1044 & N2043;
  assign N2056 = N948 & N2055;
  assign N2057 = N955 | N2056;
  assign N2058 = N2057 | N2044;
  assign N2059 = req_port_i[1] & N962;
  assign N2060 = N2058 | N2059;
  assign N2061 = N2060 | N966;
  assign N2062 = N2061 | N970;
  assign N2063 = N2062 | N974;
  assign N2064 = N2063 | N978;
  assign N2065 = N2064 | N982;
  assign N2066 = N2065 | N986;
  assign N2067 = ~N2066;
  assign N2068 = N955 & N2033;
  assign N2069 = N947 & N2068;
  assign N2070 = N989 & N2069;
  assign N2071 = N987 & N2068;
  assign N2072 = N2070 | N2071;
  assign N2073 = N962 & N2033;
  assign N2074 = req_port_i[1] & N2073;
  assign N2075 = N2072 | N2074;
  assign N2076 = N966 & N2033;
  assign N2077 = N950 & N2076;
  assign N2078 = N1888 & N2077;
  assign N2079 = N2075 | N2078;
  assign N2080 = N970 & N2033;
  assign N2081 = N950 & N2080;
  assign N2082 = N1888 & N2081;
  assign N2083 = N2079 | N2082;
  assign N2084 = mshr_index_matches_i & N2080;
  assign N2085 = N2083 | N2084;
  assign N2086 = N974 & N2033;
  assign N2087 = req_port_i[1] & N2086;
  assign N2088 = N2085 | N2087;
  assign N2089 = N978 & N2033;
  assign N2090 = N1883 & N2089;
  assign N2091 = N1878 & N2090;
  assign N2092 = N1874 & N2091;
  assign N2093 = N2088 | N2092;
  assign N2094 = N982 & N2033;
  assign N2095 = N1886 & N2094;
  assign N2096 = N2093 | N2095;
  assign N2097 = N986 & N2033;
  assign N2098 = N1955 & N2097;
  assign N2099 = N2096 | N2098;
  assign N2100 = ~N2099;
  assign N2101 = N987 & N955;
  assign N2102 = N1047 & N2055;
  assign N2103 = N2101 | N2102;
  assign N2104 = N2103 | N2044;
  assign N2105 = N2104 | N2059;
  assign N2106 = N2105 | N966;
  assign N2107 = N2106 | N970;
  assign N2108 = N2107 | N974;
  assign N2109 = N2108 | N978;
  assign N2110 = critical_word_valid_i & N982;
  assign N2111 = N1887 & N2110;
  assign N2112 = N2109 | N2111;
  assign N2113 = N1886 & N982;
  assign N2114 = N2112 | N2113;
  assign N2115 = N2114 | N986;
  assign N2116 = ~N2115;
  assign N2117 = N987 & N955;
  assign N2118 = N2117 | N2102;
  assign N2119 = N2118 | N2044;
  assign N2120 = N2119 | N2059;
  assign N2121 = N2120 | N966;
  assign N2122 = N2121 | N970;
  assign N2123 = N2122 | N974;
  assign N2124 = N2123 | N978;
  assign N2125 = critical_word_valid_i & N982;
  assign N2126 = N1887 & N2125;
  assign N2127 = N2124 | N2126;
  assign N2128 = N1886 & N982;
  assign N2129 = N2127 | N2128;
  assign N2130 = N2129 | N986;
  assign N2131 = ~N2130;
  assign N2132 = N2117 | N2059;
  assign N2133 = N2132 | N966;
  assign N2134 = N2133 | N970;
  assign N2135 = req_port_i[1] & N974;
  assign N2136 = N2134 | N2135;
  assign N2137 = N2136 | N978;
  assign N2138 = N2137 | N2126;
  assign N2139 = N2138 | N2128;
  assign N2140 = N2139 | N986;
  assign N2141 = ~N2140;
  assign N2142 = N2101 | N2046;
  assign N2143 = N2142 | N966;
  assign N2144 = N2143 | N970;
  assign N2145 = N2144 | N2135;
  assign N2146 = N2145 | N978;
  assign N2147 = N2146 | N2126;
  assign N2148 = N2147 | N2113;
  assign N2149 = N2148 | N986;
  assign N2150 = ~N2149;
  assign N2151 = N2146 | N2111;
  assign N2152 = N2151 | N2113;
  assign N2153 = N2152 | N986;
  assign N2154 = ~N2153;
  assign N2155 = N2104 | N2046;
  assign N2156 = N2155 | N966;
  assign N2157 = N2156 | N970;
  assign N2158 = N2157 | N974;
  assign N2159 = N2158 | N978;
  assign N2160 = N2159 | N2111;
  assign N2161 = N2160 | N2113;
  assign N2162 = N2161 | N986;
  assign N2163 = ~N2162;
  assign N2164 = N1045 & N2039;
  assign N2165 = N2103 | N2164;
  assign N2166 = N2165 | N2046;
  assign N2167 = N2166 | N966;
  assign N2168 = N2167 | N970;
  assign N2169 = N2168 | N974;
  assign N2170 = N2169 | N978;
  assign N2171 = N2170 | N2111;
  assign N2172 = N2171 | N2113;
  assign N2173 = N2172 | N986;
  assign N2174 = ~N2173;
  assign N2175 = N1047 & N2040;
  assign N2176 = N2101 | N2175;
  assign N2177 = N2176 | N2164;
  assign N2178 = N2177 | N2046;
  assign N2179 = N2178 | N966;
  assign N2180 = N2179 | N970;
  assign N2181 = N2180 | N974;
  assign N2182 = N2181 | N978;
  assign N2183 = N2182 | N2111;
  assign N2184 = N2183 | N2113;
  assign N2185 = N2184 | N986;
  assign N2186 = ~N2185;
  assign N2187 = N947 & N955;
  assign N2188 = N989 & N2187;
  assign N2189 = N2188 | N2101;
  assign N2190 = N2189 | N2046;
  assign N2191 = N2190 | N966;
  assign N2192 = N2191 | N970;
  assign N2193 = N2192 | N974;
  assign N2194 = N2193 | N978;
  assign N2195 = req_port_i[13] & N2110;
  assign N2196 = N1888 & N2195;
  assign N2197 = N2194 | N2196;
  assign N2198 = N2197 | N2111;
  assign N2199 = N2198 | N2113;
  assign N2200 = N2199 | N986;
  assign N2201 = ~N2200;

endmodule