module rvtwoscomp_WIDTH32
(
  din,
  dout
);

  input [31:0] din;
  output [31:0] dout;
  wire [31:0] dout;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557;
  assign dout[0] = din[0];
  assign dout[1] = (N0)? N32 :
                   (N31)? din[1] : 1'b0;
  assign N0 = din[0];
  assign dout[2] = (N1)? N35 :
                   (N34)? din[2] : 1'b0;
  assign N1 = N33;
  assign dout[3] = (N2)? N38 :
                   (N37)? din[3] : 1'b0;
  assign N2 = N36;
  assign dout[4] = (N3)? N41 :
                   (N40)? din[4] : 1'b0;
  assign N3 = N39;
  assign dout[5] = (N4)? N44 :
                   (N43)? din[5] : 1'b0;
  assign N4 = N42;
  assign dout[6] = (N5)? N47 :
                   (N46)? din[6] : 1'b0;
  assign N5 = N45;
  assign dout[7] = (N6)? N50 :
                   (N49)? din[7] : 1'b0;
  assign N6 = N48;
  assign dout[8] = (N7)? N53 :
                   (N52)? din[8] : 1'b0;
  assign N7 = N51;
  assign dout[9] = (N8)? N56 :
                   (N55)? din[9] : 1'b0;
  assign N8 = N54;
  assign dout[10] = (N9)? N59 :
                    (N58)? din[10] : 1'b0;
  assign N9 = N57;
  assign dout[11] = (N10)? N62 :
                    (N61)? din[11] : 1'b0;
  assign N10 = N60;
  assign dout[12] = (N11)? N65 :
                    (N64)? din[12] : 1'b0;
  assign N11 = N63;
  assign dout[13] = (N12)? N68 :
                    (N67)? din[13] : 1'b0;
  assign N12 = N66;
  assign dout[14] = (N13)? N71 :
                    (N70)? din[14] : 1'b0;
  assign N13 = N69;
  assign dout[15] = (N14)? N74 :
                    (N73)? din[15] : 1'b0;
  assign N14 = N72;
  assign dout[16] = (N15)? N77 :
                    (N76)? din[16] : 1'b0;
  assign N15 = N75;
  assign dout[17] = (N16)? N80 :
                    (N79)? din[17] : 1'b0;
  assign N16 = N78;
  assign dout[18] = (N17)? N83 :
                    (N82)? din[18] : 1'b0;
  assign N17 = N81;
  assign dout[19] = (N18)? N86 :
                    (N85)? din[19] : 1'b0;
  assign N18 = N84;
  assign dout[20] = (N19)? N89 :
                    (N88)? din[20] : 1'b0;
  assign N19 = N87;
  assign dout[21] = (N20)? N92 :
                    (N91)? din[21] : 1'b0;
  assign N20 = N90;
  assign dout[22] = (N21)? N95 :
                    (N94)? din[22] : 1'b0;
  assign N21 = N93;
  assign dout[23] = (N22)? N98 :
                    (N97)? din[23] : 1'b0;
  assign N22 = N96;
  assign dout[24] = (N23)? N101 :
                    (N100)? din[24] : 1'b0;
  assign N23 = N99;
  assign dout[25] = (N24)? N104 :
                    (N103)? din[25] : 1'b0;
  assign N24 = N102;
  assign dout[26] = (N25)? N107 :
                    (N106)? din[26] : 1'b0;
  assign N25 = N105;
  assign dout[27] = (N26)? N110 :
                    (N109)? din[27] : 1'b0;
  assign N26 = N108;
  assign dout[28] = (N27)? N113 :
                    (N112)? din[28] : 1'b0;
  assign N27 = N111;
  assign dout[29] = (N28)? N116 :
                    (N115)? din[29] : 1'b0;
  assign N28 = N114;
  assign dout[30] = (N29)? N119 :
                    (N118)? din[30] : 1'b0;
  assign N29 = N117;
  assign dout[31] = (N30)? N122 :
                    (N121)? din[31] : 1'b0;
  assign N30 = N120;
  assign N31 = ~din[0];
  assign N32 = ~din[1];
  assign N33 = din[1] | din[0];
  assign N34 = ~N33;
  assign N35 = ~din[2];
  assign N36 = N123 | din[0];
  assign N123 = din[2] | din[1];
  assign N37 = ~N36;
  assign N38 = ~din[3];
  assign N39 = N125 | din[0];
  assign N125 = N124 | din[1];
  assign N124 = din[3] | din[2];
  assign N40 = ~N39;
  assign N41 = ~din[4];
  assign N42 = N128 | din[0];
  assign N128 = N127 | din[1];
  assign N127 = N126 | din[2];
  assign N126 = din[4] | din[3];
  assign N43 = ~N42;
  assign N44 = ~din[5];
  assign N45 = N132 | din[0];
  assign N132 = N131 | din[1];
  assign N131 = N130 | din[2];
  assign N130 = N129 | din[3];
  assign N129 = din[5] | din[4];
  assign N46 = ~N45;
  assign N47 = ~din[6];
  assign N48 = N137 | din[0];
  assign N137 = N136 | din[1];
  assign N136 = N135 | din[2];
  assign N135 = N134 | din[3];
  assign N134 = N133 | din[4];
  assign N133 = din[6] | din[5];
  assign N49 = ~N48;
  assign N50 = ~din[7];
  assign N51 = N143 | din[0];
  assign N143 = N142 | din[1];
  assign N142 = N141 | din[2];
  assign N141 = N140 | din[3];
  assign N140 = N139 | din[4];
  assign N139 = N138 | din[5];
  assign N138 = din[7] | din[6];
  assign N52 = ~N51;
  assign N53 = ~din[8];
  assign N54 = N150 | din[0];
  assign N150 = N149 | din[1];
  assign N149 = N148 | din[2];
  assign N148 = N147 | din[3];
  assign N147 = N146 | din[4];
  assign N146 = N145 | din[5];
  assign N145 = N144 | din[6];
  assign N144 = din[8] | din[7];
  assign N55 = ~N54;
  assign N56 = ~din[9];
  assign N57 = N158 | din[0];
  assign N158 = N157 | din[1];
  assign N157 = N156 | din[2];
  assign N156 = N155 | din[3];
  assign N155 = N154 | din[4];
  assign N154 = N153 | din[5];
  assign N153 = N152 | din[6];
  assign N152 = N151 | din[7];
  assign N151 = din[9] | din[8];
  assign N58 = ~N57;
  assign N59 = ~din[10];
  assign N60 = N167 | din[0];
  assign N167 = N166 | din[1];
  assign N166 = N165 | din[2];
  assign N165 = N164 | din[3];
  assign N164 = N163 | din[4];
  assign N163 = N162 | din[5];
  assign N162 = N161 | din[6];
  assign N161 = N160 | din[7];
  assign N160 = N159 | din[8];
  assign N159 = din[10] | din[9];
  assign N61 = ~N60;
  assign N62 = ~din[11];
  assign N63 = N177 | din[0];
  assign N177 = N176 | din[1];
  assign N176 = N175 | din[2];
  assign N175 = N174 | din[3];
  assign N174 = N173 | din[4];
  assign N173 = N172 | din[5];
  assign N172 = N171 | din[6];
  assign N171 = N170 | din[7];
  assign N170 = N169 | din[8];
  assign N169 = N168 | din[9];
  assign N168 = din[11] | din[10];
  assign N64 = ~N63;
  assign N65 = ~din[12];
  assign N66 = N188 | din[0];
  assign N188 = N187 | din[1];
  assign N187 = N186 | din[2];
  assign N186 = N185 | din[3];
  assign N185 = N184 | din[4];
  assign N184 = N183 | din[5];
  assign N183 = N182 | din[6];
  assign N182 = N181 | din[7];
  assign N181 = N180 | din[8];
  assign N180 = N179 | din[9];
  assign N179 = N178 | din[10];
  assign N178 = din[12] | din[11];
  assign N67 = ~N66;
  assign N68 = ~din[13];
  assign N69 = N200 | din[0];
  assign N200 = N199 | din[1];
  assign N199 = N198 | din[2];
  assign N198 = N197 | din[3];
  assign N197 = N196 | din[4];
  assign N196 = N195 | din[5];
  assign N195 = N194 | din[6];
  assign N194 = N193 | din[7];
  assign N193 = N192 | din[8];
  assign N192 = N191 | din[9];
  assign N191 = N190 | din[10];
  assign N190 = N189 | din[11];
  assign N189 = din[13] | din[12];
  assign N70 = ~N69;
  assign N71 = ~din[14];
  assign N72 = N213 | din[0];
  assign N213 = N212 | din[1];
  assign N212 = N211 | din[2];
  assign N211 = N210 | din[3];
  assign N210 = N209 | din[4];
  assign N209 = N208 | din[5];
  assign N208 = N207 | din[6];
  assign N207 = N206 | din[7];
  assign N206 = N205 | din[8];
  assign N205 = N204 | din[9];
  assign N204 = N203 | din[10];
  assign N203 = N202 | din[11];
  assign N202 = N201 | din[12];
  assign N201 = din[14] | din[13];
  assign N73 = ~N72;
  assign N74 = ~din[15];
  assign N75 = N227 | din[0];
  assign N227 = N226 | din[1];
  assign N226 = N225 | din[2];
  assign N225 = N224 | din[3];
  assign N224 = N223 | din[4];
  assign N223 = N222 | din[5];
  assign N222 = N221 | din[6];
  assign N221 = N220 | din[7];
  assign N220 = N219 | din[8];
  assign N219 = N218 | din[9];
  assign N218 = N217 | din[10];
  assign N217 = N216 | din[11];
  assign N216 = N215 | din[12];
  assign N215 = N214 | din[13];
  assign N214 = din[15] | din[14];
  assign N76 = ~N75;
  assign N77 = ~din[16];
  assign N78 = N242 | din[0];
  assign N242 = N241 | din[1];
  assign N241 = N240 | din[2];
  assign N240 = N239 | din[3];
  assign N239 = N238 | din[4];
  assign N238 = N237 | din[5];
  assign N237 = N236 | din[6];
  assign N236 = N235 | din[7];
  assign N235 = N234 | din[8];
  assign N234 = N233 | din[9];
  assign N233 = N232 | din[10];
  assign N232 = N231 | din[11];
  assign N231 = N230 | din[12];
  assign N230 = N229 | din[13];
  assign N229 = N228 | din[14];
  assign N228 = din[16] | din[15];
  assign N79 = ~N78;
  assign N80 = ~din[17];
  assign N81 = N258 | din[0];
  assign N258 = N257 | din[1];
  assign N257 = N256 | din[2];
  assign N256 = N255 | din[3];
  assign N255 = N254 | din[4];
  assign N254 = N253 | din[5];
  assign N253 = N252 | din[6];
  assign N252 = N251 | din[7];
  assign N251 = N250 | din[8];
  assign N250 = N249 | din[9];
  assign N249 = N248 | din[10];
  assign N248 = N247 | din[11];
  assign N247 = N246 | din[12];
  assign N246 = N245 | din[13];
  assign N245 = N244 | din[14];
  assign N244 = N243 | din[15];
  assign N243 = din[17] | din[16];
  assign N82 = ~N81;
  assign N83 = ~din[18];
  assign N84 = N275 | din[0];
  assign N275 = N274 | din[1];
  assign N274 = N273 | din[2];
  assign N273 = N272 | din[3];
  assign N272 = N271 | din[4];
  assign N271 = N270 | din[5];
  assign N270 = N269 | din[6];
  assign N269 = N268 | din[7];
  assign N268 = N267 | din[8];
  assign N267 = N266 | din[9];
  assign N266 = N265 | din[10];
  assign N265 = N264 | din[11];
  assign N264 = N263 | din[12];
  assign N263 = N262 | din[13];
  assign N262 = N261 | din[14];
  assign N261 = N260 | din[15];
  assign N260 = N259 | din[16];
  assign N259 = din[18] | din[17];
  assign N85 = ~N84;
  assign N86 = ~din[19];
  assign N87 = N293 | din[0];
  assign N293 = N292 | din[1];
  assign N292 = N291 | din[2];
  assign N291 = N290 | din[3];
  assign N290 = N289 | din[4];
  assign N289 = N288 | din[5];
  assign N288 = N287 | din[6];
  assign N287 = N286 | din[7];
  assign N286 = N285 | din[8];
  assign N285 = N284 | din[9];
  assign N284 = N283 | din[10];
  assign N283 = N282 | din[11];
  assign N282 = N281 | din[12];
  assign N281 = N280 | din[13];
  assign N280 = N279 | din[14];
  assign N279 = N278 | din[15];
  assign N278 = N277 | din[16];
  assign N277 = N276 | din[17];
  assign N276 = din[19] | din[18];
  assign N88 = ~N87;
  assign N89 = ~din[20];
  assign N90 = N312 | din[0];
  assign N312 = N311 | din[1];
  assign N311 = N310 | din[2];
  assign N310 = N309 | din[3];
  assign N309 = N308 | din[4];
  assign N308 = N307 | din[5];
  assign N307 = N306 | din[6];
  assign N306 = N305 | din[7];
  assign N305 = N304 | din[8];
  assign N304 = N303 | din[9];
  assign N303 = N302 | din[10];
  assign N302 = N301 | din[11];
  assign N301 = N300 | din[12];
  assign N300 = N299 | din[13];
  assign N299 = N298 | din[14];
  assign N298 = N297 | din[15];
  assign N297 = N296 | din[16];
  assign N296 = N295 | din[17];
  assign N295 = N294 | din[18];
  assign N294 = din[20] | din[19];
  assign N91 = ~N90;
  assign N92 = ~din[21];
  assign N93 = N332 | din[0];
  assign N332 = N331 | din[1];
  assign N331 = N330 | din[2];
  assign N330 = N329 | din[3];
  assign N329 = N328 | din[4];
  assign N328 = N327 | din[5];
  assign N327 = N326 | din[6];
  assign N326 = N325 | din[7];
  assign N325 = N324 | din[8];
  assign N324 = N323 | din[9];
  assign N323 = N322 | din[10];
  assign N322 = N321 | din[11];
  assign N321 = N320 | din[12];
  assign N320 = N319 | din[13];
  assign N319 = N318 | din[14];
  assign N318 = N317 | din[15];
  assign N317 = N316 | din[16];
  assign N316 = N315 | din[17];
  assign N315 = N314 | din[18];
  assign N314 = N313 | din[19];
  assign N313 = din[21] | din[20];
  assign N94 = ~N93;
  assign N95 = ~din[22];
  assign N96 = N353 | din[0];
  assign N353 = N352 | din[1];
  assign N352 = N351 | din[2];
  assign N351 = N350 | din[3];
  assign N350 = N349 | din[4];
  assign N349 = N348 | din[5];
  assign N348 = N347 | din[6];
  assign N347 = N346 | din[7];
  assign N346 = N345 | din[8];
  assign N345 = N344 | din[9];
  assign N344 = N343 | din[10];
  assign N343 = N342 | din[11];
  assign N342 = N341 | din[12];
  assign N341 = N340 | din[13];
  assign N340 = N339 | din[14];
  assign N339 = N338 | din[15];
  assign N338 = N337 | din[16];
  assign N337 = N336 | din[17];
  assign N336 = N335 | din[18];
  assign N335 = N334 | din[19];
  assign N334 = N333 | din[20];
  assign N333 = din[22] | din[21];
  assign N97 = ~N96;
  assign N98 = ~din[23];
  assign N99 = N375 | din[0];
  assign N375 = N374 | din[1];
  assign N374 = N373 | din[2];
  assign N373 = N372 | din[3];
  assign N372 = N371 | din[4];
  assign N371 = N370 | din[5];
  assign N370 = N369 | din[6];
  assign N369 = N368 | din[7];
  assign N368 = N367 | din[8];
  assign N367 = N366 | din[9];
  assign N366 = N365 | din[10];
  assign N365 = N364 | din[11];
  assign N364 = N363 | din[12];
  assign N363 = N362 | din[13];
  assign N362 = N361 | din[14];
  assign N361 = N360 | din[15];
  assign N360 = N359 | din[16];
  assign N359 = N358 | din[17];
  assign N358 = N357 | din[18];
  assign N357 = N356 | din[19];
  assign N356 = N355 | din[20];
  assign N355 = N354 | din[21];
  assign N354 = din[23] | din[22];
  assign N100 = ~N99;
  assign N101 = ~din[24];
  assign N102 = N398 | din[0];
  assign N398 = N397 | din[1];
  assign N397 = N396 | din[2];
  assign N396 = N395 | din[3];
  assign N395 = N394 | din[4];
  assign N394 = N393 | din[5];
  assign N393 = N392 | din[6];
  assign N392 = N391 | din[7];
  assign N391 = N390 | din[8];
  assign N390 = N389 | din[9];
  assign N389 = N388 | din[10];
  assign N388 = N387 | din[11];
  assign N387 = N386 | din[12];
  assign N386 = N385 | din[13];
  assign N385 = N384 | din[14];
  assign N384 = N383 | din[15];
  assign N383 = N382 | din[16];
  assign N382 = N381 | din[17];
  assign N381 = N380 | din[18];
  assign N380 = N379 | din[19];
  assign N379 = N378 | din[20];
  assign N378 = N377 | din[21];
  assign N377 = N376 | din[22];
  assign N376 = din[24] | din[23];
  assign N103 = ~N102;
  assign N104 = ~din[25];
  assign N105 = N422 | din[0];
  assign N422 = N421 | din[1];
  assign N421 = N420 | din[2];
  assign N420 = N419 | din[3];
  assign N419 = N418 | din[4];
  assign N418 = N417 | din[5];
  assign N417 = N416 | din[6];
  assign N416 = N415 | din[7];
  assign N415 = N414 | din[8];
  assign N414 = N413 | din[9];
  assign N413 = N412 | din[10];
  assign N412 = N411 | din[11];
  assign N411 = N410 | din[12];
  assign N410 = N409 | din[13];
  assign N409 = N408 | din[14];
  assign N408 = N407 | din[15];
  assign N407 = N406 | din[16];
  assign N406 = N405 | din[17];
  assign N405 = N404 | din[18];
  assign N404 = N403 | din[19];
  assign N403 = N402 | din[20];
  assign N402 = N401 | din[21];
  assign N401 = N400 | din[22];
  assign N400 = N399 | din[23];
  assign N399 = din[25] | din[24];
  assign N106 = ~N105;
  assign N107 = ~din[26];
  assign N108 = N447 | din[0];
  assign N447 = N446 | din[1];
  assign N446 = N445 | din[2];
  assign N445 = N444 | din[3];
  assign N444 = N443 | din[4];
  assign N443 = N442 | din[5];
  assign N442 = N441 | din[6];
  assign N441 = N440 | din[7];
  assign N440 = N439 | din[8];
  assign N439 = N438 | din[9];
  assign N438 = N437 | din[10];
  assign N437 = N436 | din[11];
  assign N436 = N435 | din[12];
  assign N435 = N434 | din[13];
  assign N434 = N433 | din[14];
  assign N433 = N432 | din[15];
  assign N432 = N431 | din[16];
  assign N431 = N430 | din[17];
  assign N430 = N429 | din[18];
  assign N429 = N428 | din[19];
  assign N428 = N427 | din[20];
  assign N427 = N426 | din[21];
  assign N426 = N425 | din[22];
  assign N425 = N424 | din[23];
  assign N424 = N423 | din[24];
  assign N423 = din[26] | din[25];
  assign N109 = ~N108;
  assign N110 = ~din[27];
  assign N111 = N473 | din[0];
  assign N473 = N472 | din[1];
  assign N472 = N471 | din[2];
  assign N471 = N470 | din[3];
  assign N470 = N469 | din[4];
  assign N469 = N468 | din[5];
  assign N468 = N467 | din[6];
  assign N467 = N466 | din[7];
  assign N466 = N465 | din[8];
  assign N465 = N464 | din[9];
  assign N464 = N463 | din[10];
  assign N463 = N462 | din[11];
  assign N462 = N461 | din[12];
  assign N461 = N460 | din[13];
  assign N460 = N459 | din[14];
  assign N459 = N458 | din[15];
  assign N458 = N457 | din[16];
  assign N457 = N456 | din[17];
  assign N456 = N455 | din[18];
  assign N455 = N454 | din[19];
  assign N454 = N453 | din[20];
  assign N453 = N452 | din[21];
  assign N452 = N451 | din[22];
  assign N451 = N450 | din[23];
  assign N450 = N449 | din[24];
  assign N449 = N448 | din[25];
  assign N448 = din[27] | din[26];
  assign N112 = ~N111;
  assign N113 = ~din[28];
  assign N114 = N500 | din[0];
  assign N500 = N499 | din[1];
  assign N499 = N498 | din[2];
  assign N498 = N497 | din[3];
  assign N497 = N496 | din[4];
  assign N496 = N495 | din[5];
  assign N495 = N494 | din[6];
  assign N494 = N493 | din[7];
  assign N493 = N492 | din[8];
  assign N492 = N491 | din[9];
  assign N491 = N490 | din[10];
  assign N490 = N489 | din[11];
  assign N489 = N488 | din[12];
  assign N488 = N487 | din[13];
  assign N487 = N486 | din[14];
  assign N486 = N485 | din[15];
  assign N485 = N484 | din[16];
  assign N484 = N483 | din[17];
  assign N483 = N482 | din[18];
  assign N482 = N481 | din[19];
  assign N481 = N480 | din[20];
  assign N480 = N479 | din[21];
  assign N479 = N478 | din[22];
  assign N478 = N477 | din[23];
  assign N477 = N476 | din[24];
  assign N476 = N475 | din[25];
  assign N475 = N474 | din[26];
  assign N474 = din[28] | din[27];
  assign N115 = ~N114;
  assign N116 = ~din[29];
  assign N117 = N528 | din[0];
  assign N528 = N527 | din[1];
  assign N527 = N526 | din[2];
  assign N526 = N525 | din[3];
  assign N525 = N524 | din[4];
  assign N524 = N523 | din[5];
  assign N523 = N522 | din[6];
  assign N522 = N521 | din[7];
  assign N521 = N520 | din[8];
  assign N520 = N519 | din[9];
  assign N519 = N518 | din[10];
  assign N518 = N517 | din[11];
  assign N517 = N516 | din[12];
  assign N516 = N515 | din[13];
  assign N515 = N514 | din[14];
  assign N514 = N513 | din[15];
  assign N513 = N512 | din[16];
  assign N512 = N511 | din[17];
  assign N511 = N510 | din[18];
  assign N510 = N509 | din[19];
  assign N509 = N508 | din[20];
  assign N508 = N507 | din[21];
  assign N507 = N506 | din[22];
  assign N506 = N505 | din[23];
  assign N505 = N504 | din[24];
  assign N504 = N503 | din[25];
  assign N503 = N502 | din[26];
  assign N502 = N501 | din[27];
  assign N501 = din[29] | din[28];
  assign N118 = ~N117;
  assign N119 = ~din[30];
  assign N120 = N557 | din[0];
  assign N557 = N556 | din[1];
  assign N556 = N555 | din[2];
  assign N555 = N554 | din[3];
  assign N554 = N553 | din[4];
  assign N553 = N552 | din[5];
  assign N552 = N551 | din[6];
  assign N551 = N550 | din[7];
  assign N550 = N549 | din[8];
  assign N549 = N548 | din[9];
  assign N548 = N547 | din[10];
  assign N547 = N546 | din[11];
  assign N546 = N545 | din[12];
  assign N545 = N544 | din[13];
  assign N544 = N543 | din[14];
  assign N543 = N542 | din[15];
  assign N542 = N541 | din[16];
  assign N541 = N540 | din[17];
  assign N540 = N539 | din[18];
  assign N539 = N538 | din[19];
  assign N538 = N537 | din[20];
  assign N537 = N536 | din[21];
  assign N536 = N535 | din[22];
  assign N535 = N534 | din[23];
  assign N534 = N533 | din[24];
  assign N533 = N532 | din[25];
  assign N532 = N531 | din[26];
  assign N531 = N530 | din[27];
  assign N530 = N529 | din[28];
  assign N529 = din[30] | din[29];
  assign N121 = ~N120;
  assign N122 = ~din[31];

endmodule