module bit_counter(clk, rs, count_right, do_popcnt, is_32bit, datalen, result);
  reg [63:0] _000_;
  reg [64:0] _001_;
  wire _002_;
  wire _003_;
  wire [63:0] _004_;
  wire _005_;
  wire [31:0] _006_;
  wire [63:0] _007_;
  wire [63:0] _008_;
  wire [64:0] _009_;
  wire [63:0] _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire [63:0] _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  reg [3:0] _327_;
  reg _328_;
  reg [31:0] _329_;
  wire [1:0] _330_;
  wire [1:0] _331_;
  wire [1:0] _332_;
  wire [1:0] _333_;
  wire [1:0] _334_;
  wire [1:0] _335_;
  wire [1:0] _336_;
  wire [1:0] _337_;
  wire [1:0] _338_;
  wire [1:0] _339_;
  wire [1:0] _340_;
  wire [1:0] _341_;
  wire [1:0] _342_;
  wire [1:0] _343_;
  wire [1:0] _344_;
  wire [1:0] _345_;
  wire [1:0] _346_;
  wire [1:0] _347_;
  wire [1:0] _348_;
  wire [1:0] _349_;
  wire [1:0] _350_;
  wire [1:0] _351_;
  wire [1:0] _352_;
  wire [1:0] _353_;
  wire [1:0] _354_;
  wire [1:0] _355_;
  wire [1:0] _356_;
  wire [1:0] _357_;
  wire [1:0] _358_;
  wire [1:0] _359_;
  wire [1:0] _360_;
  wire [1:0] _361_;
  wire [2:0] _362_;
  wire [2:0] _363_;
  wire [2:0] _364_;
  wire [2:0] _365_;
  wire [2:0] _366_;
  wire [2:0] _367_;
  wire [2:0] _368_;
  wire [2:0] _369_;
  wire [2:0] _370_;
  wire [2:0] _371_;
  wire [2:0] _372_;
  wire [2:0] _373_;
  wire [2:0] _374_;
  wire [2:0] _375_;
  wire [2:0] _376_;
  wire [2:0] _377_;
  wire [3:0] _378_;
  wire [3:0] _379_;
  wire [3:0] _380_;
  wire [3:0] _381_;
  wire [3:0] _382_;
  wire [3:0] _383_;
  wire [3:0] _384_;
  wire [3:0] _385_;
  wire [5:0] _386_;
  wire [5:0] _387_;
  wire [5:0] _388_;
  wire [5:0] _389_;
  wire [5:0] _390_;
  wire [5:0] _391_;
  wire _392_;
  wire _393_;
  wire [6:0] _394_;
  wire [5:0] _395_;
  wire _396_;
  wire [5:0] _397_;
  wire [3:0] _398_;
  wire [2:0] _399_;
  wire [3:0] _400_;
  wire [3:0] _401_;
  wire [3:0] _402_;
  wire [3:0] _403_;
  wire [1:0] _404_;
  wire [3:0] _405_;
  wire [3:0] _406_;
  wire [3:0] _407_;
  wire _408_;
  wire [63:0] _409_;
  wire [5:0] bitnum;
  input clk;
  wire clk;
  wire [63:0] cntz;
  input count_right;
  wire count_right;
  input [3:0] datalen;
  wire [3:0] datalen;
  wire [3:0] dlen_r;
  input do_popcnt;
  wire do_popcnt;
  wire [63:0] \edge ;
  wire [63:0] inp;
  wire [63:0] inp_r;
  input is_32bit;
  wire is_32bit;
  wire [63:0] onehot;
  wire [63:0] pc2;
  wire [11:0] pc32;
  wire [47:0] pc4;
  wire [31:0] pc8;
  wire [31:0] pc8_r;
  wire pcnt_r;
  wire [63:0] popcnt;
  output [63:0] result;
  wire [63:0] result;
  input [63:0] rs;
  wire [63:0] rs;
  wire [64:0] sum;
  wire [64:0] sum_r;
  always @(posedge clk)
    _000_ <= inp;
  always @(posedge clk)
    _001_ <= sum;
  assign _002_ = ~ is_32bit;
  assign _003_ = ~ count_right;
  assign _004_ = _003_ ? { rs[0], rs[1], rs[2], rs[3], rs[4], rs[5], rs[6], rs[7], rs[8], rs[9], rs[10], rs[11], rs[12], rs[13], rs[14], rs[15], rs[16], rs[17], rs[18], rs[19], rs[20], rs[21], rs[22], rs[23], rs[24], rs[25], rs[26], rs[27], rs[28], rs[29], rs[30], rs[31], rs[32], rs[33], rs[34], rs[35], rs[36], rs[37], rs[38], rs[39], rs[40], rs[41], rs[42], rs[43], rs[44], rs[45], rs[46], rs[47], rs[48], rs[49], rs[50], rs[51], rs[52], rs[53], rs[54], rs[55], rs[56], rs[57], rs[58], rs[59], rs[60], rs[61], rs[62], rs[63] } : rs;
  assign _005_ = ~ count_right;
  assign _006_ = _005_ ? { rs[0], rs[1], rs[2], rs[3], rs[4], rs[5], rs[6], rs[7], rs[8], rs[9], rs[10], rs[11], rs[12], rs[13], rs[14], rs[15], rs[16], rs[17], rs[18], rs[19], rs[20], rs[21], rs[22], rs[23], rs[24], rs[25], rs[26], rs[27], rs[28], rs[29], rs[30], rs[31] } : rs[31:0];
  assign _007_ = _002_ ? _004_ : { 32'hffffffff, _006_ };
  assign _008_ = ~ inp;
  assign _009_ = { 1'h0, _008_ } + 65'h00000000000000001;
  assign _010_ = sum_r[63:0] | inp_r;
  assign _011_ = ~ \edge [0];
  assign _012_ = \edge [1] & _011_;
  assign _013_ = 1'h0 | _012_;
  assign _014_ = ~ \edge [2];
  assign _015_ = \edge [3] & _014_;
  assign _016_ = _013_ | _015_;
  assign _017_ = ~ \edge [4];
  assign _018_ = \edge [5] & _017_;
  assign _019_ = _016_ | _018_;
  assign _020_ = ~ \edge [6];
  assign _021_ = \edge [7] & _020_;
  assign _022_ = _019_ | _021_;
  assign _023_ = ~ \edge [8];
  assign _024_ = \edge [9] & _023_;
  assign _025_ = _022_ | _024_;
  assign _026_ = ~ \edge [10];
  assign _027_ = \edge [11] & _026_;
  assign _028_ = _025_ | _027_;
  assign _029_ = ~ \edge [12];
  assign _030_ = \edge [13] & _029_;
  assign _031_ = _028_ | _030_;
  assign _032_ = ~ \edge [14];
  assign _033_ = \edge [15] & _032_;
  assign _034_ = _031_ | _033_;
  assign _035_ = ~ \edge [16];
  assign _036_ = \edge [17] & _035_;
  assign _037_ = _034_ | _036_;
  assign _038_ = ~ \edge [18];
  assign _039_ = \edge [19] & _038_;
  assign _040_ = _037_ | _039_;
  assign _041_ = ~ \edge [20];
  assign _042_ = \edge [21] & _041_;
  assign _043_ = _040_ | _042_;
  assign _044_ = ~ \edge [22];
  assign _045_ = \edge [23] & _044_;
  assign _046_ = _043_ | _045_;
  assign _047_ = ~ \edge [24];
  assign _048_ = \edge [25] & _047_;
  assign _049_ = _046_ | _048_;
  assign _050_ = ~ \edge [26];
  assign _051_ = \edge [27] & _050_;
  assign _052_ = _049_ | _051_;
  assign _053_ = ~ \edge [28];
  assign _054_ = \edge [29] & _053_;
  assign _055_ = _052_ | _054_;
  assign _056_ = ~ \edge [30];
  assign _057_ = \edge [31] & _056_;
  assign _058_ = _055_ | _057_;
  assign _059_ = ~ \edge [32];
  assign _060_ = \edge [33] & _059_;
  assign _061_ = _058_ | _060_;
  assign _062_ = ~ \edge [34];
  assign _063_ = \edge [35] & _062_;
  assign _064_ = _061_ | _063_;
  assign _065_ = ~ \edge [36];
  assign _066_ = \edge [37] & _065_;
  assign _067_ = _064_ | _066_;
  assign _068_ = ~ \edge [38];
  assign _069_ = \edge [39] & _068_;
  assign _070_ = _067_ | _069_;
  assign _071_ = ~ \edge [40];
  assign _072_ = \edge [41] & _071_;
  assign _073_ = _070_ | _072_;
  assign _074_ = ~ \edge [42];
  assign _075_ = \edge [43] & _074_;
  assign _076_ = _073_ | _075_;
  assign _077_ = ~ \edge [44];
  assign _078_ = \edge [45] & _077_;
  assign _079_ = _076_ | _078_;
  assign _080_ = ~ \edge [46];
  assign _081_ = \edge [47] & _080_;
  assign _082_ = _079_ | _081_;
  assign _083_ = ~ \edge [48];
  assign _084_ = \edge [49] & _083_;
  assign _085_ = _082_ | _084_;
  assign _086_ = ~ \edge [50];
  assign _087_ = \edge [51] & _086_;
  assign _088_ = _085_ | _087_;
  assign _089_ = ~ \edge [52];
  assign _090_ = \edge [53] & _089_;
  assign _091_ = _088_ | _090_;
  assign _092_ = ~ \edge [54];
  assign _093_ = \edge [55] & _092_;
  assign _094_ = _091_ | _093_;
  assign _095_ = ~ \edge [56];
  assign _096_ = \edge [57] & _095_;
  assign _097_ = _094_ | _096_;
  assign _098_ = ~ \edge [58];
  assign _099_ = \edge [59] & _098_;
  assign _100_ = _097_ | _099_;
  assign _101_ = ~ \edge [60];
  assign _102_ = \edge [61] & _101_;
  assign _103_ = _100_ | _102_;
  assign _104_ = ~ \edge [62];
  assign _105_ = \edge [63] & _104_;
  assign _106_ = _103_ | _105_;
  assign _107_ = ~ \edge [1];
  assign _108_ = \edge [3] & _107_;
  assign _109_ = 1'h0 | _108_;
  assign _110_ = ~ \edge [5];
  assign _111_ = \edge [7] & _110_;
  assign _112_ = _109_ | _111_;
  assign _113_ = ~ \edge [9];
  assign _114_ = \edge [11] & _113_;
  assign _115_ = _112_ | _114_;
  assign _116_ = ~ \edge [13];
  assign _117_ = \edge [15] & _116_;
  assign _118_ = _115_ | _117_;
  assign _119_ = ~ \edge [17];
  assign _120_ = \edge [19] & _119_;
  assign _121_ = _118_ | _120_;
  assign _122_ = ~ \edge [21];
  assign _123_ = \edge [23] & _122_;
  assign _124_ = _121_ | _123_;
  assign _125_ = ~ \edge [25];
  assign _126_ = \edge [27] & _125_;
  assign _127_ = _124_ | _126_;
  assign _128_ = ~ \edge [29];
  assign _129_ = \edge [31] & _128_;
  assign _130_ = _127_ | _129_;
  assign _131_ = ~ \edge [33];
  assign _132_ = \edge [35] & _131_;
  assign _133_ = _130_ | _132_;
  assign _134_ = ~ \edge [37];
  assign _135_ = \edge [39] & _134_;
  assign _136_ = _133_ | _135_;
  assign _137_ = ~ \edge [41];
  assign _138_ = \edge [43] & _137_;
  assign _139_ = _136_ | _138_;
  assign _140_ = ~ \edge [45];
  assign _141_ = \edge [47] & _140_;
  assign _142_ = _139_ | _141_;
  assign _143_ = ~ \edge [49];
  assign _144_ = \edge [51] & _143_;
  assign _145_ = _142_ | _144_;
  assign _146_ = ~ \edge [53];
  assign _147_ = \edge [55] & _146_;
  assign _148_ = _145_ | _147_;
  assign _149_ = ~ \edge [57];
  assign _150_ = \edge [59] & _149_;
  assign _151_ = _148_ | _150_;
  assign _152_ = ~ \edge [61];
  assign _153_ = \edge [63] & _152_;
  assign _154_ = _151_ | _153_;
  assign _155_ = ~ \edge [3];
  assign _156_ = \edge [7] & _155_;
  assign _157_ = 1'h0 | _156_;
  assign _158_ = ~ \edge [11];
  assign _159_ = \edge [15] & _158_;
  assign _160_ = _157_ | _159_;
  assign _161_ = ~ \edge [19];
  assign _162_ = \edge [23] & _161_;
  assign _163_ = _160_ | _162_;
  assign _164_ = ~ \edge [27];
  assign _165_ = \edge [31] & _164_;
  assign _166_ = _163_ | _165_;
  assign _167_ = ~ \edge [35];
  assign _168_ = \edge [39] & _167_;
  assign _169_ = _166_ | _168_;
  assign _170_ = ~ \edge [43];
  assign _171_ = \edge [47] & _170_;
  assign _172_ = _169_ | _171_;
  assign _173_ = ~ \edge [51];
  assign _174_ = \edge [55] & _173_;
  assign _175_ = _172_ | _174_;
  assign _176_ = ~ \edge [59];
  assign _177_ = \edge [63] & _176_;
  assign _178_ = _175_ | _177_;
  assign _179_ = ~ \edge [7];
  assign _180_ = \edge [15] & _179_;
  assign _181_ = 1'h0 | _180_;
  assign _182_ = ~ \edge [23];
  assign _183_ = \edge [31] & _182_;
  assign _184_ = _181_ | _183_;
  assign _185_ = ~ \edge [39];
  assign _186_ = \edge [47] & _185_;
  assign _187_ = _184_ | _186_;
  assign _188_ = ~ \edge [55];
  assign _189_ = \edge [63] & _188_;
  assign _190_ = _187_ | _189_;
  assign _191_ = ~ \edge [15];
  assign _192_ = \edge [31] & _191_;
  assign _193_ = 1'h0 | _192_;
  assign _194_ = ~ \edge [47];
  assign _195_ = \edge [63] & _194_;
  assign _196_ = _193_ | _195_;
  assign _197_ = ~ \edge [31];
  assign _198_ = \edge [63] & _197_;
  assign _199_ = 1'h0 | _198_;
  assign _200_ = sum_r[63:0] & inp_r;
  assign _201_ = | onehot[1];
  assign _202_ = 1'h0 | _201_;
  assign _203_ = | onehot[3];
  assign _204_ = _202_ | _203_;
  assign _205_ = | onehot[5];
  assign _206_ = _204_ | _205_;
  assign _207_ = | onehot[7];
  assign _208_ = _206_ | _207_;
  assign _209_ = | onehot[9];
  assign _210_ = _208_ | _209_;
  assign _211_ = | onehot[11];
  assign _212_ = _210_ | _211_;
  assign _213_ = | onehot[13];
  assign _214_ = _212_ | _213_;
  assign _215_ = | onehot[15];
  assign _216_ = _214_ | _215_;
  assign _217_ = | onehot[17];
  assign _218_ = _216_ | _217_;
  assign _219_ = | onehot[19];
  assign _220_ = _218_ | _219_;
  assign _221_ = | onehot[21];
  assign _222_ = _220_ | _221_;
  assign _223_ = | onehot[23];
  assign _224_ = _222_ | _223_;
  assign _225_ = | onehot[25];
  assign _226_ = _224_ | _225_;
  assign _227_ = | onehot[27];
  assign _228_ = _226_ | _227_;
  assign _229_ = | onehot[29];
  assign _230_ = _228_ | _229_;
  assign _231_ = | onehot[31];
  assign _232_ = _230_ | _231_;
  assign _233_ = | onehot[33];
  assign _234_ = _232_ | _233_;
  assign _235_ = | onehot[35];
  assign _236_ = _234_ | _235_;
  assign _237_ = | onehot[37];
  assign _238_ = _236_ | _237_;
  assign _239_ = | onehot[39];
  assign _240_ = _238_ | _239_;
  assign _241_ = | onehot[41];
  assign _242_ = _240_ | _241_;
  assign _243_ = | onehot[43];
  assign _244_ = _242_ | _243_;
  assign _245_ = | onehot[45];
  assign _246_ = _244_ | _245_;
  assign _247_ = | onehot[47];
  assign _248_ = _246_ | _247_;
  assign _249_ = | onehot[49];
  assign _250_ = _248_ | _249_;
  assign _251_ = | onehot[51];
  assign _252_ = _250_ | _251_;
  assign _253_ = | onehot[53];
  assign _254_ = _252_ | _253_;
  assign _255_ = | onehot[55];
  assign _256_ = _254_ | _255_;
  assign _257_ = | onehot[57];
  assign _258_ = _256_ | _257_;
  assign _259_ = | onehot[59];
  assign _260_ = _258_ | _259_;
  assign _261_ = | onehot[61];
  assign _262_ = _260_ | _261_;
  assign _263_ = | onehot[63];
  assign _264_ = _262_ | _263_;
  assign _265_ = | onehot[3:2];
  assign _266_ = 1'h0 | _265_;
  assign _267_ = | onehot[7:6];
  assign _268_ = _266_ | _267_;
  assign _269_ = | onehot[11:10];
  assign _270_ = _268_ | _269_;
  assign _271_ = | onehot[15:14];
  assign _272_ = _270_ | _271_;
  assign _273_ = | onehot[19:18];
  assign _274_ = _272_ | _273_;
  assign _275_ = | onehot[23:22];
  assign _276_ = _274_ | _275_;
  assign _277_ = | onehot[27:26];
  assign _278_ = _276_ | _277_;
  assign _279_ = | onehot[31:30];
  assign _280_ = _278_ | _279_;
  assign _281_ = | onehot[35:34];
  assign _282_ = _280_ | _281_;
  assign _283_ = | onehot[39:38];
  assign _284_ = _282_ | _283_;
  assign _285_ = | onehot[43:42];
  assign _286_ = _284_ | _285_;
  assign _287_ = | onehot[47:46];
  assign _288_ = _286_ | _287_;
  assign _289_ = | onehot[51:50];
  assign _290_ = _288_ | _289_;
  assign _291_ = | onehot[55:54];
  assign _292_ = _290_ | _291_;
  assign _293_ = | onehot[59:58];
  assign _294_ = _292_ | _293_;
  assign _295_ = | onehot[63:62];
  assign _296_ = _294_ | _295_;
  assign _297_ = | onehot[7:4];
  assign _298_ = 1'h0 | _297_;
  assign _299_ = | onehot[15:12];
  assign _300_ = _298_ | _299_;
  assign _301_ = | onehot[23:20];
  assign _302_ = _300_ | _301_;
  assign _303_ = | onehot[31:28];
  assign _304_ = _302_ | _303_;
  assign _305_ = | onehot[39:36];
  assign _306_ = _304_ | _305_;
  assign _307_ = | onehot[47:44];
  assign _308_ = _306_ | _307_;
  assign _309_ = | onehot[55:52];
  assign _310_ = _308_ | _309_;
  assign _311_ = | onehot[63:60];
  assign _312_ = _310_ | _311_;
  assign _313_ = | onehot[15:8];
  assign _314_ = 1'h0 | _313_;
  assign _315_ = | onehot[31:24];
  assign _316_ = _314_ | _315_;
  assign _317_ = | onehot[47:40];
  assign _318_ = _316_ | _317_;
  assign _319_ = | onehot[63:56];
  assign _320_ = _318_ | _319_;
  assign _321_ = | onehot[31:16];
  assign _322_ = 1'h0 | _321_;
  assign _323_ = | onehot[63:48];
  assign _324_ = _322_ | _323_;
  assign _325_ = | onehot[63:32];
  assign _326_ = 1'h0 | _325_;
  always @(posedge clk)
    _327_ <= datalen;
  always @(posedge clk)
    _328_ <= do_popcnt;
  always @(posedge clk)
    _329_ <= pc8;
  assign _330_ = { 1'h0, rs[0] } + { 1'h0, rs[1] };
  assign _331_ = { 1'h0, rs[2] } + { 1'h0, rs[3] };
  assign _332_ = { 1'h0, rs[4] } + { 1'h0, rs[5] };
  assign _333_ = { 1'h0, rs[6] } + { 1'h0, rs[7] };
  assign _334_ = { 1'h0, rs[8] } + { 1'h0, rs[9] };
  assign _335_ = { 1'h0, rs[10] } + { 1'h0, rs[11] };
  assign _336_ = { 1'h0, rs[12] } + { 1'h0, rs[13] };
  assign _337_ = { 1'h0, rs[14] } + { 1'h0, rs[15] };
  assign _338_ = { 1'h0, rs[16] } + { 1'h0, rs[17] };
  assign _339_ = { 1'h0, rs[18] } + { 1'h0, rs[19] };
  assign _340_ = { 1'h0, rs[20] } + { 1'h0, rs[21] };
  assign _341_ = { 1'h0, rs[22] } + { 1'h0, rs[23] };
  assign _342_ = { 1'h0, rs[24] } + { 1'h0, rs[25] };
  assign _343_ = { 1'h0, rs[26] } + { 1'h0, rs[27] };
  assign _344_ = { 1'h0, rs[28] } + { 1'h0, rs[29] };
  assign _345_ = { 1'h0, rs[30] } + { 1'h0, rs[31] };
  assign _346_ = { 1'h0, rs[32] } + { 1'h0, rs[33] };
  assign _347_ = { 1'h0, rs[34] } + { 1'h0, rs[35] };
  assign _348_ = { 1'h0, rs[36] } + { 1'h0, rs[37] };
  assign _349_ = { 1'h0, rs[38] } + { 1'h0, rs[39] };
  assign _350_ = { 1'h0, rs[40] } + { 1'h0, rs[41] };
  assign _351_ = { 1'h0, rs[42] } + { 1'h0, rs[43] };
  assign _352_ = { 1'h0, rs[44] } + { 1'h0, rs[45] };
  assign _353_ = { 1'h0, rs[46] } + { 1'h0, rs[47] };
  assign _354_ = { 1'h0, rs[48] } + { 1'h0, rs[49] };
  assign _355_ = { 1'h0, rs[50] } + { 1'h0, rs[51] };
  assign _356_ = { 1'h0, rs[52] } + { 1'h0, rs[53] };
  assign _357_ = { 1'h0, rs[54] } + { 1'h0, rs[55] };
  assign _358_ = { 1'h0, rs[56] } + { 1'h0, rs[57] };
  assign _359_ = { 1'h0, rs[58] } + { 1'h0, rs[59] };
  assign _360_ = { 1'h0, rs[60] } + { 1'h0, rs[61] };
  assign _361_ = { 1'h0, rs[62] } + { 1'h0, rs[63] };
  assign _362_ = { 1'h0, pc2[63:62] } + { 1'h0, pc2[61:60] };
  assign _363_ = { 1'h0, pc2[59:58] } + { 1'h0, pc2[57:56] };
  assign _364_ = { 1'h0, pc2[55:54] } + { 1'h0, pc2[53:52] };
  assign _365_ = { 1'h0, pc2[51:50] } + { 1'h0, pc2[49:48] };
  assign _366_ = { 1'h0, pc2[47:46] } + { 1'h0, pc2[45:44] };
  assign _367_ = { 1'h0, pc2[43:42] } + { 1'h0, pc2[41:40] };
  assign _368_ = { 1'h0, pc2[39:38] } + { 1'h0, pc2[37:36] };
  assign _369_ = { 1'h0, pc2[35:34] } + { 1'h0, pc2[33:32] };
  assign _370_ = { 1'h0, pc2[31:30] } + { 1'h0, pc2[29:28] };
  assign _371_ = { 1'h0, pc2[27:26] } + { 1'h0, pc2[25:24] };
  assign _372_ = { 1'h0, pc2[23:22] } + { 1'h0, pc2[21:20] };
  assign _373_ = { 1'h0, pc2[19:18] } + { 1'h0, pc2[17:16] };
  assign _374_ = { 1'h0, pc2[15:14] } + { 1'h0, pc2[13:12] };
  assign _375_ = { 1'h0, pc2[11:10] } + { 1'h0, pc2[9:8] };
  assign _376_ = { 1'h0, pc2[7:6] } + { 1'h0, pc2[5:4] };
  assign _377_ = { 1'h0, pc2[3:2] } + { 1'h0, pc2[1:0] };
  assign _378_ = { 1'h0, pc4[47:45] } + { 1'h0, pc4[44:42] };
  assign _379_ = { 1'h0, pc4[41:39] } + { 1'h0, pc4[38:36] };
  assign _380_ = { 1'h0, pc4[35:33] } + { 1'h0, pc4[32:30] };
  assign _381_ = { 1'h0, pc4[29:27] } + { 1'h0, pc4[26:24] };
  assign _382_ = { 1'h0, pc4[23:21] } + { 1'h0, pc4[20:18] };
  assign _383_ = { 1'h0, pc4[17:15] } + { 1'h0, pc4[14:12] };
  assign _384_ = { 1'h0, pc4[11:9] } + { 1'h0, pc4[8:6] };
  assign _385_ = { 1'h0, pc4[5:3] } + { 1'h0, pc4[2:0] };
  assign _386_ = { 2'h0, pc8_r[31:28] } + { 2'h0, pc8_r[27:24] };
  assign _387_ = _386_ + { 2'h0, pc8_r[23:20] };
  assign _388_ = _387_ + { 2'h0, pc8_r[19:16] };
  assign _389_ = { 2'h0, pc8_r[15:12] } + { 2'h0, pc8_r[11:8] };
  assign _390_ = _389_ + { 2'h0, pc8_r[7:4] };
  assign _391_ = _390_ + { 2'h0, pc8_r[3:0] };
  assign _392_ = dlen_r[3:2] == 2'h0;
  assign _393_ = ~ dlen_r[3];
  assign _394_ = { 1'h0, pc32[11:6] } + { 1'h0, pc32[5:0] };
  assign _395_ = _393_ ? pc32[11:6] : _394_[5:0];
  assign _396_ = _393_ ? 1'h0 : _394_[6];
  assign _397_ = _393_ ? pc32[5:0] : 6'h00;
  assign _398_ = _392_ ? pc8_r[31:28] : _395_[3:0];
  assign _399_ = _392_ ? 3'h0 : { _396_, _395_[5:4] };
  assign _400_ = _392_ ? pc8_r[27:24] : 4'h0;
  assign _401_ = _392_ ? pc8_r[23:20] : 4'h0;
  assign _402_ = _392_ ? pc8_r[19:16] : 4'h0;
  assign _403_ = _392_ ? pc8_r[15:12] : _397_[3:0];
  assign _404_ = _392_ ? 2'h0 : _397_[5:4];
  assign _405_ = _392_ ? pc8_r[11:8] : 4'h0;
  assign _406_ = _392_ ? pc8_r[7:4] : 4'h0;
  assign _407_ = _392_ ? pc8_r[3:0] : 4'h0;
  assign _408_ = ~ pcnt_r;
  assign _409_ = _408_ ? cntz : popcnt;
  assign inp = _007_;
  assign inp_r = _000_;
  assign sum = _009_;
  assign sum_r = _001_;
  assign onehot = _200_;
  assign \edge  = _010_;
  assign bitnum = { _199_, _196_, _190_, _178_, _296_, _264_ };
  assign cntz = { 57'h000000000000000, sum_r[64], bitnum };
  assign dlen_r = _327_;
  assign pcnt_r = _328_;
  assign pc2 = { _330_, _331_, _332_, _333_, _334_, _335_, _336_, _337_, _338_, _339_, _340_, _341_, _342_, _343_, _344_, _345_, _346_, _347_, _348_, _349_, _350_, _351_, _352_, _353_, _354_, _355_, _356_, _357_, _358_, _359_, _360_, _361_ };
  assign pc4 = { _362_, _363_, _364_, _365_, _366_, _367_, _368_, _369_, _370_, _371_, _372_, _373_, _374_, _375_, _376_, _377_ };
  assign pc8 = { _378_, _379_, _380_, _381_, _382_, _383_, _384_, _385_ };
  assign pc8_r = _329_;
  assign pc32 = { _388_, _391_ };
  assign popcnt = { 4'h0, _407_, 4'h0, _406_, 4'h0, _405_, 2'h0, _404_, _403_, 4'h0, _402_, 4'h0, _401_, 4'h0, _400_, 1'h0, _399_, _398_ };
  assign result = _409_;
endmodule