module HellaCacheArbiter
(
  clk,
  io_requestor_2_req_ready,
  io_requestor_2_req_valid,
  io_requestor_2_req_bits_addr,
  io_requestor_2_req_bits_tag,
  io_requestor_2_req_bits_cmd,
  io_requestor_2_req_bits_typ,
  io_requestor_2_req_bits_kill,
  io_requestor_2_req_bits_phys,
  io_requestor_2_req_bits_data,
  io_requestor_2_resp_valid,
  io_requestor_2_resp_bits_addr,
  io_requestor_2_resp_bits_tag,
  io_requestor_2_resp_bits_cmd,
  io_requestor_2_resp_bits_typ,
  io_requestor_2_resp_bits_data,
  io_requestor_2_resp_bits_nack,
  io_requestor_2_resp_bits_replay,
  io_requestor_2_resp_bits_has_data,
  io_requestor_2_resp_bits_data_word_bypass,
  io_requestor_2_resp_bits_store_data,
  io_requestor_2_replay_next_valid,
  io_requestor_2_replay_next_bits,
  io_requestor_2_xcpt_ma_ld,
  io_requestor_2_xcpt_ma_st,
  io_requestor_2_xcpt_pf_ld,
  io_requestor_2_xcpt_pf_st,
  io_requestor_2_ordered,
  io_requestor_1_req_ready,
  io_requestor_1_req_valid,
  io_requestor_1_req_bits_addr,
  io_requestor_1_req_bits_tag,
  io_requestor_1_req_bits_cmd,
  io_requestor_1_req_bits_typ,
  io_requestor_1_req_bits_kill,
  io_requestor_1_req_bits_phys,
  io_requestor_1_req_bits_data,
  io_requestor_1_resp_valid,
  io_requestor_1_resp_bits_addr,
  io_requestor_1_resp_bits_tag,
  io_requestor_1_resp_bits_cmd,
  io_requestor_1_resp_bits_typ,
  io_requestor_1_resp_bits_data,
  io_requestor_1_resp_bits_nack,
  io_requestor_1_resp_bits_replay,
  io_requestor_1_resp_bits_has_data,
  io_requestor_1_resp_bits_data_word_bypass,
  io_requestor_1_resp_bits_store_data,
  io_requestor_1_replay_next_valid,
  io_requestor_1_replay_next_bits,
  io_requestor_1_xcpt_ma_ld,
  io_requestor_1_xcpt_ma_st,
  io_requestor_1_xcpt_pf_ld,
  io_requestor_1_xcpt_pf_st,
  io_requestor_1_invalidate_lr,
  io_requestor_1_ordered,
  io_requestor_0_req_ready,
  io_requestor_0_req_valid,
  io_requestor_0_req_bits_addr,
  io_requestor_0_req_bits_tag,
  io_requestor_0_req_bits_cmd,
  io_requestor_0_req_bits_typ,
  io_requestor_0_req_bits_kill,
  io_requestor_0_req_bits_phys,
  io_requestor_0_req_bits_data,
  io_requestor_0_resp_valid,
  io_requestor_0_resp_bits_addr,
  io_requestor_0_resp_bits_tag,
  io_requestor_0_resp_bits_cmd,
  io_requestor_0_resp_bits_typ,
  io_requestor_0_resp_bits_data,
  io_requestor_0_resp_bits_nack,
  io_requestor_0_resp_bits_replay,
  io_requestor_0_resp_bits_has_data,
  io_requestor_0_resp_bits_data_word_bypass,
  io_requestor_0_resp_bits_store_data,
  io_requestor_0_replay_next_valid,
  io_requestor_0_replay_next_bits,
  io_requestor_0_xcpt_ma_ld,
  io_requestor_0_xcpt_ma_st,
  io_requestor_0_xcpt_pf_ld,
  io_requestor_0_xcpt_pf_st,
  io_requestor_0_ordered,
  io_mem_req_ready,
  io_mem_req_valid,
  io_mem_req_bits_addr,
  io_mem_req_bits_tag,
  io_mem_req_bits_cmd,
  io_mem_req_bits_typ,
  io_mem_req_bits_kill,
  io_mem_req_bits_phys,
  io_mem_req_bits_data,
  io_mem_resp_valid,
  io_mem_resp_bits_addr,
  io_mem_resp_bits_tag,
  io_mem_resp_bits_cmd,
  io_mem_resp_bits_typ,
  io_mem_resp_bits_data,
  io_mem_resp_bits_nack,
  io_mem_resp_bits_replay,
  io_mem_resp_bits_has_data,
  io_mem_resp_bits_data_word_bypass,
  io_mem_resp_bits_store_data,
  io_mem_replay_next_valid,
  io_mem_replay_next_bits,
  io_mem_xcpt_ma_ld,
  io_mem_xcpt_ma_st,
  io_mem_xcpt_pf_ld,
  io_mem_xcpt_pf_st,
  io_mem_ordered
);

  input [39:0] io_requestor_2_req_bits_addr;
  input [9:0] io_requestor_2_req_bits_tag;
  input [4:0] io_requestor_2_req_bits_cmd;
  input [2:0] io_requestor_2_req_bits_typ;
  input [63:0] io_requestor_2_req_bits_data;
  output [39:0] io_requestor_2_resp_bits_addr;
  output [9:0] io_requestor_2_resp_bits_tag;
  output [4:0] io_requestor_2_resp_bits_cmd;
  output [2:0] io_requestor_2_resp_bits_typ;
  output [63:0] io_requestor_2_resp_bits_data;
  output [63:0] io_requestor_2_resp_bits_data_word_bypass;
  output [63:0] io_requestor_2_resp_bits_store_data;
  output [9:0] io_requestor_2_replay_next_bits;
  input [39:0] io_requestor_1_req_bits_addr;
  input [9:0] io_requestor_1_req_bits_tag;
  input [4:0] io_requestor_1_req_bits_cmd;
  input [2:0] io_requestor_1_req_bits_typ;
  input [63:0] io_requestor_1_req_bits_data;
  output [39:0] io_requestor_1_resp_bits_addr;
  output [9:0] io_requestor_1_resp_bits_tag;
  output [4:0] io_requestor_1_resp_bits_cmd;
  output [2:0] io_requestor_1_resp_bits_typ;
  output [63:0] io_requestor_1_resp_bits_data;
  output [63:0] io_requestor_1_resp_bits_data_word_bypass;
  output [63:0] io_requestor_1_resp_bits_store_data;
  output [9:0] io_requestor_1_replay_next_bits;
  input [39:0] io_requestor_0_req_bits_addr;
  input [9:0] io_requestor_0_req_bits_tag;
  input [4:0] io_requestor_0_req_bits_cmd;
  input [2:0] io_requestor_0_req_bits_typ;
  input [63:0] io_requestor_0_req_bits_data;
  output [39:0] io_requestor_0_resp_bits_addr;
  output [9:0] io_requestor_0_resp_bits_tag;
  output [4:0] io_requestor_0_resp_bits_cmd;
  output [2:0] io_requestor_0_resp_bits_typ;
  output [63:0] io_requestor_0_resp_bits_data;
  output [63:0] io_requestor_0_resp_bits_data_word_bypass;
  output [63:0] io_requestor_0_resp_bits_store_data;
  output [9:0] io_requestor_0_replay_next_bits;
  output [39:0] io_mem_req_bits_addr;
  output [9:0] io_mem_req_bits_tag;
  output [4:0] io_mem_req_bits_cmd;
  output [2:0] io_mem_req_bits_typ;
  output [63:0] io_mem_req_bits_data;
  input [39:0] io_mem_resp_bits_addr;
  input [9:0] io_mem_resp_bits_tag;
  input [4:0] io_mem_resp_bits_cmd;
  input [2:0] io_mem_resp_bits_typ;
  input [63:0] io_mem_resp_bits_data;
  input [63:0] io_mem_resp_bits_data_word_bypass;
  input [63:0] io_mem_resp_bits_store_data;
  input [9:0] io_mem_replay_next_bits;
  input clk;
  input io_requestor_2_req_valid;
  input io_requestor_2_req_bits_kill;
  input io_requestor_2_req_bits_phys;
  input io_requestor_1_req_valid;
  input io_requestor_1_req_bits_kill;
  input io_requestor_1_req_bits_phys;
  input io_requestor_1_invalidate_lr;
  input io_requestor_0_req_valid;
  input io_requestor_0_req_bits_kill;
  input io_requestor_0_req_bits_phys;
  input io_mem_req_ready;
  input io_mem_resp_valid;
  input io_mem_resp_bits_nack;
  input io_mem_resp_bits_replay;
  input io_mem_resp_bits_has_data;
  input io_mem_replay_next_valid;
  input io_mem_xcpt_ma_ld;
  input io_mem_xcpt_ma_st;
  input io_mem_xcpt_pf_ld;
  input io_mem_xcpt_pf_st;
  input io_mem_ordered;
  output io_requestor_2_req_ready;
  output io_requestor_2_resp_valid;
  output io_requestor_2_resp_bits_nack;
  output io_requestor_2_resp_bits_replay;
  output io_requestor_2_resp_bits_has_data;
  output io_requestor_2_replay_next_valid;
  output io_requestor_2_xcpt_ma_ld;
  output io_requestor_2_xcpt_ma_st;
  output io_requestor_2_xcpt_pf_ld;
  output io_requestor_2_xcpt_pf_st;
  output io_requestor_2_ordered;
  output io_requestor_1_req_ready;
  output io_requestor_1_resp_valid;
  output io_requestor_1_resp_bits_nack;
  output io_requestor_1_resp_bits_replay;
  output io_requestor_1_resp_bits_has_data;
  output io_requestor_1_replay_next_valid;
  output io_requestor_1_xcpt_ma_ld;
  output io_requestor_1_xcpt_ma_st;
  output io_requestor_1_xcpt_pf_ld;
  output io_requestor_1_xcpt_pf_st;
  output io_requestor_1_ordered;
  output io_requestor_0_req_ready;
  output io_requestor_0_resp_valid;
  output io_requestor_0_resp_bits_nack;
  output io_requestor_0_resp_bits_replay;
  output io_requestor_0_resp_bits_has_data;
  output io_requestor_0_replay_next_valid;
  output io_requestor_0_xcpt_ma_ld;
  output io_requestor_0_xcpt_ma_st;
  output io_requestor_0_xcpt_pf_ld;
  output io_requestor_0_xcpt_pf_st;
  output io_requestor_0_ordered;
  output io_mem_req_valid;
  output io_mem_req_bits_kill;
  output io_mem_req_bits_phys;
  wire [39:0] io_requestor_2_resp_bits_addr,io_requestor_1_resp_bits_addr,
  io_requestor_0_resp_bits_addr,io_mem_req_bits_addr,T16;
  wire [9:0] io_requestor_2_resp_bits_tag,io_requestor_2_replay_next_bits,
  io_requestor_1_resp_bits_tag,io_requestor_1_replay_next_bits,io_requestor_0_resp_bits_tag,
  io_requestor_0_replay_next_bits,io_mem_req_bits_tag,T11;
  wire [4:0] io_requestor_2_resp_bits_cmd,io_requestor_1_resp_bits_cmd,
  io_requestor_0_resp_bits_cmd,io_mem_req_bits_cmd,T9;
  wire [2:0] io_requestor_2_resp_bits_typ,io_requestor_1_resp_bits_typ,
  io_requestor_0_resp_bits_typ,io_mem_req_bits_typ,T7;
  wire [63:0] io_requestor_2_resp_bits_data,io_requestor_2_resp_bits_data_word_bypass,
  io_requestor_2_resp_bits_store_data,io_requestor_1_resp_bits_data,
  io_requestor_1_resp_bits_data_word_bypass,io_requestor_1_resp_bits_store_data,
  io_requestor_0_resp_bits_data,io_requestor_0_resp_bits_data_word_bypass,
  io_requestor_0_resp_bits_store_data,io_mem_req_bits_data,T1;
  wire io_requestor_2_req_ready,io_requestor_2_resp_valid,
  io_requestor_2_resp_bits_nack,io_requestor_2_resp_bits_replay,io_requestor_2_resp_bits_has_data,
  io_requestor_2_replay_next_valid,io_requestor_2_xcpt_ma_ld,io_requestor_2_xcpt_ma_st,
  io_requestor_2_xcpt_pf_ld,io_requestor_2_xcpt_pf_st,io_requestor_2_ordered,
  io_requestor_1_req_ready,io_requestor_1_resp_valid,io_requestor_1_resp_bits_nack,
  io_requestor_1_resp_bits_replay,io_requestor_1_resp_bits_has_data,
  io_requestor_1_replay_next_valid,io_requestor_1_xcpt_ma_ld,io_requestor_1_xcpt_ma_st,
  io_requestor_1_xcpt_pf_ld,io_requestor_1_xcpt_pf_st,io_requestor_1_ordered,io_requestor_0_req_ready,
  io_requestor_0_resp_valid,io_requestor_0_resp_bits_nack,
  io_requestor_0_resp_bits_replay,io_requestor_0_resp_bits_has_data,io_requestor_0_replay_next_valid,
  io_requestor_0_xcpt_ma_ld,io_requestor_0_xcpt_ma_st,io_requestor_0_xcpt_pf_ld,
  io_requestor_0_xcpt_pf_st,io_requestor_0_ordered,io_mem_req_valid,io_mem_req_bits_kill,
  io_mem_req_bits_phys,N0,N1,N2,N3,N4,N5,N6,N7,io_mem_req_ready,
  io_mem_resp_bits_has_data,io_mem_xcpt_ma_ld,io_mem_xcpt_ma_st,io_mem_xcpt_pf_ld,io_mem_xcpt_pf_st,
  io_mem_ordered,N8,N9,T3,T5,N10,N11,T18,T40,T52,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27;
  reg r_valid_1,r_valid_0;
  assign io_requestor_2_resp_bits_tag[8] = 1'b0;
  assign io_requestor_2_resp_bits_tag[9] = 1'b0;
  assign io_requestor_2_replay_next_bits[8] = 1'b0;
  assign io_requestor_2_replay_next_bits[9] = 1'b0;
  assign io_requestor_1_resp_bits_tag[8] = 1'b0;
  assign io_requestor_1_resp_bits_tag[9] = 1'b0;
  assign io_requestor_1_replay_next_bits[8] = 1'b0;
  assign io_requestor_1_replay_next_bits[9] = 1'b0;
  assign io_requestor_0_resp_bits_tag[8] = 1'b0;
  assign io_requestor_0_resp_bits_tag[9] = 1'b0;
  assign io_requestor_0_replay_next_bits[8] = 1'b0;
  assign io_requestor_0_replay_next_bits[9] = 1'b0;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_2_resp_bits_addr[39] = io_mem_resp_bits_addr[39];
  assign io_requestor_1_resp_bits_addr[39] = io_mem_resp_bits_addr[39];
  assign io_requestor_0_resp_bits_addr[39] = io_mem_resp_bits_addr[39];
  assign io_requestor_2_resp_bits_addr[38] = io_mem_resp_bits_addr[38];
  assign io_requestor_1_resp_bits_addr[38] = io_mem_resp_bits_addr[38];
  assign io_requestor_0_resp_bits_addr[38] = io_mem_resp_bits_addr[38];
  assign io_requestor_2_resp_bits_addr[37] = io_mem_resp_bits_addr[37];
  assign io_requestor_1_resp_bits_addr[37] = io_mem_resp_bits_addr[37];
  assign io_requestor_0_resp_bits_addr[37] = io_mem_resp_bits_addr[37];
  assign io_requestor_2_resp_bits_addr[36] = io_mem_resp_bits_addr[36];
  assign io_requestor_1_resp_bits_addr[36] = io_mem_resp_bits_addr[36];
  assign io_requestor_0_resp_bits_addr[36] = io_mem_resp_bits_addr[36];
  assign io_requestor_2_resp_bits_addr[35] = io_mem_resp_bits_addr[35];
  assign io_requestor_1_resp_bits_addr[35] = io_mem_resp_bits_addr[35];
  assign io_requestor_0_resp_bits_addr[35] = io_mem_resp_bits_addr[35];
  assign io_requestor_2_resp_bits_addr[34] = io_mem_resp_bits_addr[34];
  assign io_requestor_1_resp_bits_addr[34] = io_mem_resp_bits_addr[34];
  assign io_requestor_0_resp_bits_addr[34] = io_mem_resp_bits_addr[34];
  assign io_requestor_2_resp_bits_addr[33] = io_mem_resp_bits_addr[33];
  assign io_requestor_1_resp_bits_addr[33] = io_mem_resp_bits_addr[33];
  assign io_requestor_0_resp_bits_addr[33] = io_mem_resp_bits_addr[33];
  assign io_requestor_2_resp_bits_addr[32] = io_mem_resp_bits_addr[32];
  assign io_requestor_1_resp_bits_addr[32] = io_mem_resp_bits_addr[32];
  assign io_requestor_0_resp_bits_addr[32] = io_mem_resp_bits_addr[32];
  assign io_requestor_2_resp_bits_addr[31] = io_mem_resp_bits_addr[31];
  assign io_requestor_1_resp_bits_addr[31] = io_mem_resp_bits_addr[31];
  assign io_requestor_0_resp_bits_addr[31] = io_mem_resp_bits_addr[31];
  assign io_requestor_2_resp_bits_addr[30] = io_mem_resp_bits_addr[30];
  assign io_requestor_1_resp_bits_addr[30] = io_mem_resp_bits_addr[30];
  assign io_requestor_0_resp_bits_addr[30] = io_mem_resp_bits_addr[30];
  assign io_requestor_2_resp_bits_addr[29] = io_mem_resp_bits_addr[29];
  assign io_requestor_1_resp_bits_addr[29] = io_mem_resp_bits_addr[29];
  assign io_requestor_0_resp_bits_addr[29] = io_mem_resp_bits_addr[29];
  assign io_requestor_2_resp_bits_addr[28] = io_mem_resp_bits_addr[28];
  assign io_requestor_1_resp_bits_addr[28] = io_mem_resp_bits_addr[28];
  assign io_requestor_0_resp_bits_addr[28] = io_mem_resp_bits_addr[28];
  assign io_requestor_2_resp_bits_addr[27] = io_mem_resp_bits_addr[27];
  assign io_requestor_1_resp_bits_addr[27] = io_mem_resp_bits_addr[27];
  assign io_requestor_0_resp_bits_addr[27] = io_mem_resp_bits_addr[27];
  assign io_requestor_2_resp_bits_addr[26] = io_mem_resp_bits_addr[26];
  assign io_requestor_1_resp_bits_addr[26] = io_mem_resp_bits_addr[26];
  assign io_requestor_0_resp_bits_addr[26] = io_mem_resp_bits_addr[26];
  assign io_requestor_2_resp_bits_addr[25] = io_mem_resp_bits_addr[25];
  assign io_requestor_1_resp_bits_addr[25] = io_mem_resp_bits_addr[25];
  assign io_requestor_0_resp_bits_addr[25] = io_mem_resp_bits_addr[25];
  assign io_requestor_2_resp_bits_addr[24] = io_mem_resp_bits_addr[24];
  assign io_requestor_1_resp_bits_addr[24] = io_mem_resp_bits_addr[24];
  assign io_requestor_0_resp_bits_addr[24] = io_mem_resp_bits_addr[24];
  assign io_requestor_2_resp_bits_addr[23] = io_mem_resp_bits_addr[23];
  assign io_requestor_1_resp_bits_addr[23] = io_mem_resp_bits_addr[23];
  assign io_requestor_0_resp_bits_addr[23] = io_mem_resp_bits_addr[23];
  assign io_requestor_2_resp_bits_addr[22] = io_mem_resp_bits_addr[22];
  assign io_requestor_1_resp_bits_addr[22] = io_mem_resp_bits_addr[22];
  assign io_requestor_0_resp_bits_addr[22] = io_mem_resp_bits_addr[22];
  assign io_requestor_2_resp_bits_addr[21] = io_mem_resp_bits_addr[21];
  assign io_requestor_1_resp_bits_addr[21] = io_mem_resp_bits_addr[21];
  assign io_requestor_0_resp_bits_addr[21] = io_mem_resp_bits_addr[21];
  assign io_requestor_2_resp_bits_addr[20] = io_mem_resp_bits_addr[20];
  assign io_requestor_1_resp_bits_addr[20] = io_mem_resp_bits_addr[20];
  assign io_requestor_0_resp_bits_addr[20] = io_mem_resp_bits_addr[20];
  assign io_requestor_2_resp_bits_addr[19] = io_mem_resp_bits_addr[19];
  assign io_requestor_1_resp_bits_addr[19] = io_mem_resp_bits_addr[19];
  assign io_requestor_0_resp_bits_addr[19] = io_mem_resp_bits_addr[19];
  assign io_requestor_2_resp_bits_addr[18] = io_mem_resp_bits_addr[18];
  assign io_requestor_1_resp_bits_addr[18] = io_mem_resp_bits_addr[18];
  assign io_requestor_0_resp_bits_addr[18] = io_mem_resp_bits_addr[18];
  assign io_requestor_2_resp_bits_addr[17] = io_mem_resp_bits_addr[17];
  assign io_requestor_1_resp_bits_addr[17] = io_mem_resp_bits_addr[17];
  assign io_requestor_0_resp_bits_addr[17] = io_mem_resp_bits_addr[17];
  assign io_requestor_2_resp_bits_addr[16] = io_mem_resp_bits_addr[16];
  assign io_requestor_1_resp_bits_addr[16] = io_mem_resp_bits_addr[16];
  assign io_requestor_0_resp_bits_addr[16] = io_mem_resp_bits_addr[16];
  assign io_requestor_2_resp_bits_addr[15] = io_mem_resp_bits_addr[15];
  assign io_requestor_1_resp_bits_addr[15] = io_mem_resp_bits_addr[15];
  assign io_requestor_0_resp_bits_addr[15] = io_mem_resp_bits_addr[15];
  assign io_requestor_2_resp_bits_addr[14] = io_mem_resp_bits_addr[14];
  assign io_requestor_1_resp_bits_addr[14] = io_mem_resp_bits_addr[14];
  assign io_requestor_0_resp_bits_addr[14] = io_mem_resp_bits_addr[14];
  assign io_requestor_2_resp_bits_addr[13] = io_mem_resp_bits_addr[13];
  assign io_requestor_1_resp_bits_addr[13] = io_mem_resp_bits_addr[13];
  assign io_requestor_0_resp_bits_addr[13] = io_mem_resp_bits_addr[13];
  assign io_requestor_2_resp_bits_addr[12] = io_mem_resp_bits_addr[12];
  assign io_requestor_1_resp_bits_addr[12] = io_mem_resp_bits_addr[12];
  assign io_requestor_0_resp_bits_addr[12] = io_mem_resp_bits_addr[12];
  assign io_requestor_2_resp_bits_addr[11] = io_mem_resp_bits_addr[11];
  assign io_requestor_1_resp_bits_addr[11] = io_mem_resp_bits_addr[11];
  assign io_requestor_0_resp_bits_addr[11] = io_mem_resp_bits_addr[11];
  assign io_requestor_2_resp_bits_addr[10] = io_mem_resp_bits_addr[10];
  assign io_requestor_1_resp_bits_addr[10] = io_mem_resp_bits_addr[10];
  assign io_requestor_0_resp_bits_addr[10] = io_mem_resp_bits_addr[10];
  assign io_requestor_2_resp_bits_addr[9] = io_mem_resp_bits_addr[9];
  assign io_requestor_1_resp_bits_addr[9] = io_mem_resp_bits_addr[9];
  assign io_requestor_0_resp_bits_addr[9] = io_mem_resp_bits_addr[9];
  assign io_requestor_2_resp_bits_addr[8] = io_mem_resp_bits_addr[8];
  assign io_requestor_1_resp_bits_addr[8] = io_mem_resp_bits_addr[8];
  assign io_requestor_0_resp_bits_addr[8] = io_mem_resp_bits_addr[8];
  assign io_requestor_2_resp_bits_addr[7] = io_mem_resp_bits_addr[7];
  assign io_requestor_1_resp_bits_addr[7] = io_mem_resp_bits_addr[7];
  assign io_requestor_0_resp_bits_addr[7] = io_mem_resp_bits_addr[7];
  assign io_requestor_2_resp_bits_addr[6] = io_mem_resp_bits_addr[6];
  assign io_requestor_1_resp_bits_addr[6] = io_mem_resp_bits_addr[6];
  assign io_requestor_0_resp_bits_addr[6] = io_mem_resp_bits_addr[6];
  assign io_requestor_2_resp_bits_addr[5] = io_mem_resp_bits_addr[5];
  assign io_requestor_1_resp_bits_addr[5] = io_mem_resp_bits_addr[5];
  assign io_requestor_0_resp_bits_addr[5] = io_mem_resp_bits_addr[5];
  assign io_requestor_2_resp_bits_addr[4] = io_mem_resp_bits_addr[4];
  assign io_requestor_1_resp_bits_addr[4] = io_mem_resp_bits_addr[4];
  assign io_requestor_0_resp_bits_addr[4] = io_mem_resp_bits_addr[4];
  assign io_requestor_2_resp_bits_addr[3] = io_mem_resp_bits_addr[3];
  assign io_requestor_1_resp_bits_addr[3] = io_mem_resp_bits_addr[3];
  assign io_requestor_0_resp_bits_addr[3] = io_mem_resp_bits_addr[3];
  assign io_requestor_2_resp_bits_addr[2] = io_mem_resp_bits_addr[2];
  assign io_requestor_1_resp_bits_addr[2] = io_mem_resp_bits_addr[2];
  assign io_requestor_0_resp_bits_addr[2] = io_mem_resp_bits_addr[2];
  assign io_requestor_2_resp_bits_addr[1] = io_mem_resp_bits_addr[1];
  assign io_requestor_1_resp_bits_addr[1] = io_mem_resp_bits_addr[1];
  assign io_requestor_0_resp_bits_addr[1] = io_mem_resp_bits_addr[1];
  assign io_requestor_2_resp_bits_addr[0] = io_mem_resp_bits_addr[0];
  assign io_requestor_1_resp_bits_addr[0] = io_mem_resp_bits_addr[0];
  assign io_requestor_0_resp_bits_addr[0] = io_mem_resp_bits_addr[0];
  assign io_requestor_2_resp_bits_tag[7] = io_mem_resp_bits_tag[9];
  assign io_requestor_1_resp_bits_tag[7] = io_mem_resp_bits_tag[9];
  assign io_requestor_0_resp_bits_tag[7] = io_mem_resp_bits_tag[9];
  assign io_requestor_2_resp_bits_tag[6] = io_mem_resp_bits_tag[8];
  assign io_requestor_1_resp_bits_tag[6] = io_mem_resp_bits_tag[8];
  assign io_requestor_0_resp_bits_tag[6] = io_mem_resp_bits_tag[8];
  assign io_requestor_2_resp_bits_tag[5] = io_mem_resp_bits_tag[7];
  assign io_requestor_1_resp_bits_tag[5] = io_mem_resp_bits_tag[7];
  assign io_requestor_0_resp_bits_tag[5] = io_mem_resp_bits_tag[7];
  assign io_requestor_2_resp_bits_tag[4] = io_mem_resp_bits_tag[6];
  assign io_requestor_1_resp_bits_tag[4] = io_mem_resp_bits_tag[6];
  assign io_requestor_0_resp_bits_tag[4] = io_mem_resp_bits_tag[6];
  assign io_requestor_2_resp_bits_tag[3] = io_mem_resp_bits_tag[5];
  assign io_requestor_1_resp_bits_tag[3] = io_mem_resp_bits_tag[5];
  assign io_requestor_0_resp_bits_tag[3] = io_mem_resp_bits_tag[5];
  assign io_requestor_2_resp_bits_tag[2] = io_mem_resp_bits_tag[4];
  assign io_requestor_1_resp_bits_tag[2] = io_mem_resp_bits_tag[4];
  assign io_requestor_0_resp_bits_tag[2] = io_mem_resp_bits_tag[4];
  assign io_requestor_2_resp_bits_tag[1] = io_mem_resp_bits_tag[3];
  assign io_requestor_1_resp_bits_tag[1] = io_mem_resp_bits_tag[3];
  assign io_requestor_0_resp_bits_tag[1] = io_mem_resp_bits_tag[3];
  assign io_requestor_2_resp_bits_tag[0] = io_mem_resp_bits_tag[2];
  assign io_requestor_1_resp_bits_tag[0] = io_mem_resp_bits_tag[2];
  assign io_requestor_0_resp_bits_tag[0] = io_mem_resp_bits_tag[2];
  assign io_requestor_2_resp_bits_cmd[4] = io_mem_resp_bits_cmd[4];
  assign io_requestor_1_resp_bits_cmd[4] = io_mem_resp_bits_cmd[4];
  assign io_requestor_0_resp_bits_cmd[4] = io_mem_resp_bits_cmd[4];
  assign io_requestor_2_resp_bits_cmd[3] = io_mem_resp_bits_cmd[3];
  assign io_requestor_1_resp_bits_cmd[3] = io_mem_resp_bits_cmd[3];
  assign io_requestor_0_resp_bits_cmd[3] = io_mem_resp_bits_cmd[3];
  assign io_requestor_2_resp_bits_cmd[2] = io_mem_resp_bits_cmd[2];
  assign io_requestor_1_resp_bits_cmd[2] = io_mem_resp_bits_cmd[2];
  assign io_requestor_0_resp_bits_cmd[2] = io_mem_resp_bits_cmd[2];
  assign io_requestor_2_resp_bits_cmd[1] = io_mem_resp_bits_cmd[1];
  assign io_requestor_1_resp_bits_cmd[1] = io_mem_resp_bits_cmd[1];
  assign io_requestor_0_resp_bits_cmd[1] = io_mem_resp_bits_cmd[1];
  assign io_requestor_2_resp_bits_cmd[0] = io_mem_resp_bits_cmd[0];
  assign io_requestor_1_resp_bits_cmd[0] = io_mem_resp_bits_cmd[0];
  assign io_requestor_0_resp_bits_cmd[0] = io_mem_resp_bits_cmd[0];
  assign io_requestor_2_resp_bits_typ[2] = io_mem_resp_bits_typ[2];
  assign io_requestor_1_resp_bits_typ[2] = io_mem_resp_bits_typ[2];
  assign io_requestor_0_resp_bits_typ[2] = io_mem_resp_bits_typ[2];
  assign io_requestor_2_resp_bits_typ[1] = io_mem_resp_bits_typ[1];
  assign io_requestor_1_resp_bits_typ[1] = io_mem_resp_bits_typ[1];
  assign io_requestor_0_resp_bits_typ[1] = io_mem_resp_bits_typ[1];
  assign io_requestor_2_resp_bits_typ[0] = io_mem_resp_bits_typ[0];
  assign io_requestor_1_resp_bits_typ[0] = io_mem_resp_bits_typ[0];
  assign io_requestor_0_resp_bits_typ[0] = io_mem_resp_bits_typ[0];
  assign io_requestor_2_resp_bits_data[63] = io_mem_resp_bits_data[63];
  assign io_requestor_1_resp_bits_data[63] = io_mem_resp_bits_data[63];
  assign io_requestor_0_resp_bits_data[63] = io_mem_resp_bits_data[63];
  assign io_requestor_2_resp_bits_data[62] = io_mem_resp_bits_data[62];
  assign io_requestor_1_resp_bits_data[62] = io_mem_resp_bits_data[62];
  assign io_requestor_0_resp_bits_data[62] = io_mem_resp_bits_data[62];
  assign io_requestor_2_resp_bits_data[61] = io_mem_resp_bits_data[61];
  assign io_requestor_1_resp_bits_data[61] = io_mem_resp_bits_data[61];
  assign io_requestor_0_resp_bits_data[61] = io_mem_resp_bits_data[61];
  assign io_requestor_2_resp_bits_data[60] = io_mem_resp_bits_data[60];
  assign io_requestor_1_resp_bits_data[60] = io_mem_resp_bits_data[60];
  assign io_requestor_0_resp_bits_data[60] = io_mem_resp_bits_data[60];
  assign io_requestor_2_resp_bits_data[59] = io_mem_resp_bits_data[59];
  assign io_requestor_1_resp_bits_data[59] = io_mem_resp_bits_data[59];
  assign io_requestor_0_resp_bits_data[59] = io_mem_resp_bits_data[59];
  assign io_requestor_2_resp_bits_data[58] = io_mem_resp_bits_data[58];
  assign io_requestor_1_resp_bits_data[58] = io_mem_resp_bits_data[58];
  assign io_requestor_0_resp_bits_data[58] = io_mem_resp_bits_data[58];
  assign io_requestor_2_resp_bits_data[57] = io_mem_resp_bits_data[57];
  assign io_requestor_1_resp_bits_data[57] = io_mem_resp_bits_data[57];
  assign io_requestor_0_resp_bits_data[57] = io_mem_resp_bits_data[57];
  assign io_requestor_2_resp_bits_data[56] = io_mem_resp_bits_data[56];
  assign io_requestor_1_resp_bits_data[56] = io_mem_resp_bits_data[56];
  assign io_requestor_0_resp_bits_data[56] = io_mem_resp_bits_data[56];
  assign io_requestor_2_resp_bits_data[55] = io_mem_resp_bits_data[55];
  assign io_requestor_1_resp_bits_data[55] = io_mem_resp_bits_data[55];
  assign io_requestor_0_resp_bits_data[55] = io_mem_resp_bits_data[55];
  assign io_requestor_2_resp_bits_data[54] = io_mem_resp_bits_data[54];
  assign io_requestor_1_resp_bits_data[54] = io_mem_resp_bits_data[54];
  assign io_requestor_0_resp_bits_data[54] = io_mem_resp_bits_data[54];
  assign io_requestor_2_resp_bits_data[53] = io_mem_resp_bits_data[53];
  assign io_requestor_1_resp_bits_data[53] = io_mem_resp_bits_data[53];
  assign io_requestor_0_resp_bits_data[53] = io_mem_resp_bits_data[53];
  assign io_requestor_2_resp_bits_data[52] = io_mem_resp_bits_data[52];
  assign io_requestor_1_resp_bits_data[52] = io_mem_resp_bits_data[52];
  assign io_requestor_0_resp_bits_data[52] = io_mem_resp_bits_data[52];
  assign io_requestor_2_resp_bits_data[51] = io_mem_resp_bits_data[51];
  assign io_requestor_1_resp_bits_data[51] = io_mem_resp_bits_data[51];
  assign io_requestor_0_resp_bits_data[51] = io_mem_resp_bits_data[51];
  assign io_requestor_2_resp_bits_data[50] = io_mem_resp_bits_data[50];
  assign io_requestor_1_resp_bits_data[50] = io_mem_resp_bits_data[50];
  assign io_requestor_0_resp_bits_data[50] = io_mem_resp_bits_data[50];
  assign io_requestor_2_resp_bits_data[49] = io_mem_resp_bits_data[49];
  assign io_requestor_1_resp_bits_data[49] = io_mem_resp_bits_data[49];
  assign io_requestor_0_resp_bits_data[49] = io_mem_resp_bits_data[49];
  assign io_requestor_2_resp_bits_data[48] = io_mem_resp_bits_data[48];
  assign io_requestor_1_resp_bits_data[48] = io_mem_resp_bits_data[48];
  assign io_requestor_0_resp_bits_data[48] = io_mem_resp_bits_data[48];
  assign io_requestor_2_resp_bits_data[47] = io_mem_resp_bits_data[47];
  assign io_requestor_1_resp_bits_data[47] = io_mem_resp_bits_data[47];
  assign io_requestor_0_resp_bits_data[47] = io_mem_resp_bits_data[47];
  assign io_requestor_2_resp_bits_data[46] = io_mem_resp_bits_data[46];
  assign io_requestor_1_resp_bits_data[46] = io_mem_resp_bits_data[46];
  assign io_requestor_0_resp_bits_data[46] = io_mem_resp_bits_data[46];
  assign io_requestor_2_resp_bits_data[45] = io_mem_resp_bits_data[45];
  assign io_requestor_1_resp_bits_data[45] = io_mem_resp_bits_data[45];
  assign io_requestor_0_resp_bits_data[45] = io_mem_resp_bits_data[45];
  assign io_requestor_2_resp_bits_data[44] = io_mem_resp_bits_data[44];
  assign io_requestor_1_resp_bits_data[44] = io_mem_resp_bits_data[44];
  assign io_requestor_0_resp_bits_data[44] = io_mem_resp_bits_data[44];
  assign io_requestor_2_resp_bits_data[43] = io_mem_resp_bits_data[43];
  assign io_requestor_1_resp_bits_data[43] = io_mem_resp_bits_data[43];
  assign io_requestor_0_resp_bits_data[43] = io_mem_resp_bits_data[43];
  assign io_requestor_2_resp_bits_data[42] = io_mem_resp_bits_data[42];
  assign io_requestor_1_resp_bits_data[42] = io_mem_resp_bits_data[42];
  assign io_requestor_0_resp_bits_data[42] = io_mem_resp_bits_data[42];
  assign io_requestor_2_resp_bits_data[41] = io_mem_resp_bits_data[41];
  assign io_requestor_1_resp_bits_data[41] = io_mem_resp_bits_data[41];
  assign io_requestor_0_resp_bits_data[41] = io_mem_resp_bits_data[41];
  assign io_requestor_2_resp_bits_data[40] = io_mem_resp_bits_data[40];
  assign io_requestor_1_resp_bits_data[40] = io_mem_resp_bits_data[40];
  assign io_requestor_0_resp_bits_data[40] = io_mem_resp_bits_data[40];
  assign io_requestor_2_resp_bits_data[39] = io_mem_resp_bits_data[39];
  assign io_requestor_1_resp_bits_data[39] = io_mem_resp_bits_data[39];
  assign io_requestor_0_resp_bits_data[39] = io_mem_resp_bits_data[39];
  assign io_requestor_2_resp_bits_data[38] = io_mem_resp_bits_data[38];
  assign io_requestor_1_resp_bits_data[38] = io_mem_resp_bits_data[38];
  assign io_requestor_0_resp_bits_data[38] = io_mem_resp_bits_data[38];
  assign io_requestor_2_resp_bits_data[37] = io_mem_resp_bits_data[37];
  assign io_requestor_1_resp_bits_data[37] = io_mem_resp_bits_data[37];
  assign io_requestor_0_resp_bits_data[37] = io_mem_resp_bits_data[37];
  assign io_requestor_2_resp_bits_data[36] = io_mem_resp_bits_data[36];
  assign io_requestor_1_resp_bits_data[36] = io_mem_resp_bits_data[36];
  assign io_requestor_0_resp_bits_data[36] = io_mem_resp_bits_data[36];
  assign io_requestor_2_resp_bits_data[35] = io_mem_resp_bits_data[35];
  assign io_requestor_1_resp_bits_data[35] = io_mem_resp_bits_data[35];
  assign io_requestor_0_resp_bits_data[35] = io_mem_resp_bits_data[35];
  assign io_requestor_2_resp_bits_data[34] = io_mem_resp_bits_data[34];
  assign io_requestor_1_resp_bits_data[34] = io_mem_resp_bits_data[34];
  assign io_requestor_0_resp_bits_data[34] = io_mem_resp_bits_data[34];
  assign io_requestor_2_resp_bits_data[33] = io_mem_resp_bits_data[33];
  assign io_requestor_1_resp_bits_data[33] = io_mem_resp_bits_data[33];
  assign io_requestor_0_resp_bits_data[33] = io_mem_resp_bits_data[33];
  assign io_requestor_2_resp_bits_data[32] = io_mem_resp_bits_data[32];
  assign io_requestor_1_resp_bits_data[32] = io_mem_resp_bits_data[32];
  assign io_requestor_0_resp_bits_data[32] = io_mem_resp_bits_data[32];
  assign io_requestor_2_resp_bits_data[31] = io_mem_resp_bits_data[31];
  assign io_requestor_1_resp_bits_data[31] = io_mem_resp_bits_data[31];
  assign io_requestor_0_resp_bits_data[31] = io_mem_resp_bits_data[31];
  assign io_requestor_2_resp_bits_data[30] = io_mem_resp_bits_data[30];
  assign io_requestor_1_resp_bits_data[30] = io_mem_resp_bits_data[30];
  assign io_requestor_0_resp_bits_data[30] = io_mem_resp_bits_data[30];
  assign io_requestor_2_resp_bits_data[29] = io_mem_resp_bits_data[29];
  assign io_requestor_1_resp_bits_data[29] = io_mem_resp_bits_data[29];
  assign io_requestor_0_resp_bits_data[29] = io_mem_resp_bits_data[29];
  assign io_requestor_2_resp_bits_data[28] = io_mem_resp_bits_data[28];
  assign io_requestor_1_resp_bits_data[28] = io_mem_resp_bits_data[28];
  assign io_requestor_0_resp_bits_data[28] = io_mem_resp_bits_data[28];
  assign io_requestor_2_resp_bits_data[27] = io_mem_resp_bits_data[27];
  assign io_requestor_1_resp_bits_data[27] = io_mem_resp_bits_data[27];
  assign io_requestor_0_resp_bits_data[27] = io_mem_resp_bits_data[27];
  assign io_requestor_2_resp_bits_data[26] = io_mem_resp_bits_data[26];
  assign io_requestor_1_resp_bits_data[26] = io_mem_resp_bits_data[26];
  assign io_requestor_0_resp_bits_data[26] = io_mem_resp_bits_data[26];
  assign io_requestor_2_resp_bits_data[25] = io_mem_resp_bits_data[25];
  assign io_requestor_1_resp_bits_data[25] = io_mem_resp_bits_data[25];
  assign io_requestor_0_resp_bits_data[25] = io_mem_resp_bits_data[25];
  assign io_requestor_2_resp_bits_data[24] = io_mem_resp_bits_data[24];
  assign io_requestor_1_resp_bits_data[24] = io_mem_resp_bits_data[24];
  assign io_requestor_0_resp_bits_data[24] = io_mem_resp_bits_data[24];
  assign io_requestor_2_resp_bits_data[23] = io_mem_resp_bits_data[23];
  assign io_requestor_1_resp_bits_data[23] = io_mem_resp_bits_data[23];
  assign io_requestor_0_resp_bits_data[23] = io_mem_resp_bits_data[23];
  assign io_requestor_2_resp_bits_data[22] = io_mem_resp_bits_data[22];
  assign io_requestor_1_resp_bits_data[22] = io_mem_resp_bits_data[22];
  assign io_requestor_0_resp_bits_data[22] = io_mem_resp_bits_data[22];
  assign io_requestor_2_resp_bits_data[21] = io_mem_resp_bits_data[21];
  assign io_requestor_1_resp_bits_data[21] = io_mem_resp_bits_data[21];
  assign io_requestor_0_resp_bits_data[21] = io_mem_resp_bits_data[21];
  assign io_requestor_2_resp_bits_data[20] = io_mem_resp_bits_data[20];
  assign io_requestor_1_resp_bits_data[20] = io_mem_resp_bits_data[20];
  assign io_requestor_0_resp_bits_data[20] = io_mem_resp_bits_data[20];
  assign io_requestor_2_resp_bits_data[19] = io_mem_resp_bits_data[19];
  assign io_requestor_1_resp_bits_data[19] = io_mem_resp_bits_data[19];
  assign io_requestor_0_resp_bits_data[19] = io_mem_resp_bits_data[19];
  assign io_requestor_2_resp_bits_data[18] = io_mem_resp_bits_data[18];
  assign io_requestor_1_resp_bits_data[18] = io_mem_resp_bits_data[18];
  assign io_requestor_0_resp_bits_data[18] = io_mem_resp_bits_data[18];
  assign io_requestor_2_resp_bits_data[17] = io_mem_resp_bits_data[17];
  assign io_requestor_1_resp_bits_data[17] = io_mem_resp_bits_data[17];
  assign io_requestor_0_resp_bits_data[17] = io_mem_resp_bits_data[17];
  assign io_requestor_2_resp_bits_data[16] = io_mem_resp_bits_data[16];
  assign io_requestor_1_resp_bits_data[16] = io_mem_resp_bits_data[16];
  assign io_requestor_0_resp_bits_data[16] = io_mem_resp_bits_data[16];
  assign io_requestor_2_resp_bits_data[15] = io_mem_resp_bits_data[15];
  assign io_requestor_1_resp_bits_data[15] = io_mem_resp_bits_data[15];
  assign io_requestor_0_resp_bits_data[15] = io_mem_resp_bits_data[15];
  assign io_requestor_2_resp_bits_data[14] = io_mem_resp_bits_data[14];
  assign io_requestor_1_resp_bits_data[14] = io_mem_resp_bits_data[14];
  assign io_requestor_0_resp_bits_data[14] = io_mem_resp_bits_data[14];
  assign io_requestor_2_resp_bits_data[13] = io_mem_resp_bits_data[13];
  assign io_requestor_1_resp_bits_data[13] = io_mem_resp_bits_data[13];
  assign io_requestor_0_resp_bits_data[13] = io_mem_resp_bits_data[13];
  assign io_requestor_2_resp_bits_data[12] = io_mem_resp_bits_data[12];
  assign io_requestor_1_resp_bits_data[12] = io_mem_resp_bits_data[12];
  assign io_requestor_0_resp_bits_data[12] = io_mem_resp_bits_data[12];
  assign io_requestor_2_resp_bits_data[11] = io_mem_resp_bits_data[11];
  assign io_requestor_1_resp_bits_data[11] = io_mem_resp_bits_data[11];
  assign io_requestor_0_resp_bits_data[11] = io_mem_resp_bits_data[11];
  assign io_requestor_2_resp_bits_data[10] = io_mem_resp_bits_data[10];
  assign io_requestor_1_resp_bits_data[10] = io_mem_resp_bits_data[10];
  assign io_requestor_0_resp_bits_data[10] = io_mem_resp_bits_data[10];
  assign io_requestor_2_resp_bits_data[9] = io_mem_resp_bits_data[9];
  assign io_requestor_1_resp_bits_data[9] = io_mem_resp_bits_data[9];
  assign io_requestor_0_resp_bits_data[9] = io_mem_resp_bits_data[9];
  assign io_requestor_2_resp_bits_data[8] = io_mem_resp_bits_data[8];
  assign io_requestor_1_resp_bits_data[8] = io_mem_resp_bits_data[8];
  assign io_requestor_0_resp_bits_data[8] = io_mem_resp_bits_data[8];
  assign io_requestor_2_resp_bits_data[7] = io_mem_resp_bits_data[7];
  assign io_requestor_1_resp_bits_data[7] = io_mem_resp_bits_data[7];
  assign io_requestor_0_resp_bits_data[7] = io_mem_resp_bits_data[7];
  assign io_requestor_2_resp_bits_data[6] = io_mem_resp_bits_data[6];
  assign io_requestor_1_resp_bits_data[6] = io_mem_resp_bits_data[6];
  assign io_requestor_0_resp_bits_data[6] = io_mem_resp_bits_data[6];
  assign io_requestor_2_resp_bits_data[5] = io_mem_resp_bits_data[5];
  assign io_requestor_1_resp_bits_data[5] = io_mem_resp_bits_data[5];
  assign io_requestor_0_resp_bits_data[5] = io_mem_resp_bits_data[5];
  assign io_requestor_2_resp_bits_data[4] = io_mem_resp_bits_data[4];
  assign io_requestor_1_resp_bits_data[4] = io_mem_resp_bits_data[4];
  assign io_requestor_0_resp_bits_data[4] = io_mem_resp_bits_data[4];
  assign io_requestor_2_resp_bits_data[3] = io_mem_resp_bits_data[3];
  assign io_requestor_1_resp_bits_data[3] = io_mem_resp_bits_data[3];
  assign io_requestor_0_resp_bits_data[3] = io_mem_resp_bits_data[3];
  assign io_requestor_2_resp_bits_data[2] = io_mem_resp_bits_data[2];
  assign io_requestor_1_resp_bits_data[2] = io_mem_resp_bits_data[2];
  assign io_requestor_0_resp_bits_data[2] = io_mem_resp_bits_data[2];
  assign io_requestor_2_resp_bits_data[1] = io_mem_resp_bits_data[1];
  assign io_requestor_1_resp_bits_data[1] = io_mem_resp_bits_data[1];
  assign io_requestor_0_resp_bits_data[1] = io_mem_resp_bits_data[1];
  assign io_requestor_2_resp_bits_data[0] = io_mem_resp_bits_data[0];
  assign io_requestor_1_resp_bits_data[0] = io_mem_resp_bits_data[0];
  assign io_requestor_0_resp_bits_data[0] = io_mem_resp_bits_data[0];
  assign io_requestor_2_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_2_resp_bits_data_word_bypass[63] = io_mem_resp_bits_data_word_bypass[63];
  assign io_requestor_1_resp_bits_data_word_bypass[63] = io_mem_resp_bits_data_word_bypass[63];
  assign io_requestor_0_resp_bits_data_word_bypass[63] = io_mem_resp_bits_data_word_bypass[63];
  assign io_requestor_2_resp_bits_data_word_bypass[62] = io_mem_resp_bits_data_word_bypass[62];
  assign io_requestor_1_resp_bits_data_word_bypass[62] = io_mem_resp_bits_data_word_bypass[62];
  assign io_requestor_0_resp_bits_data_word_bypass[62] = io_mem_resp_bits_data_word_bypass[62];
  assign io_requestor_2_resp_bits_data_word_bypass[61] = io_mem_resp_bits_data_word_bypass[61];
  assign io_requestor_1_resp_bits_data_word_bypass[61] = io_mem_resp_bits_data_word_bypass[61];
  assign io_requestor_0_resp_bits_data_word_bypass[61] = io_mem_resp_bits_data_word_bypass[61];
  assign io_requestor_2_resp_bits_data_word_bypass[60] = io_mem_resp_bits_data_word_bypass[60];
  assign io_requestor_1_resp_bits_data_word_bypass[60] = io_mem_resp_bits_data_word_bypass[60];
  assign io_requestor_0_resp_bits_data_word_bypass[60] = io_mem_resp_bits_data_word_bypass[60];
  assign io_requestor_2_resp_bits_data_word_bypass[59] = io_mem_resp_bits_data_word_bypass[59];
  assign io_requestor_1_resp_bits_data_word_bypass[59] = io_mem_resp_bits_data_word_bypass[59];
  assign io_requestor_0_resp_bits_data_word_bypass[59] = io_mem_resp_bits_data_word_bypass[59];
  assign io_requestor_2_resp_bits_data_word_bypass[58] = io_mem_resp_bits_data_word_bypass[58];
  assign io_requestor_1_resp_bits_data_word_bypass[58] = io_mem_resp_bits_data_word_bypass[58];
  assign io_requestor_0_resp_bits_data_word_bypass[58] = io_mem_resp_bits_data_word_bypass[58];
  assign io_requestor_2_resp_bits_data_word_bypass[57] = io_mem_resp_bits_data_word_bypass[57];
  assign io_requestor_1_resp_bits_data_word_bypass[57] = io_mem_resp_bits_data_word_bypass[57];
  assign io_requestor_0_resp_bits_data_word_bypass[57] = io_mem_resp_bits_data_word_bypass[57];
  assign io_requestor_2_resp_bits_data_word_bypass[56] = io_mem_resp_bits_data_word_bypass[56];
  assign io_requestor_1_resp_bits_data_word_bypass[56] = io_mem_resp_bits_data_word_bypass[56];
  assign io_requestor_0_resp_bits_data_word_bypass[56] = io_mem_resp_bits_data_word_bypass[56];
  assign io_requestor_2_resp_bits_data_word_bypass[55] = io_mem_resp_bits_data_word_bypass[55];
  assign io_requestor_1_resp_bits_data_word_bypass[55] = io_mem_resp_bits_data_word_bypass[55];
  assign io_requestor_0_resp_bits_data_word_bypass[55] = io_mem_resp_bits_data_word_bypass[55];
  assign io_requestor_2_resp_bits_data_word_bypass[54] = io_mem_resp_bits_data_word_bypass[54];
  assign io_requestor_1_resp_bits_data_word_bypass[54] = io_mem_resp_bits_data_word_bypass[54];
  assign io_requestor_0_resp_bits_data_word_bypass[54] = io_mem_resp_bits_data_word_bypass[54];
  assign io_requestor_2_resp_bits_data_word_bypass[53] = io_mem_resp_bits_data_word_bypass[53];
  assign io_requestor_1_resp_bits_data_word_bypass[53] = io_mem_resp_bits_data_word_bypass[53];
  assign io_requestor_0_resp_bits_data_word_bypass[53] = io_mem_resp_bits_data_word_bypass[53];
  assign io_requestor_2_resp_bits_data_word_bypass[52] = io_mem_resp_bits_data_word_bypass[52];
  assign io_requestor_1_resp_bits_data_word_bypass[52] = io_mem_resp_bits_data_word_bypass[52];
  assign io_requestor_0_resp_bits_data_word_bypass[52] = io_mem_resp_bits_data_word_bypass[52];
  assign io_requestor_2_resp_bits_data_word_bypass[51] = io_mem_resp_bits_data_word_bypass[51];
  assign io_requestor_1_resp_bits_data_word_bypass[51] = io_mem_resp_bits_data_word_bypass[51];
  assign io_requestor_0_resp_bits_data_word_bypass[51] = io_mem_resp_bits_data_word_bypass[51];
  assign io_requestor_2_resp_bits_data_word_bypass[50] = io_mem_resp_bits_data_word_bypass[50];
  assign io_requestor_1_resp_bits_data_word_bypass[50] = io_mem_resp_bits_data_word_bypass[50];
  assign io_requestor_0_resp_bits_data_word_bypass[50] = io_mem_resp_bits_data_word_bypass[50];
  assign io_requestor_2_resp_bits_data_word_bypass[49] = io_mem_resp_bits_data_word_bypass[49];
  assign io_requestor_1_resp_bits_data_word_bypass[49] = io_mem_resp_bits_data_word_bypass[49];
  assign io_requestor_0_resp_bits_data_word_bypass[49] = io_mem_resp_bits_data_word_bypass[49];
  assign io_requestor_2_resp_bits_data_word_bypass[48] = io_mem_resp_bits_data_word_bypass[48];
  assign io_requestor_1_resp_bits_data_word_bypass[48] = io_mem_resp_bits_data_word_bypass[48];
  assign io_requestor_0_resp_bits_data_word_bypass[48] = io_mem_resp_bits_data_word_bypass[48];
  assign io_requestor_2_resp_bits_data_word_bypass[47] = io_mem_resp_bits_data_word_bypass[47];
  assign io_requestor_1_resp_bits_data_word_bypass[47] = io_mem_resp_bits_data_word_bypass[47];
  assign io_requestor_0_resp_bits_data_word_bypass[47] = io_mem_resp_bits_data_word_bypass[47];
  assign io_requestor_2_resp_bits_data_word_bypass[46] = io_mem_resp_bits_data_word_bypass[46];
  assign io_requestor_1_resp_bits_data_word_bypass[46] = io_mem_resp_bits_data_word_bypass[46];
  assign io_requestor_0_resp_bits_data_word_bypass[46] = io_mem_resp_bits_data_word_bypass[46];
  assign io_requestor_2_resp_bits_data_word_bypass[45] = io_mem_resp_bits_data_word_bypass[45];
  assign io_requestor_1_resp_bits_data_word_bypass[45] = io_mem_resp_bits_data_word_bypass[45];
  assign io_requestor_0_resp_bits_data_word_bypass[45] = io_mem_resp_bits_data_word_bypass[45];
  assign io_requestor_2_resp_bits_data_word_bypass[44] = io_mem_resp_bits_data_word_bypass[44];
  assign io_requestor_1_resp_bits_data_word_bypass[44] = io_mem_resp_bits_data_word_bypass[44];
  assign io_requestor_0_resp_bits_data_word_bypass[44] = io_mem_resp_bits_data_word_bypass[44];
  assign io_requestor_2_resp_bits_data_word_bypass[43] = io_mem_resp_bits_data_word_bypass[43];
  assign io_requestor_1_resp_bits_data_word_bypass[43] = io_mem_resp_bits_data_word_bypass[43];
  assign io_requestor_0_resp_bits_data_word_bypass[43] = io_mem_resp_bits_data_word_bypass[43];
  assign io_requestor_2_resp_bits_data_word_bypass[42] = io_mem_resp_bits_data_word_bypass[42];
  assign io_requestor_1_resp_bits_data_word_bypass[42] = io_mem_resp_bits_data_word_bypass[42];
  assign io_requestor_0_resp_bits_data_word_bypass[42] = io_mem_resp_bits_data_word_bypass[42];
  assign io_requestor_2_resp_bits_data_word_bypass[41] = io_mem_resp_bits_data_word_bypass[41];
  assign io_requestor_1_resp_bits_data_word_bypass[41] = io_mem_resp_bits_data_word_bypass[41];
  assign io_requestor_0_resp_bits_data_word_bypass[41] = io_mem_resp_bits_data_word_bypass[41];
  assign io_requestor_2_resp_bits_data_word_bypass[40] = io_mem_resp_bits_data_word_bypass[40];
  assign io_requestor_1_resp_bits_data_word_bypass[40] = io_mem_resp_bits_data_word_bypass[40];
  assign io_requestor_0_resp_bits_data_word_bypass[40] = io_mem_resp_bits_data_word_bypass[40];
  assign io_requestor_2_resp_bits_data_word_bypass[39] = io_mem_resp_bits_data_word_bypass[39];
  assign io_requestor_1_resp_bits_data_word_bypass[39] = io_mem_resp_bits_data_word_bypass[39];
  assign io_requestor_0_resp_bits_data_word_bypass[39] = io_mem_resp_bits_data_word_bypass[39];
  assign io_requestor_2_resp_bits_data_word_bypass[38] = io_mem_resp_bits_data_word_bypass[38];
  assign io_requestor_1_resp_bits_data_word_bypass[38] = io_mem_resp_bits_data_word_bypass[38];
  assign io_requestor_0_resp_bits_data_word_bypass[38] = io_mem_resp_bits_data_word_bypass[38];
  assign io_requestor_2_resp_bits_data_word_bypass[37] = io_mem_resp_bits_data_word_bypass[37];
  assign io_requestor_1_resp_bits_data_word_bypass[37] = io_mem_resp_bits_data_word_bypass[37];
  assign io_requestor_0_resp_bits_data_word_bypass[37] = io_mem_resp_bits_data_word_bypass[37];
  assign io_requestor_2_resp_bits_data_word_bypass[36] = io_mem_resp_bits_data_word_bypass[36];
  assign io_requestor_1_resp_bits_data_word_bypass[36] = io_mem_resp_bits_data_word_bypass[36];
  assign io_requestor_0_resp_bits_data_word_bypass[36] = io_mem_resp_bits_data_word_bypass[36];
  assign io_requestor_2_resp_bits_data_word_bypass[35] = io_mem_resp_bits_data_word_bypass[35];
  assign io_requestor_1_resp_bits_data_word_bypass[35] = io_mem_resp_bits_data_word_bypass[35];
  assign io_requestor_0_resp_bits_data_word_bypass[35] = io_mem_resp_bits_data_word_bypass[35];
  assign io_requestor_2_resp_bits_data_word_bypass[34] = io_mem_resp_bits_data_word_bypass[34];
  assign io_requestor_1_resp_bits_data_word_bypass[34] = io_mem_resp_bits_data_word_bypass[34];
  assign io_requestor_0_resp_bits_data_word_bypass[34] = io_mem_resp_bits_data_word_bypass[34];
  assign io_requestor_2_resp_bits_data_word_bypass[33] = io_mem_resp_bits_data_word_bypass[33];
  assign io_requestor_1_resp_bits_data_word_bypass[33] = io_mem_resp_bits_data_word_bypass[33];
  assign io_requestor_0_resp_bits_data_word_bypass[33] = io_mem_resp_bits_data_word_bypass[33];
  assign io_requestor_2_resp_bits_data_word_bypass[32] = io_mem_resp_bits_data_word_bypass[32];
  assign io_requestor_1_resp_bits_data_word_bypass[32] = io_mem_resp_bits_data_word_bypass[32];
  assign io_requestor_0_resp_bits_data_word_bypass[32] = io_mem_resp_bits_data_word_bypass[32];
  assign io_requestor_2_resp_bits_data_word_bypass[31] = io_mem_resp_bits_data_word_bypass[31];
  assign io_requestor_1_resp_bits_data_word_bypass[31] = io_mem_resp_bits_data_word_bypass[31];
  assign io_requestor_0_resp_bits_data_word_bypass[31] = io_mem_resp_bits_data_word_bypass[31];
  assign io_requestor_2_resp_bits_data_word_bypass[30] = io_mem_resp_bits_data_word_bypass[30];
  assign io_requestor_1_resp_bits_data_word_bypass[30] = io_mem_resp_bits_data_word_bypass[30];
  assign io_requestor_0_resp_bits_data_word_bypass[30] = io_mem_resp_bits_data_word_bypass[30];
  assign io_requestor_2_resp_bits_data_word_bypass[29] = io_mem_resp_bits_data_word_bypass[29];
  assign io_requestor_1_resp_bits_data_word_bypass[29] = io_mem_resp_bits_data_word_bypass[29];
  assign io_requestor_0_resp_bits_data_word_bypass[29] = io_mem_resp_bits_data_word_bypass[29];
  assign io_requestor_2_resp_bits_data_word_bypass[28] = io_mem_resp_bits_data_word_bypass[28];
  assign io_requestor_1_resp_bits_data_word_bypass[28] = io_mem_resp_bits_data_word_bypass[28];
  assign io_requestor_0_resp_bits_data_word_bypass[28] = io_mem_resp_bits_data_word_bypass[28];
  assign io_requestor_2_resp_bits_data_word_bypass[27] = io_mem_resp_bits_data_word_bypass[27];
  assign io_requestor_1_resp_bits_data_word_bypass[27] = io_mem_resp_bits_data_word_bypass[27];
  assign io_requestor_0_resp_bits_data_word_bypass[27] = io_mem_resp_bits_data_word_bypass[27];
  assign io_requestor_2_resp_bits_data_word_bypass[26] = io_mem_resp_bits_data_word_bypass[26];
  assign io_requestor_1_resp_bits_data_word_bypass[26] = io_mem_resp_bits_data_word_bypass[26];
  assign io_requestor_0_resp_bits_data_word_bypass[26] = io_mem_resp_bits_data_word_bypass[26];
  assign io_requestor_2_resp_bits_data_word_bypass[25] = io_mem_resp_bits_data_word_bypass[25];
  assign io_requestor_1_resp_bits_data_word_bypass[25] = io_mem_resp_bits_data_word_bypass[25];
  assign io_requestor_0_resp_bits_data_word_bypass[25] = io_mem_resp_bits_data_word_bypass[25];
  assign io_requestor_2_resp_bits_data_word_bypass[24] = io_mem_resp_bits_data_word_bypass[24];
  assign io_requestor_1_resp_bits_data_word_bypass[24] = io_mem_resp_bits_data_word_bypass[24];
  assign io_requestor_0_resp_bits_data_word_bypass[24] = io_mem_resp_bits_data_word_bypass[24];
  assign io_requestor_2_resp_bits_data_word_bypass[23] = io_mem_resp_bits_data_word_bypass[23];
  assign io_requestor_1_resp_bits_data_word_bypass[23] = io_mem_resp_bits_data_word_bypass[23];
  assign io_requestor_0_resp_bits_data_word_bypass[23] = io_mem_resp_bits_data_word_bypass[23];
  assign io_requestor_2_resp_bits_data_word_bypass[22] = io_mem_resp_bits_data_word_bypass[22];
  assign io_requestor_1_resp_bits_data_word_bypass[22] = io_mem_resp_bits_data_word_bypass[22];
  assign io_requestor_0_resp_bits_data_word_bypass[22] = io_mem_resp_bits_data_word_bypass[22];
  assign io_requestor_2_resp_bits_data_word_bypass[21] = io_mem_resp_bits_data_word_bypass[21];
  assign io_requestor_1_resp_bits_data_word_bypass[21] = io_mem_resp_bits_data_word_bypass[21];
  assign io_requestor_0_resp_bits_data_word_bypass[21] = io_mem_resp_bits_data_word_bypass[21];
  assign io_requestor_2_resp_bits_data_word_bypass[20] = io_mem_resp_bits_data_word_bypass[20];
  assign io_requestor_1_resp_bits_data_word_bypass[20] = io_mem_resp_bits_data_word_bypass[20];
  assign io_requestor_0_resp_bits_data_word_bypass[20] = io_mem_resp_bits_data_word_bypass[20];
  assign io_requestor_2_resp_bits_data_word_bypass[19] = io_mem_resp_bits_data_word_bypass[19];
  assign io_requestor_1_resp_bits_data_word_bypass[19] = io_mem_resp_bits_data_word_bypass[19];
  assign io_requestor_0_resp_bits_data_word_bypass[19] = io_mem_resp_bits_data_word_bypass[19];
  assign io_requestor_2_resp_bits_data_word_bypass[18] = io_mem_resp_bits_data_word_bypass[18];
  assign io_requestor_1_resp_bits_data_word_bypass[18] = io_mem_resp_bits_data_word_bypass[18];
  assign io_requestor_0_resp_bits_data_word_bypass[18] = io_mem_resp_bits_data_word_bypass[18];
  assign io_requestor_2_resp_bits_data_word_bypass[17] = io_mem_resp_bits_data_word_bypass[17];
  assign io_requestor_1_resp_bits_data_word_bypass[17] = io_mem_resp_bits_data_word_bypass[17];
  assign io_requestor_0_resp_bits_data_word_bypass[17] = io_mem_resp_bits_data_word_bypass[17];
  assign io_requestor_2_resp_bits_data_word_bypass[16] = io_mem_resp_bits_data_word_bypass[16];
  assign io_requestor_1_resp_bits_data_word_bypass[16] = io_mem_resp_bits_data_word_bypass[16];
  assign io_requestor_0_resp_bits_data_word_bypass[16] = io_mem_resp_bits_data_word_bypass[16];
  assign io_requestor_2_resp_bits_data_word_bypass[15] = io_mem_resp_bits_data_word_bypass[15];
  assign io_requestor_1_resp_bits_data_word_bypass[15] = io_mem_resp_bits_data_word_bypass[15];
  assign io_requestor_0_resp_bits_data_word_bypass[15] = io_mem_resp_bits_data_word_bypass[15];
  assign io_requestor_2_resp_bits_data_word_bypass[14] = io_mem_resp_bits_data_word_bypass[14];
  assign io_requestor_1_resp_bits_data_word_bypass[14] = io_mem_resp_bits_data_word_bypass[14];
  assign io_requestor_0_resp_bits_data_word_bypass[14] = io_mem_resp_bits_data_word_bypass[14];
  assign io_requestor_2_resp_bits_data_word_bypass[13] = io_mem_resp_bits_data_word_bypass[13];
  assign io_requestor_1_resp_bits_data_word_bypass[13] = io_mem_resp_bits_data_word_bypass[13];
  assign io_requestor_0_resp_bits_data_word_bypass[13] = io_mem_resp_bits_data_word_bypass[13];
  assign io_requestor_2_resp_bits_data_word_bypass[12] = io_mem_resp_bits_data_word_bypass[12];
  assign io_requestor_1_resp_bits_data_word_bypass[12] = io_mem_resp_bits_data_word_bypass[12];
  assign io_requestor_0_resp_bits_data_word_bypass[12] = io_mem_resp_bits_data_word_bypass[12];
  assign io_requestor_2_resp_bits_data_word_bypass[11] = io_mem_resp_bits_data_word_bypass[11];
  assign io_requestor_1_resp_bits_data_word_bypass[11] = io_mem_resp_bits_data_word_bypass[11];
  assign io_requestor_0_resp_bits_data_word_bypass[11] = io_mem_resp_bits_data_word_bypass[11];
  assign io_requestor_2_resp_bits_data_word_bypass[10] = io_mem_resp_bits_data_word_bypass[10];
  assign io_requestor_1_resp_bits_data_word_bypass[10] = io_mem_resp_bits_data_word_bypass[10];
  assign io_requestor_0_resp_bits_data_word_bypass[10] = io_mem_resp_bits_data_word_bypass[10];
  assign io_requestor_2_resp_bits_data_word_bypass[9] = io_mem_resp_bits_data_word_bypass[9];
  assign io_requestor_1_resp_bits_data_word_bypass[9] = io_mem_resp_bits_data_word_bypass[9];
  assign io_requestor_0_resp_bits_data_word_bypass[9] = io_mem_resp_bits_data_word_bypass[9];
  assign io_requestor_2_resp_bits_data_word_bypass[8] = io_mem_resp_bits_data_word_bypass[8];
  assign io_requestor_1_resp_bits_data_word_bypass[8] = io_mem_resp_bits_data_word_bypass[8];
  assign io_requestor_0_resp_bits_data_word_bypass[8] = io_mem_resp_bits_data_word_bypass[8];
  assign io_requestor_2_resp_bits_data_word_bypass[7] = io_mem_resp_bits_data_word_bypass[7];
  assign io_requestor_1_resp_bits_data_word_bypass[7] = io_mem_resp_bits_data_word_bypass[7];
  assign io_requestor_0_resp_bits_data_word_bypass[7] = io_mem_resp_bits_data_word_bypass[7];
  assign io_requestor_2_resp_bits_data_word_bypass[6] = io_mem_resp_bits_data_word_bypass[6];
  assign io_requestor_1_resp_bits_data_word_bypass[6] = io_mem_resp_bits_data_word_bypass[6];
  assign io_requestor_0_resp_bits_data_word_bypass[6] = io_mem_resp_bits_data_word_bypass[6];
  assign io_requestor_2_resp_bits_data_word_bypass[5] = io_mem_resp_bits_data_word_bypass[5];
  assign io_requestor_1_resp_bits_data_word_bypass[5] = io_mem_resp_bits_data_word_bypass[5];
  assign io_requestor_0_resp_bits_data_word_bypass[5] = io_mem_resp_bits_data_word_bypass[5];
  assign io_requestor_2_resp_bits_data_word_bypass[4] = io_mem_resp_bits_data_word_bypass[4];
  assign io_requestor_1_resp_bits_data_word_bypass[4] = io_mem_resp_bits_data_word_bypass[4];
  assign io_requestor_0_resp_bits_data_word_bypass[4] = io_mem_resp_bits_data_word_bypass[4];
  assign io_requestor_2_resp_bits_data_word_bypass[3] = io_mem_resp_bits_data_word_bypass[3];
  assign io_requestor_1_resp_bits_data_word_bypass[3] = io_mem_resp_bits_data_word_bypass[3];
  assign io_requestor_0_resp_bits_data_word_bypass[3] = io_mem_resp_bits_data_word_bypass[3];
  assign io_requestor_2_resp_bits_data_word_bypass[2] = io_mem_resp_bits_data_word_bypass[2];
  assign io_requestor_1_resp_bits_data_word_bypass[2] = io_mem_resp_bits_data_word_bypass[2];
  assign io_requestor_0_resp_bits_data_word_bypass[2] = io_mem_resp_bits_data_word_bypass[2];
  assign io_requestor_2_resp_bits_data_word_bypass[1] = io_mem_resp_bits_data_word_bypass[1];
  assign io_requestor_1_resp_bits_data_word_bypass[1] = io_mem_resp_bits_data_word_bypass[1];
  assign io_requestor_0_resp_bits_data_word_bypass[1] = io_mem_resp_bits_data_word_bypass[1];
  assign io_requestor_2_resp_bits_data_word_bypass[0] = io_mem_resp_bits_data_word_bypass[0];
  assign io_requestor_1_resp_bits_data_word_bypass[0] = io_mem_resp_bits_data_word_bypass[0];
  assign io_requestor_0_resp_bits_data_word_bypass[0] = io_mem_resp_bits_data_word_bypass[0];
  assign io_requestor_2_resp_bits_store_data[63] = io_mem_resp_bits_store_data[63];
  assign io_requestor_1_resp_bits_store_data[63] = io_mem_resp_bits_store_data[63];
  assign io_requestor_0_resp_bits_store_data[63] = io_mem_resp_bits_store_data[63];
  assign io_requestor_2_resp_bits_store_data[62] = io_mem_resp_bits_store_data[62];
  assign io_requestor_1_resp_bits_store_data[62] = io_mem_resp_bits_store_data[62];
  assign io_requestor_0_resp_bits_store_data[62] = io_mem_resp_bits_store_data[62];
  assign io_requestor_2_resp_bits_store_data[61] = io_mem_resp_bits_store_data[61];
  assign io_requestor_1_resp_bits_store_data[61] = io_mem_resp_bits_store_data[61];
  assign io_requestor_0_resp_bits_store_data[61] = io_mem_resp_bits_store_data[61];
  assign io_requestor_2_resp_bits_store_data[60] = io_mem_resp_bits_store_data[60];
  assign io_requestor_1_resp_bits_store_data[60] = io_mem_resp_bits_store_data[60];
  assign io_requestor_0_resp_bits_store_data[60] = io_mem_resp_bits_store_data[60];
  assign io_requestor_2_resp_bits_store_data[59] = io_mem_resp_bits_store_data[59];
  assign io_requestor_1_resp_bits_store_data[59] = io_mem_resp_bits_store_data[59];
  assign io_requestor_0_resp_bits_store_data[59] = io_mem_resp_bits_store_data[59];
  assign io_requestor_2_resp_bits_store_data[58] = io_mem_resp_bits_store_data[58];
  assign io_requestor_1_resp_bits_store_data[58] = io_mem_resp_bits_store_data[58];
  assign io_requestor_0_resp_bits_store_data[58] = io_mem_resp_bits_store_data[58];
  assign io_requestor_2_resp_bits_store_data[57] = io_mem_resp_bits_store_data[57];
  assign io_requestor_1_resp_bits_store_data[57] = io_mem_resp_bits_store_data[57];
  assign io_requestor_0_resp_bits_store_data[57] = io_mem_resp_bits_store_data[57];
  assign io_requestor_2_resp_bits_store_data[56] = io_mem_resp_bits_store_data[56];
  assign io_requestor_1_resp_bits_store_data[56] = io_mem_resp_bits_store_data[56];
  assign io_requestor_0_resp_bits_store_data[56] = io_mem_resp_bits_store_data[56];
  assign io_requestor_2_resp_bits_store_data[55] = io_mem_resp_bits_store_data[55];
  assign io_requestor_1_resp_bits_store_data[55] = io_mem_resp_bits_store_data[55];
  assign io_requestor_0_resp_bits_store_data[55] = io_mem_resp_bits_store_data[55];
  assign io_requestor_2_resp_bits_store_data[54] = io_mem_resp_bits_store_data[54];
  assign io_requestor_1_resp_bits_store_data[54] = io_mem_resp_bits_store_data[54];
  assign io_requestor_0_resp_bits_store_data[54] = io_mem_resp_bits_store_data[54];
  assign io_requestor_2_resp_bits_store_data[53] = io_mem_resp_bits_store_data[53];
  assign io_requestor_1_resp_bits_store_data[53] = io_mem_resp_bits_store_data[53];
  assign io_requestor_0_resp_bits_store_data[53] = io_mem_resp_bits_store_data[53];
  assign io_requestor_2_resp_bits_store_data[52] = io_mem_resp_bits_store_data[52];
  assign io_requestor_1_resp_bits_store_data[52] = io_mem_resp_bits_store_data[52];
  assign io_requestor_0_resp_bits_store_data[52] = io_mem_resp_bits_store_data[52];
  assign io_requestor_2_resp_bits_store_data[51] = io_mem_resp_bits_store_data[51];
  assign io_requestor_1_resp_bits_store_data[51] = io_mem_resp_bits_store_data[51];
  assign io_requestor_0_resp_bits_store_data[51] = io_mem_resp_bits_store_data[51];
  assign io_requestor_2_resp_bits_store_data[50] = io_mem_resp_bits_store_data[50];
  assign io_requestor_1_resp_bits_store_data[50] = io_mem_resp_bits_store_data[50];
  assign io_requestor_0_resp_bits_store_data[50] = io_mem_resp_bits_store_data[50];
  assign io_requestor_2_resp_bits_store_data[49] = io_mem_resp_bits_store_data[49];
  assign io_requestor_1_resp_bits_store_data[49] = io_mem_resp_bits_store_data[49];
  assign io_requestor_0_resp_bits_store_data[49] = io_mem_resp_bits_store_data[49];
  assign io_requestor_2_resp_bits_store_data[48] = io_mem_resp_bits_store_data[48];
  assign io_requestor_1_resp_bits_store_data[48] = io_mem_resp_bits_store_data[48];
  assign io_requestor_0_resp_bits_store_data[48] = io_mem_resp_bits_store_data[48];
  assign io_requestor_2_resp_bits_store_data[47] = io_mem_resp_bits_store_data[47];
  assign io_requestor_1_resp_bits_store_data[47] = io_mem_resp_bits_store_data[47];
  assign io_requestor_0_resp_bits_store_data[47] = io_mem_resp_bits_store_data[47];
  assign io_requestor_2_resp_bits_store_data[46] = io_mem_resp_bits_store_data[46];
  assign io_requestor_1_resp_bits_store_data[46] = io_mem_resp_bits_store_data[46];
  assign io_requestor_0_resp_bits_store_data[46] = io_mem_resp_bits_store_data[46];
  assign io_requestor_2_resp_bits_store_data[45] = io_mem_resp_bits_store_data[45];
  assign io_requestor_1_resp_bits_store_data[45] = io_mem_resp_bits_store_data[45];
  assign io_requestor_0_resp_bits_store_data[45] = io_mem_resp_bits_store_data[45];
  assign io_requestor_2_resp_bits_store_data[44] = io_mem_resp_bits_store_data[44];
  assign io_requestor_1_resp_bits_store_data[44] = io_mem_resp_bits_store_data[44];
  assign io_requestor_0_resp_bits_store_data[44] = io_mem_resp_bits_store_data[44];
  assign io_requestor_2_resp_bits_store_data[43] = io_mem_resp_bits_store_data[43];
  assign io_requestor_1_resp_bits_store_data[43] = io_mem_resp_bits_store_data[43];
  assign io_requestor_0_resp_bits_store_data[43] = io_mem_resp_bits_store_data[43];
  assign io_requestor_2_resp_bits_store_data[42] = io_mem_resp_bits_store_data[42];
  assign io_requestor_1_resp_bits_store_data[42] = io_mem_resp_bits_store_data[42];
  assign io_requestor_0_resp_bits_store_data[42] = io_mem_resp_bits_store_data[42];
  assign io_requestor_2_resp_bits_store_data[41] = io_mem_resp_bits_store_data[41];
  assign io_requestor_1_resp_bits_store_data[41] = io_mem_resp_bits_store_data[41];
  assign io_requestor_0_resp_bits_store_data[41] = io_mem_resp_bits_store_data[41];
  assign io_requestor_2_resp_bits_store_data[40] = io_mem_resp_bits_store_data[40];
  assign io_requestor_1_resp_bits_store_data[40] = io_mem_resp_bits_store_data[40];
  assign io_requestor_0_resp_bits_store_data[40] = io_mem_resp_bits_store_data[40];
  assign io_requestor_2_resp_bits_store_data[39] = io_mem_resp_bits_store_data[39];
  assign io_requestor_1_resp_bits_store_data[39] = io_mem_resp_bits_store_data[39];
  assign io_requestor_0_resp_bits_store_data[39] = io_mem_resp_bits_store_data[39];
  assign io_requestor_2_resp_bits_store_data[38] = io_mem_resp_bits_store_data[38];
  assign io_requestor_1_resp_bits_store_data[38] = io_mem_resp_bits_store_data[38];
  assign io_requestor_0_resp_bits_store_data[38] = io_mem_resp_bits_store_data[38];
  assign io_requestor_2_resp_bits_store_data[37] = io_mem_resp_bits_store_data[37];
  assign io_requestor_1_resp_bits_store_data[37] = io_mem_resp_bits_store_data[37];
  assign io_requestor_0_resp_bits_store_data[37] = io_mem_resp_bits_store_data[37];
  assign io_requestor_2_resp_bits_store_data[36] = io_mem_resp_bits_store_data[36];
  assign io_requestor_1_resp_bits_store_data[36] = io_mem_resp_bits_store_data[36];
  assign io_requestor_0_resp_bits_store_data[36] = io_mem_resp_bits_store_data[36];
  assign io_requestor_2_resp_bits_store_data[35] = io_mem_resp_bits_store_data[35];
  assign io_requestor_1_resp_bits_store_data[35] = io_mem_resp_bits_store_data[35];
  assign io_requestor_0_resp_bits_store_data[35] = io_mem_resp_bits_store_data[35];
  assign io_requestor_2_resp_bits_store_data[34] = io_mem_resp_bits_store_data[34];
  assign io_requestor_1_resp_bits_store_data[34] = io_mem_resp_bits_store_data[34];
  assign io_requestor_0_resp_bits_store_data[34] = io_mem_resp_bits_store_data[34];
  assign io_requestor_2_resp_bits_store_data[33] = io_mem_resp_bits_store_data[33];
  assign io_requestor_1_resp_bits_store_data[33] = io_mem_resp_bits_store_data[33];
  assign io_requestor_0_resp_bits_store_data[33] = io_mem_resp_bits_store_data[33];
  assign io_requestor_2_resp_bits_store_data[32] = io_mem_resp_bits_store_data[32];
  assign io_requestor_1_resp_bits_store_data[32] = io_mem_resp_bits_store_data[32];
  assign io_requestor_0_resp_bits_store_data[32] = io_mem_resp_bits_store_data[32];
  assign io_requestor_2_resp_bits_store_data[31] = io_mem_resp_bits_store_data[31];
  assign io_requestor_1_resp_bits_store_data[31] = io_mem_resp_bits_store_data[31];
  assign io_requestor_0_resp_bits_store_data[31] = io_mem_resp_bits_store_data[31];
  assign io_requestor_2_resp_bits_store_data[30] = io_mem_resp_bits_store_data[30];
  assign io_requestor_1_resp_bits_store_data[30] = io_mem_resp_bits_store_data[30];
  assign io_requestor_0_resp_bits_store_data[30] = io_mem_resp_bits_store_data[30];
  assign io_requestor_2_resp_bits_store_data[29] = io_mem_resp_bits_store_data[29];
  assign io_requestor_1_resp_bits_store_data[29] = io_mem_resp_bits_store_data[29];
  assign io_requestor_0_resp_bits_store_data[29] = io_mem_resp_bits_store_data[29];
  assign io_requestor_2_resp_bits_store_data[28] = io_mem_resp_bits_store_data[28];
  assign io_requestor_1_resp_bits_store_data[28] = io_mem_resp_bits_store_data[28];
  assign io_requestor_0_resp_bits_store_data[28] = io_mem_resp_bits_store_data[28];
  assign io_requestor_2_resp_bits_store_data[27] = io_mem_resp_bits_store_data[27];
  assign io_requestor_1_resp_bits_store_data[27] = io_mem_resp_bits_store_data[27];
  assign io_requestor_0_resp_bits_store_data[27] = io_mem_resp_bits_store_data[27];
  assign io_requestor_2_resp_bits_store_data[26] = io_mem_resp_bits_store_data[26];
  assign io_requestor_1_resp_bits_store_data[26] = io_mem_resp_bits_store_data[26];
  assign io_requestor_0_resp_bits_store_data[26] = io_mem_resp_bits_store_data[26];
  assign io_requestor_2_resp_bits_store_data[25] = io_mem_resp_bits_store_data[25];
  assign io_requestor_1_resp_bits_store_data[25] = io_mem_resp_bits_store_data[25];
  assign io_requestor_0_resp_bits_store_data[25] = io_mem_resp_bits_store_data[25];
  assign io_requestor_2_resp_bits_store_data[24] = io_mem_resp_bits_store_data[24];
  assign io_requestor_1_resp_bits_store_data[24] = io_mem_resp_bits_store_data[24];
  assign io_requestor_0_resp_bits_store_data[24] = io_mem_resp_bits_store_data[24];
  assign io_requestor_2_resp_bits_store_data[23] = io_mem_resp_bits_store_data[23];
  assign io_requestor_1_resp_bits_store_data[23] = io_mem_resp_bits_store_data[23];
  assign io_requestor_0_resp_bits_store_data[23] = io_mem_resp_bits_store_data[23];
  assign io_requestor_2_resp_bits_store_data[22] = io_mem_resp_bits_store_data[22];
  assign io_requestor_1_resp_bits_store_data[22] = io_mem_resp_bits_store_data[22];
  assign io_requestor_0_resp_bits_store_data[22] = io_mem_resp_bits_store_data[22];
  assign io_requestor_2_resp_bits_store_data[21] = io_mem_resp_bits_store_data[21];
  assign io_requestor_1_resp_bits_store_data[21] = io_mem_resp_bits_store_data[21];
  assign io_requestor_0_resp_bits_store_data[21] = io_mem_resp_bits_store_data[21];
  assign io_requestor_2_resp_bits_store_data[20] = io_mem_resp_bits_store_data[20];
  assign io_requestor_1_resp_bits_store_data[20] = io_mem_resp_bits_store_data[20];
  assign io_requestor_0_resp_bits_store_data[20] = io_mem_resp_bits_store_data[20];
  assign io_requestor_2_resp_bits_store_data[19] = io_mem_resp_bits_store_data[19];
  assign io_requestor_1_resp_bits_store_data[19] = io_mem_resp_bits_store_data[19];
  assign io_requestor_0_resp_bits_store_data[19] = io_mem_resp_bits_store_data[19];
  assign io_requestor_2_resp_bits_store_data[18] = io_mem_resp_bits_store_data[18];
  assign io_requestor_1_resp_bits_store_data[18] = io_mem_resp_bits_store_data[18];
  assign io_requestor_0_resp_bits_store_data[18] = io_mem_resp_bits_store_data[18];
  assign io_requestor_2_resp_bits_store_data[17] = io_mem_resp_bits_store_data[17];
  assign io_requestor_1_resp_bits_store_data[17] = io_mem_resp_bits_store_data[17];
  assign io_requestor_0_resp_bits_store_data[17] = io_mem_resp_bits_store_data[17];
  assign io_requestor_2_resp_bits_store_data[16] = io_mem_resp_bits_store_data[16];
  assign io_requestor_1_resp_bits_store_data[16] = io_mem_resp_bits_store_data[16];
  assign io_requestor_0_resp_bits_store_data[16] = io_mem_resp_bits_store_data[16];
  assign io_requestor_2_resp_bits_store_data[15] = io_mem_resp_bits_store_data[15];
  assign io_requestor_1_resp_bits_store_data[15] = io_mem_resp_bits_store_data[15];
  assign io_requestor_0_resp_bits_store_data[15] = io_mem_resp_bits_store_data[15];
  assign io_requestor_2_resp_bits_store_data[14] = io_mem_resp_bits_store_data[14];
  assign io_requestor_1_resp_bits_store_data[14] = io_mem_resp_bits_store_data[14];
  assign io_requestor_0_resp_bits_store_data[14] = io_mem_resp_bits_store_data[14];
  assign io_requestor_2_resp_bits_store_data[13] = io_mem_resp_bits_store_data[13];
  assign io_requestor_1_resp_bits_store_data[13] = io_mem_resp_bits_store_data[13];
  assign io_requestor_0_resp_bits_store_data[13] = io_mem_resp_bits_store_data[13];
  assign io_requestor_2_resp_bits_store_data[12] = io_mem_resp_bits_store_data[12];
  assign io_requestor_1_resp_bits_store_data[12] = io_mem_resp_bits_store_data[12];
  assign io_requestor_0_resp_bits_store_data[12] = io_mem_resp_bits_store_data[12];
  assign io_requestor_2_resp_bits_store_data[11] = io_mem_resp_bits_store_data[11];
  assign io_requestor_1_resp_bits_store_data[11] = io_mem_resp_bits_store_data[11];
  assign io_requestor_0_resp_bits_store_data[11] = io_mem_resp_bits_store_data[11];
  assign io_requestor_2_resp_bits_store_data[10] = io_mem_resp_bits_store_data[10];
  assign io_requestor_1_resp_bits_store_data[10] = io_mem_resp_bits_store_data[10];
  assign io_requestor_0_resp_bits_store_data[10] = io_mem_resp_bits_store_data[10];
  assign io_requestor_2_resp_bits_store_data[9] = io_mem_resp_bits_store_data[9];
  assign io_requestor_1_resp_bits_store_data[9] = io_mem_resp_bits_store_data[9];
  assign io_requestor_0_resp_bits_store_data[9] = io_mem_resp_bits_store_data[9];
  assign io_requestor_2_resp_bits_store_data[8] = io_mem_resp_bits_store_data[8];
  assign io_requestor_1_resp_bits_store_data[8] = io_mem_resp_bits_store_data[8];
  assign io_requestor_0_resp_bits_store_data[8] = io_mem_resp_bits_store_data[8];
  assign io_requestor_2_resp_bits_store_data[7] = io_mem_resp_bits_store_data[7];
  assign io_requestor_1_resp_bits_store_data[7] = io_mem_resp_bits_store_data[7];
  assign io_requestor_0_resp_bits_store_data[7] = io_mem_resp_bits_store_data[7];
  assign io_requestor_2_resp_bits_store_data[6] = io_mem_resp_bits_store_data[6];
  assign io_requestor_1_resp_bits_store_data[6] = io_mem_resp_bits_store_data[6];
  assign io_requestor_0_resp_bits_store_data[6] = io_mem_resp_bits_store_data[6];
  assign io_requestor_2_resp_bits_store_data[5] = io_mem_resp_bits_store_data[5];
  assign io_requestor_1_resp_bits_store_data[5] = io_mem_resp_bits_store_data[5];
  assign io_requestor_0_resp_bits_store_data[5] = io_mem_resp_bits_store_data[5];
  assign io_requestor_2_resp_bits_store_data[4] = io_mem_resp_bits_store_data[4];
  assign io_requestor_1_resp_bits_store_data[4] = io_mem_resp_bits_store_data[4];
  assign io_requestor_0_resp_bits_store_data[4] = io_mem_resp_bits_store_data[4];
  assign io_requestor_2_resp_bits_store_data[3] = io_mem_resp_bits_store_data[3];
  assign io_requestor_1_resp_bits_store_data[3] = io_mem_resp_bits_store_data[3];
  assign io_requestor_0_resp_bits_store_data[3] = io_mem_resp_bits_store_data[3];
  assign io_requestor_2_resp_bits_store_data[2] = io_mem_resp_bits_store_data[2];
  assign io_requestor_1_resp_bits_store_data[2] = io_mem_resp_bits_store_data[2];
  assign io_requestor_0_resp_bits_store_data[2] = io_mem_resp_bits_store_data[2];
  assign io_requestor_2_resp_bits_store_data[1] = io_mem_resp_bits_store_data[1];
  assign io_requestor_1_resp_bits_store_data[1] = io_mem_resp_bits_store_data[1];
  assign io_requestor_0_resp_bits_store_data[1] = io_mem_resp_bits_store_data[1];
  assign io_requestor_2_resp_bits_store_data[0] = io_mem_resp_bits_store_data[0];
  assign io_requestor_1_resp_bits_store_data[0] = io_mem_resp_bits_store_data[0];
  assign io_requestor_0_resp_bits_store_data[0] = io_mem_resp_bits_store_data[0];
  assign io_requestor_2_replay_next_bits[7] = io_mem_replay_next_bits[9];
  assign io_requestor_1_replay_next_bits[7] = io_mem_replay_next_bits[9];
  assign io_requestor_0_replay_next_bits[7] = io_mem_replay_next_bits[9];
  assign io_requestor_2_replay_next_bits[6] = io_mem_replay_next_bits[8];
  assign io_requestor_1_replay_next_bits[6] = io_mem_replay_next_bits[8];
  assign io_requestor_0_replay_next_bits[6] = io_mem_replay_next_bits[8];
  assign io_requestor_2_replay_next_bits[5] = io_mem_replay_next_bits[7];
  assign io_requestor_1_replay_next_bits[5] = io_mem_replay_next_bits[7];
  assign io_requestor_0_replay_next_bits[5] = io_mem_replay_next_bits[7];
  assign io_requestor_2_replay_next_bits[4] = io_mem_replay_next_bits[6];
  assign io_requestor_1_replay_next_bits[4] = io_mem_replay_next_bits[6];
  assign io_requestor_0_replay_next_bits[4] = io_mem_replay_next_bits[6];
  assign io_requestor_2_replay_next_bits[3] = io_mem_replay_next_bits[5];
  assign io_requestor_1_replay_next_bits[3] = io_mem_replay_next_bits[5];
  assign io_requestor_0_replay_next_bits[3] = io_mem_replay_next_bits[5];
  assign io_requestor_2_replay_next_bits[2] = io_mem_replay_next_bits[4];
  assign io_requestor_1_replay_next_bits[2] = io_mem_replay_next_bits[4];
  assign io_requestor_0_replay_next_bits[2] = io_mem_replay_next_bits[4];
  assign io_requestor_2_replay_next_bits[1] = io_mem_replay_next_bits[3];
  assign io_requestor_1_replay_next_bits[1] = io_mem_replay_next_bits[3];
  assign io_requestor_0_replay_next_bits[1] = io_mem_replay_next_bits[3];
  assign io_requestor_2_replay_next_bits[0] = io_mem_replay_next_bits[2];
  assign io_requestor_1_replay_next_bits[0] = io_mem_replay_next_bits[2];
  assign io_requestor_0_replay_next_bits[0] = io_mem_replay_next_bits[2];
  assign io_requestor_2_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_2_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_2_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_2_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_2_ordered = io_mem_ordered;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_0_ordered = io_mem_ordered;

  always @(posedge clk) begin
    if(1'b1) begin
      r_valid_1 <= io_requestor_1_req_valid;
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      r_valid_0 <= io_requestor_0_req_valid;
    end 
  end

  assign N12 = ~io_mem_resp_bits_tag[1];
  assign N13 = io_mem_resp_bits_tag[0] | N12;
  assign N14 = ~N13;
  assign N15 = ~io_mem_replay_next_bits[1];
  assign N16 = io_mem_replay_next_bits[0] | N15;
  assign N17 = ~N16;
  assign N18 = ~io_mem_resp_bits_tag[0];
  assign N19 = N18 | io_mem_resp_bits_tag[1];
  assign N20 = ~N19;
  assign N21 = ~io_mem_replay_next_bits[0];
  assign N22 = N21 | io_mem_replay_next_bits[1];
  assign N23 = ~N22;
  assign N24 = io_mem_resp_bits_tag[0] | io_mem_resp_bits_tag[1];
  assign N25 = ~N24;
  assign N26 = io_mem_replay_next_bits[0] | io_mem_replay_next_bits[1];
  assign N27 = ~N26;
  assign io_mem_req_bits_data = (N0)? io_requestor_0_req_bits_data : 
                                (N1)? T1 : 1'b0;
  assign N0 = r_valid_0;
  assign N1 = N8;
  assign T1 = (N2)? io_requestor_1_req_bits_data : 
              (N3)? io_requestor_2_req_bits_data : 1'b0;
  assign N2 = r_valid_1;
  assign N3 = N9;
  assign io_mem_req_bits_phys = (N4)? io_requestor_0_req_bits_phys : 
                                (N5)? T3 : 1'b0;
  assign N4 = io_requestor_0_req_valid;
  assign N5 = N10;
  assign T3 = (N6)? io_requestor_1_req_bits_phys : 
              (N7)? io_requestor_2_req_bits_phys : 1'b0;
  assign N6 = T11[0];
  assign N7 = T11[1];
  assign io_mem_req_bits_kill = (N0)? io_requestor_0_req_bits_kill : 
                                (N1)? T5 : 1'b0;
  assign T5 = (N2)? io_requestor_1_req_bits_kill : 
              (N3)? io_requestor_2_req_bits_kill : 1'b0;
  assign io_mem_req_bits_typ = (N4)? io_requestor_0_req_bits_typ : 
                               (N5)? T7 : 1'b0;
  assign T7 = (N6)? io_requestor_1_req_bits_typ : 
              (N7)? io_requestor_2_req_bits_typ : 1'b0;
  assign io_mem_req_bits_cmd = (N4)? io_requestor_0_req_bits_cmd : 
                               (N5)? T9 : 1'b0;
  assign T9 = (N6)? io_requestor_1_req_bits_cmd : 
              (N7)? io_requestor_2_req_bits_cmd : 1'b0;
  assign io_mem_req_bits_tag = (N4)? { io_requestor_0_req_bits_tag[7:0], 1'b0, 1'b0 } : 
                               (N5)? T11 : 1'b0;
  assign T11[9:2] = (N6)? io_requestor_1_req_bits_tag[7:0] : 
                    (N7)? io_requestor_2_req_bits_tag[7:0] : 1'b0;
  assign io_mem_req_bits_addr = (N4)? io_requestor_0_req_bits_addr : 
                                (N5)? T16 : 1'b0;
  assign T16 = (N6)? io_requestor_1_req_bits_addr : 
               (N7)? io_requestor_2_req_bits_addr : 1'b0;
  assign N8 = ~r_valid_0;
  assign N9 = ~r_valid_1;
  assign N10 = ~io_requestor_0_req_valid;
  assign N11 = ~io_requestor_1_req_valid;
  assign T11[0] = io_requestor_1_req_valid;
  assign T11[1] = N11;
  assign io_mem_req_valid = T18 | io_requestor_2_req_valid;
  assign T18 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_replay_next_valid = io_mem_replay_next_valid & N27;
  assign io_requestor_0_resp_bits_replay = io_mem_resp_bits_replay & N25;
  assign io_requestor_0_resp_bits_nack = io_mem_resp_bits_nack & N25;
  assign io_requestor_0_resp_valid = io_mem_resp_valid & N25;
  assign io_requestor_1_replay_next_valid = io_mem_replay_next_valid & N23;
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay & N20;
  assign io_requestor_1_resp_bits_nack = io_mem_resp_bits_nack & N20;
  assign io_requestor_1_resp_valid = io_mem_resp_valid & N20;
  assign io_requestor_1_req_ready = io_mem_req_ready & T40;
  assign T40 = ~io_requestor_0_req_valid;
  assign io_requestor_2_replay_next_valid = io_mem_replay_next_valid & N17;
  assign io_requestor_2_resp_bits_replay = io_mem_resp_bits_replay & N14;
  assign io_requestor_2_resp_bits_nack = io_mem_resp_bits_nack & N14;
  assign io_requestor_2_resp_valid = io_mem_resp_valid & N14;
  assign io_requestor_2_req_ready = io_requestor_1_req_ready & T52;
  assign T52 = ~io_requestor_1_req_valid;

endmodule