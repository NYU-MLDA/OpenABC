module bsg_array_concentrate_static_1b_128
(
  i,
  o
);

  input [639:0] i;
  output [511:0] o;
  wire [511:0] o;
  assign o[511] = i[639];
  assign o[510] = i[638];
  assign o[509] = i[637];
  assign o[508] = i[636];
  assign o[507] = i[635];
  assign o[506] = i[634];
  assign o[505] = i[633];
  assign o[504] = i[632];
  assign o[503] = i[631];
  assign o[502] = i[630];
  assign o[501] = i[629];
  assign o[500] = i[628];
  assign o[499] = i[627];
  assign o[498] = i[626];
  assign o[497] = i[625];
  assign o[496] = i[624];
  assign o[495] = i[623];
  assign o[494] = i[622];
  assign o[493] = i[621];
  assign o[492] = i[620];
  assign o[491] = i[619];
  assign o[490] = i[618];
  assign o[489] = i[617];
  assign o[488] = i[616];
  assign o[487] = i[615];
  assign o[486] = i[614];
  assign o[485] = i[613];
  assign o[484] = i[612];
  assign o[483] = i[611];
  assign o[482] = i[610];
  assign o[481] = i[609];
  assign o[480] = i[608];
  assign o[479] = i[607];
  assign o[478] = i[606];
  assign o[477] = i[605];
  assign o[476] = i[604];
  assign o[475] = i[603];
  assign o[474] = i[602];
  assign o[473] = i[601];
  assign o[472] = i[600];
  assign o[471] = i[599];
  assign o[470] = i[598];
  assign o[469] = i[597];
  assign o[468] = i[596];
  assign o[467] = i[595];
  assign o[466] = i[594];
  assign o[465] = i[593];
  assign o[464] = i[592];
  assign o[463] = i[591];
  assign o[462] = i[590];
  assign o[461] = i[589];
  assign o[460] = i[588];
  assign o[459] = i[587];
  assign o[458] = i[586];
  assign o[457] = i[585];
  assign o[456] = i[584];
  assign o[455] = i[583];
  assign o[454] = i[582];
  assign o[453] = i[581];
  assign o[452] = i[580];
  assign o[451] = i[579];
  assign o[450] = i[578];
  assign o[449] = i[577];
  assign o[448] = i[576];
  assign o[447] = i[575];
  assign o[446] = i[574];
  assign o[445] = i[573];
  assign o[444] = i[572];
  assign o[443] = i[571];
  assign o[442] = i[570];
  assign o[441] = i[569];
  assign o[440] = i[568];
  assign o[439] = i[567];
  assign o[438] = i[566];
  assign o[437] = i[565];
  assign o[436] = i[564];
  assign o[435] = i[563];
  assign o[434] = i[562];
  assign o[433] = i[561];
  assign o[432] = i[560];
  assign o[431] = i[559];
  assign o[430] = i[558];
  assign o[429] = i[557];
  assign o[428] = i[556];
  assign o[427] = i[555];
  assign o[426] = i[554];
  assign o[425] = i[553];
  assign o[424] = i[552];
  assign o[423] = i[551];
  assign o[422] = i[550];
  assign o[421] = i[549];
  assign o[420] = i[548];
  assign o[419] = i[547];
  assign o[418] = i[546];
  assign o[417] = i[545];
  assign o[416] = i[544];
  assign o[415] = i[543];
  assign o[414] = i[542];
  assign o[413] = i[541];
  assign o[412] = i[540];
  assign o[411] = i[539];
  assign o[410] = i[538];
  assign o[409] = i[537];
  assign o[408] = i[536];
  assign o[407] = i[535];
  assign o[406] = i[534];
  assign o[405] = i[533];
  assign o[404] = i[532];
  assign o[403] = i[531];
  assign o[402] = i[530];
  assign o[401] = i[529];
  assign o[400] = i[528];
  assign o[399] = i[527];
  assign o[398] = i[526];
  assign o[397] = i[525];
  assign o[396] = i[524];
  assign o[395] = i[523];
  assign o[394] = i[522];
  assign o[393] = i[521];
  assign o[392] = i[520];
  assign o[391] = i[519];
  assign o[390] = i[518];
  assign o[389] = i[517];
  assign o[388] = i[516];
  assign o[387] = i[515];
  assign o[386] = i[514];
  assign o[385] = i[513];
  assign o[384] = i[512];
  assign o[383] = i[511];
  assign o[382] = i[510];
  assign o[381] = i[509];
  assign o[380] = i[508];
  assign o[379] = i[507];
  assign o[378] = i[506];
  assign o[377] = i[505];
  assign o[376] = i[504];
  assign o[375] = i[503];
  assign o[374] = i[502];
  assign o[373] = i[501];
  assign o[372] = i[500];
  assign o[371] = i[499];
  assign o[370] = i[498];
  assign o[369] = i[497];
  assign o[368] = i[496];
  assign o[367] = i[495];
  assign o[366] = i[494];
  assign o[365] = i[493];
  assign o[364] = i[492];
  assign o[363] = i[491];
  assign o[362] = i[490];
  assign o[361] = i[489];
  assign o[360] = i[488];
  assign o[359] = i[487];
  assign o[358] = i[486];
  assign o[357] = i[485];
  assign o[356] = i[484];
  assign o[355] = i[483];
  assign o[354] = i[482];
  assign o[353] = i[481];
  assign o[352] = i[480];
  assign o[351] = i[479];
  assign o[350] = i[478];
  assign o[349] = i[477];
  assign o[348] = i[476];
  assign o[347] = i[475];
  assign o[346] = i[474];
  assign o[345] = i[473];
  assign o[344] = i[472];
  assign o[343] = i[471];
  assign o[342] = i[470];
  assign o[341] = i[469];
  assign o[340] = i[468];
  assign o[339] = i[467];
  assign o[338] = i[466];
  assign o[337] = i[465];
  assign o[336] = i[464];
  assign o[335] = i[463];
  assign o[334] = i[462];
  assign o[333] = i[461];
  assign o[332] = i[460];
  assign o[331] = i[459];
  assign o[330] = i[458];
  assign o[329] = i[457];
  assign o[328] = i[456];
  assign o[327] = i[455];
  assign o[326] = i[454];
  assign o[325] = i[453];
  assign o[324] = i[452];
  assign o[323] = i[451];
  assign o[322] = i[450];
  assign o[321] = i[449];
  assign o[320] = i[448];
  assign o[319] = i[447];
  assign o[318] = i[446];
  assign o[317] = i[445];
  assign o[316] = i[444];
  assign o[315] = i[443];
  assign o[314] = i[442];
  assign o[313] = i[441];
  assign o[312] = i[440];
  assign o[311] = i[439];
  assign o[310] = i[438];
  assign o[309] = i[437];
  assign o[308] = i[436];
  assign o[307] = i[435];
  assign o[306] = i[434];
  assign o[305] = i[433];
  assign o[304] = i[432];
  assign o[303] = i[431];
  assign o[302] = i[430];
  assign o[301] = i[429];
  assign o[300] = i[428];
  assign o[299] = i[427];
  assign o[298] = i[426];
  assign o[297] = i[425];
  assign o[296] = i[424];
  assign o[295] = i[423];
  assign o[294] = i[422];
  assign o[293] = i[421];
  assign o[292] = i[420];
  assign o[291] = i[419];
  assign o[290] = i[418];
  assign o[289] = i[417];
  assign o[288] = i[416];
  assign o[287] = i[415];
  assign o[286] = i[414];
  assign o[285] = i[413];
  assign o[284] = i[412];
  assign o[283] = i[411];
  assign o[282] = i[410];
  assign o[281] = i[409];
  assign o[280] = i[408];
  assign o[279] = i[407];
  assign o[278] = i[406];
  assign o[277] = i[405];
  assign o[276] = i[404];
  assign o[275] = i[403];
  assign o[274] = i[402];
  assign o[273] = i[401];
  assign o[272] = i[400];
  assign o[271] = i[399];
  assign o[270] = i[398];
  assign o[269] = i[397];
  assign o[268] = i[396];
  assign o[267] = i[395];
  assign o[266] = i[394];
  assign o[265] = i[393];
  assign o[264] = i[392];
  assign o[263] = i[391];
  assign o[262] = i[390];
  assign o[261] = i[389];
  assign o[260] = i[388];
  assign o[259] = i[387];
  assign o[258] = i[386];
  assign o[257] = i[385];
  assign o[256] = i[384];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule