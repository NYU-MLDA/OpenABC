module bsg_mem_1r1w_synth_width_p62_els_p64_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [61:0] w_data_i;
  input [5:0] r_addr_i;
  output [61:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [61:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294;
  wire [3967:0] mem;
  reg mem_3967_sv2v_reg,mem_3966_sv2v_reg,mem_3965_sv2v_reg,mem_3964_sv2v_reg,
  mem_3963_sv2v_reg,mem_3962_sv2v_reg,mem_3961_sv2v_reg,mem_3960_sv2v_reg,
  mem_3959_sv2v_reg,mem_3958_sv2v_reg,mem_3957_sv2v_reg,mem_3956_sv2v_reg,mem_3955_sv2v_reg,
  mem_3954_sv2v_reg,mem_3953_sv2v_reg,mem_3952_sv2v_reg,mem_3951_sv2v_reg,
  mem_3950_sv2v_reg,mem_3949_sv2v_reg,mem_3948_sv2v_reg,mem_3947_sv2v_reg,mem_3946_sv2v_reg,
  mem_3945_sv2v_reg,mem_3944_sv2v_reg,mem_3943_sv2v_reg,mem_3942_sv2v_reg,
  mem_3941_sv2v_reg,mem_3940_sv2v_reg,mem_3939_sv2v_reg,mem_3938_sv2v_reg,mem_3937_sv2v_reg,
  mem_3936_sv2v_reg,mem_3935_sv2v_reg,mem_3934_sv2v_reg,mem_3933_sv2v_reg,
  mem_3932_sv2v_reg,mem_3931_sv2v_reg,mem_3930_sv2v_reg,mem_3929_sv2v_reg,mem_3928_sv2v_reg,
  mem_3927_sv2v_reg,mem_3926_sv2v_reg,mem_3925_sv2v_reg,mem_3924_sv2v_reg,
  mem_3923_sv2v_reg,mem_3922_sv2v_reg,mem_3921_sv2v_reg,mem_3920_sv2v_reg,
  mem_3919_sv2v_reg,mem_3918_sv2v_reg,mem_3917_sv2v_reg,mem_3916_sv2v_reg,mem_3915_sv2v_reg,
  mem_3914_sv2v_reg,mem_3913_sv2v_reg,mem_3912_sv2v_reg,mem_3911_sv2v_reg,
  mem_3910_sv2v_reg,mem_3909_sv2v_reg,mem_3908_sv2v_reg,mem_3907_sv2v_reg,mem_3906_sv2v_reg,
  mem_3905_sv2v_reg,mem_3904_sv2v_reg,mem_3903_sv2v_reg,mem_3902_sv2v_reg,
  mem_3901_sv2v_reg,mem_3900_sv2v_reg,mem_3899_sv2v_reg,mem_3898_sv2v_reg,mem_3897_sv2v_reg,
  mem_3896_sv2v_reg,mem_3895_sv2v_reg,mem_3894_sv2v_reg,mem_3893_sv2v_reg,
  mem_3892_sv2v_reg,mem_3891_sv2v_reg,mem_3890_sv2v_reg,mem_3889_sv2v_reg,mem_3888_sv2v_reg,
  mem_3887_sv2v_reg,mem_3886_sv2v_reg,mem_3885_sv2v_reg,mem_3884_sv2v_reg,
  mem_3883_sv2v_reg,mem_3882_sv2v_reg,mem_3881_sv2v_reg,mem_3880_sv2v_reg,
  mem_3879_sv2v_reg,mem_3878_sv2v_reg,mem_3877_sv2v_reg,mem_3876_sv2v_reg,mem_3875_sv2v_reg,
  mem_3874_sv2v_reg,mem_3873_sv2v_reg,mem_3872_sv2v_reg,mem_3871_sv2v_reg,
  mem_3870_sv2v_reg,mem_3869_sv2v_reg,mem_3868_sv2v_reg,mem_3867_sv2v_reg,mem_3866_sv2v_reg,
  mem_3865_sv2v_reg,mem_3864_sv2v_reg,mem_3863_sv2v_reg,mem_3862_sv2v_reg,
  mem_3861_sv2v_reg,mem_3860_sv2v_reg,mem_3859_sv2v_reg,mem_3858_sv2v_reg,mem_3857_sv2v_reg,
  mem_3856_sv2v_reg,mem_3855_sv2v_reg,mem_3854_sv2v_reg,mem_3853_sv2v_reg,
  mem_3852_sv2v_reg,mem_3851_sv2v_reg,mem_3850_sv2v_reg,mem_3849_sv2v_reg,mem_3848_sv2v_reg,
  mem_3847_sv2v_reg,mem_3846_sv2v_reg,mem_3845_sv2v_reg,mem_3844_sv2v_reg,
  mem_3843_sv2v_reg,mem_3842_sv2v_reg,mem_3841_sv2v_reg,mem_3840_sv2v_reg,
  mem_3839_sv2v_reg,mem_3838_sv2v_reg,mem_3837_sv2v_reg,mem_3836_sv2v_reg,mem_3835_sv2v_reg,
  mem_3834_sv2v_reg,mem_3833_sv2v_reg,mem_3832_sv2v_reg,mem_3831_sv2v_reg,
  mem_3830_sv2v_reg,mem_3829_sv2v_reg,mem_3828_sv2v_reg,mem_3827_sv2v_reg,mem_3826_sv2v_reg,
  mem_3825_sv2v_reg,mem_3824_sv2v_reg,mem_3823_sv2v_reg,mem_3822_sv2v_reg,
  mem_3821_sv2v_reg,mem_3820_sv2v_reg,mem_3819_sv2v_reg,mem_3818_sv2v_reg,mem_3817_sv2v_reg,
  mem_3816_sv2v_reg,mem_3815_sv2v_reg,mem_3814_sv2v_reg,mem_3813_sv2v_reg,
  mem_3812_sv2v_reg,mem_3811_sv2v_reg,mem_3810_sv2v_reg,mem_3809_sv2v_reg,mem_3808_sv2v_reg,
  mem_3807_sv2v_reg,mem_3806_sv2v_reg,mem_3805_sv2v_reg,mem_3804_sv2v_reg,
  mem_3803_sv2v_reg,mem_3802_sv2v_reg,mem_3801_sv2v_reg,mem_3800_sv2v_reg,
  mem_3799_sv2v_reg,mem_3798_sv2v_reg,mem_3797_sv2v_reg,mem_3796_sv2v_reg,mem_3795_sv2v_reg,
  mem_3794_sv2v_reg,mem_3793_sv2v_reg,mem_3792_sv2v_reg,mem_3791_sv2v_reg,
  mem_3790_sv2v_reg,mem_3789_sv2v_reg,mem_3788_sv2v_reg,mem_3787_sv2v_reg,mem_3786_sv2v_reg,
  mem_3785_sv2v_reg,mem_3784_sv2v_reg,mem_3783_sv2v_reg,mem_3782_sv2v_reg,
  mem_3781_sv2v_reg,mem_3780_sv2v_reg,mem_3779_sv2v_reg,mem_3778_sv2v_reg,mem_3777_sv2v_reg,
  mem_3776_sv2v_reg,mem_3775_sv2v_reg,mem_3774_sv2v_reg,mem_3773_sv2v_reg,
  mem_3772_sv2v_reg,mem_3771_sv2v_reg,mem_3770_sv2v_reg,mem_3769_sv2v_reg,mem_3768_sv2v_reg,
  mem_3767_sv2v_reg,mem_3766_sv2v_reg,mem_3765_sv2v_reg,mem_3764_sv2v_reg,
  mem_3763_sv2v_reg,mem_3762_sv2v_reg,mem_3761_sv2v_reg,mem_3760_sv2v_reg,
  mem_3759_sv2v_reg,mem_3758_sv2v_reg,mem_3757_sv2v_reg,mem_3756_sv2v_reg,mem_3755_sv2v_reg,
  mem_3754_sv2v_reg,mem_3753_sv2v_reg,mem_3752_sv2v_reg,mem_3751_sv2v_reg,
  mem_3750_sv2v_reg,mem_3749_sv2v_reg,mem_3748_sv2v_reg,mem_3747_sv2v_reg,mem_3746_sv2v_reg,
  mem_3745_sv2v_reg,mem_3744_sv2v_reg,mem_3743_sv2v_reg,mem_3742_sv2v_reg,
  mem_3741_sv2v_reg,mem_3740_sv2v_reg,mem_3739_sv2v_reg,mem_3738_sv2v_reg,mem_3737_sv2v_reg,
  mem_3736_sv2v_reg,mem_3735_sv2v_reg,mem_3734_sv2v_reg,mem_3733_sv2v_reg,
  mem_3732_sv2v_reg,mem_3731_sv2v_reg,mem_3730_sv2v_reg,mem_3729_sv2v_reg,mem_3728_sv2v_reg,
  mem_3727_sv2v_reg,mem_3726_sv2v_reg,mem_3725_sv2v_reg,mem_3724_sv2v_reg,
  mem_3723_sv2v_reg,mem_3722_sv2v_reg,mem_3721_sv2v_reg,mem_3720_sv2v_reg,
  mem_3719_sv2v_reg,mem_3718_sv2v_reg,mem_3717_sv2v_reg,mem_3716_sv2v_reg,mem_3715_sv2v_reg,
  mem_3714_sv2v_reg,mem_3713_sv2v_reg,mem_3712_sv2v_reg,mem_3711_sv2v_reg,
  mem_3710_sv2v_reg,mem_3709_sv2v_reg,mem_3708_sv2v_reg,mem_3707_sv2v_reg,mem_3706_sv2v_reg,
  mem_3705_sv2v_reg,mem_3704_sv2v_reg,mem_3703_sv2v_reg,mem_3702_sv2v_reg,
  mem_3701_sv2v_reg,mem_3700_sv2v_reg,mem_3699_sv2v_reg,mem_3698_sv2v_reg,mem_3697_sv2v_reg,
  mem_3696_sv2v_reg,mem_3695_sv2v_reg,mem_3694_sv2v_reg,mem_3693_sv2v_reg,
  mem_3692_sv2v_reg,mem_3691_sv2v_reg,mem_3690_sv2v_reg,mem_3689_sv2v_reg,mem_3688_sv2v_reg,
  mem_3687_sv2v_reg,mem_3686_sv2v_reg,mem_3685_sv2v_reg,mem_3684_sv2v_reg,
  mem_3683_sv2v_reg,mem_3682_sv2v_reg,mem_3681_sv2v_reg,mem_3680_sv2v_reg,
  mem_3679_sv2v_reg,mem_3678_sv2v_reg,mem_3677_sv2v_reg,mem_3676_sv2v_reg,mem_3675_sv2v_reg,
  mem_3674_sv2v_reg,mem_3673_sv2v_reg,mem_3672_sv2v_reg,mem_3671_sv2v_reg,
  mem_3670_sv2v_reg,mem_3669_sv2v_reg,mem_3668_sv2v_reg,mem_3667_sv2v_reg,mem_3666_sv2v_reg,
  mem_3665_sv2v_reg,mem_3664_sv2v_reg,mem_3663_sv2v_reg,mem_3662_sv2v_reg,
  mem_3661_sv2v_reg,mem_3660_sv2v_reg,mem_3659_sv2v_reg,mem_3658_sv2v_reg,mem_3657_sv2v_reg,
  mem_3656_sv2v_reg,mem_3655_sv2v_reg,mem_3654_sv2v_reg,mem_3653_sv2v_reg,
  mem_3652_sv2v_reg,mem_3651_sv2v_reg,mem_3650_sv2v_reg,mem_3649_sv2v_reg,mem_3648_sv2v_reg,
  mem_3647_sv2v_reg,mem_3646_sv2v_reg,mem_3645_sv2v_reg,mem_3644_sv2v_reg,
  mem_3643_sv2v_reg,mem_3642_sv2v_reg,mem_3641_sv2v_reg,mem_3640_sv2v_reg,
  mem_3639_sv2v_reg,mem_3638_sv2v_reg,mem_3637_sv2v_reg,mem_3636_sv2v_reg,mem_3635_sv2v_reg,
  mem_3634_sv2v_reg,mem_3633_sv2v_reg,mem_3632_sv2v_reg,mem_3631_sv2v_reg,
  mem_3630_sv2v_reg,mem_3629_sv2v_reg,mem_3628_sv2v_reg,mem_3627_sv2v_reg,mem_3626_sv2v_reg,
  mem_3625_sv2v_reg,mem_3624_sv2v_reg,mem_3623_sv2v_reg,mem_3622_sv2v_reg,
  mem_3621_sv2v_reg,mem_3620_sv2v_reg,mem_3619_sv2v_reg,mem_3618_sv2v_reg,mem_3617_sv2v_reg,
  mem_3616_sv2v_reg,mem_3615_sv2v_reg,mem_3614_sv2v_reg,mem_3613_sv2v_reg,
  mem_3612_sv2v_reg,mem_3611_sv2v_reg,mem_3610_sv2v_reg,mem_3609_sv2v_reg,mem_3608_sv2v_reg,
  mem_3607_sv2v_reg,mem_3606_sv2v_reg,mem_3605_sv2v_reg,mem_3604_sv2v_reg,
  mem_3603_sv2v_reg,mem_3602_sv2v_reg,mem_3601_sv2v_reg,mem_3600_sv2v_reg,
  mem_3599_sv2v_reg,mem_3598_sv2v_reg,mem_3597_sv2v_reg,mem_3596_sv2v_reg,mem_3595_sv2v_reg,
  mem_3594_sv2v_reg,mem_3593_sv2v_reg,mem_3592_sv2v_reg,mem_3591_sv2v_reg,
  mem_3590_sv2v_reg,mem_3589_sv2v_reg,mem_3588_sv2v_reg,mem_3587_sv2v_reg,mem_3586_sv2v_reg,
  mem_3585_sv2v_reg,mem_3584_sv2v_reg,mem_3583_sv2v_reg,mem_3582_sv2v_reg,
  mem_3581_sv2v_reg,mem_3580_sv2v_reg,mem_3579_sv2v_reg,mem_3578_sv2v_reg,mem_3577_sv2v_reg,
  mem_3576_sv2v_reg,mem_3575_sv2v_reg,mem_3574_sv2v_reg,mem_3573_sv2v_reg,
  mem_3572_sv2v_reg,mem_3571_sv2v_reg,mem_3570_sv2v_reg,mem_3569_sv2v_reg,mem_3568_sv2v_reg,
  mem_3567_sv2v_reg,mem_3566_sv2v_reg,mem_3565_sv2v_reg,mem_3564_sv2v_reg,
  mem_3563_sv2v_reg,mem_3562_sv2v_reg,mem_3561_sv2v_reg,mem_3560_sv2v_reg,
  mem_3559_sv2v_reg,mem_3558_sv2v_reg,mem_3557_sv2v_reg,mem_3556_sv2v_reg,mem_3555_sv2v_reg,
  mem_3554_sv2v_reg,mem_3553_sv2v_reg,mem_3552_sv2v_reg,mem_3551_sv2v_reg,
  mem_3550_sv2v_reg,mem_3549_sv2v_reg,mem_3548_sv2v_reg,mem_3547_sv2v_reg,mem_3546_sv2v_reg,
  mem_3545_sv2v_reg,mem_3544_sv2v_reg,mem_3543_sv2v_reg,mem_3542_sv2v_reg,
  mem_3541_sv2v_reg,mem_3540_sv2v_reg,mem_3539_sv2v_reg,mem_3538_sv2v_reg,mem_3537_sv2v_reg,
  mem_3536_sv2v_reg,mem_3535_sv2v_reg,mem_3534_sv2v_reg,mem_3533_sv2v_reg,
  mem_3532_sv2v_reg,mem_3531_sv2v_reg,mem_3530_sv2v_reg,mem_3529_sv2v_reg,mem_3528_sv2v_reg,
  mem_3527_sv2v_reg,mem_3526_sv2v_reg,mem_3525_sv2v_reg,mem_3524_sv2v_reg,
  mem_3523_sv2v_reg,mem_3522_sv2v_reg,mem_3521_sv2v_reg,mem_3520_sv2v_reg,
  mem_3519_sv2v_reg,mem_3518_sv2v_reg,mem_3517_sv2v_reg,mem_3516_sv2v_reg,mem_3515_sv2v_reg,
  mem_3514_sv2v_reg,mem_3513_sv2v_reg,mem_3512_sv2v_reg,mem_3511_sv2v_reg,
  mem_3510_sv2v_reg,mem_3509_sv2v_reg,mem_3508_sv2v_reg,mem_3507_sv2v_reg,mem_3506_sv2v_reg,
  mem_3505_sv2v_reg,mem_3504_sv2v_reg,mem_3503_sv2v_reg,mem_3502_sv2v_reg,
  mem_3501_sv2v_reg,mem_3500_sv2v_reg,mem_3499_sv2v_reg,mem_3498_sv2v_reg,mem_3497_sv2v_reg,
  mem_3496_sv2v_reg,mem_3495_sv2v_reg,mem_3494_sv2v_reg,mem_3493_sv2v_reg,
  mem_3492_sv2v_reg,mem_3491_sv2v_reg,mem_3490_sv2v_reg,mem_3489_sv2v_reg,mem_3488_sv2v_reg,
  mem_3487_sv2v_reg,mem_3486_sv2v_reg,mem_3485_sv2v_reg,mem_3484_sv2v_reg,
  mem_3483_sv2v_reg,mem_3482_sv2v_reg,mem_3481_sv2v_reg,mem_3480_sv2v_reg,
  mem_3479_sv2v_reg,mem_3478_sv2v_reg,mem_3477_sv2v_reg,mem_3476_sv2v_reg,mem_3475_sv2v_reg,
  mem_3474_sv2v_reg,mem_3473_sv2v_reg,mem_3472_sv2v_reg,mem_3471_sv2v_reg,
  mem_3470_sv2v_reg,mem_3469_sv2v_reg,mem_3468_sv2v_reg,mem_3467_sv2v_reg,mem_3466_sv2v_reg,
  mem_3465_sv2v_reg,mem_3464_sv2v_reg,mem_3463_sv2v_reg,mem_3462_sv2v_reg,
  mem_3461_sv2v_reg,mem_3460_sv2v_reg,mem_3459_sv2v_reg,mem_3458_sv2v_reg,mem_3457_sv2v_reg,
  mem_3456_sv2v_reg,mem_3455_sv2v_reg,mem_3454_sv2v_reg,mem_3453_sv2v_reg,
  mem_3452_sv2v_reg,mem_3451_sv2v_reg,mem_3450_sv2v_reg,mem_3449_sv2v_reg,mem_3448_sv2v_reg,
  mem_3447_sv2v_reg,mem_3446_sv2v_reg,mem_3445_sv2v_reg,mem_3444_sv2v_reg,
  mem_3443_sv2v_reg,mem_3442_sv2v_reg,mem_3441_sv2v_reg,mem_3440_sv2v_reg,
  mem_3439_sv2v_reg,mem_3438_sv2v_reg,mem_3437_sv2v_reg,mem_3436_sv2v_reg,mem_3435_sv2v_reg,
  mem_3434_sv2v_reg,mem_3433_sv2v_reg,mem_3432_sv2v_reg,mem_3431_sv2v_reg,
  mem_3430_sv2v_reg,mem_3429_sv2v_reg,mem_3428_sv2v_reg,mem_3427_sv2v_reg,mem_3426_sv2v_reg,
  mem_3425_sv2v_reg,mem_3424_sv2v_reg,mem_3423_sv2v_reg,mem_3422_sv2v_reg,
  mem_3421_sv2v_reg,mem_3420_sv2v_reg,mem_3419_sv2v_reg,mem_3418_sv2v_reg,mem_3417_sv2v_reg,
  mem_3416_sv2v_reg,mem_3415_sv2v_reg,mem_3414_sv2v_reg,mem_3413_sv2v_reg,
  mem_3412_sv2v_reg,mem_3411_sv2v_reg,mem_3410_sv2v_reg,mem_3409_sv2v_reg,mem_3408_sv2v_reg,
  mem_3407_sv2v_reg,mem_3406_sv2v_reg,mem_3405_sv2v_reg,mem_3404_sv2v_reg,
  mem_3403_sv2v_reg,mem_3402_sv2v_reg,mem_3401_sv2v_reg,mem_3400_sv2v_reg,
  mem_3399_sv2v_reg,mem_3398_sv2v_reg,mem_3397_sv2v_reg,mem_3396_sv2v_reg,mem_3395_sv2v_reg,
  mem_3394_sv2v_reg,mem_3393_sv2v_reg,mem_3392_sv2v_reg,mem_3391_sv2v_reg,
  mem_3390_sv2v_reg,mem_3389_sv2v_reg,mem_3388_sv2v_reg,mem_3387_sv2v_reg,mem_3386_sv2v_reg,
  mem_3385_sv2v_reg,mem_3384_sv2v_reg,mem_3383_sv2v_reg,mem_3382_sv2v_reg,
  mem_3381_sv2v_reg,mem_3380_sv2v_reg,mem_3379_sv2v_reg,mem_3378_sv2v_reg,mem_3377_sv2v_reg,
  mem_3376_sv2v_reg,mem_3375_sv2v_reg,mem_3374_sv2v_reg,mem_3373_sv2v_reg,
  mem_3372_sv2v_reg,mem_3371_sv2v_reg,mem_3370_sv2v_reg,mem_3369_sv2v_reg,mem_3368_sv2v_reg,
  mem_3367_sv2v_reg,mem_3366_sv2v_reg,mem_3365_sv2v_reg,mem_3364_sv2v_reg,
  mem_3363_sv2v_reg,mem_3362_sv2v_reg,mem_3361_sv2v_reg,mem_3360_sv2v_reg,
  mem_3359_sv2v_reg,mem_3358_sv2v_reg,mem_3357_sv2v_reg,mem_3356_sv2v_reg,mem_3355_sv2v_reg,
  mem_3354_sv2v_reg,mem_3353_sv2v_reg,mem_3352_sv2v_reg,mem_3351_sv2v_reg,
  mem_3350_sv2v_reg,mem_3349_sv2v_reg,mem_3348_sv2v_reg,mem_3347_sv2v_reg,mem_3346_sv2v_reg,
  mem_3345_sv2v_reg,mem_3344_sv2v_reg,mem_3343_sv2v_reg,mem_3342_sv2v_reg,
  mem_3341_sv2v_reg,mem_3340_sv2v_reg,mem_3339_sv2v_reg,mem_3338_sv2v_reg,mem_3337_sv2v_reg,
  mem_3336_sv2v_reg,mem_3335_sv2v_reg,mem_3334_sv2v_reg,mem_3333_sv2v_reg,
  mem_3332_sv2v_reg,mem_3331_sv2v_reg,mem_3330_sv2v_reg,mem_3329_sv2v_reg,mem_3328_sv2v_reg,
  mem_3327_sv2v_reg,mem_3326_sv2v_reg,mem_3325_sv2v_reg,mem_3324_sv2v_reg,
  mem_3323_sv2v_reg,mem_3322_sv2v_reg,mem_3321_sv2v_reg,mem_3320_sv2v_reg,
  mem_3319_sv2v_reg,mem_3318_sv2v_reg,mem_3317_sv2v_reg,mem_3316_sv2v_reg,mem_3315_sv2v_reg,
  mem_3314_sv2v_reg,mem_3313_sv2v_reg,mem_3312_sv2v_reg,mem_3311_sv2v_reg,
  mem_3310_sv2v_reg,mem_3309_sv2v_reg,mem_3308_sv2v_reg,mem_3307_sv2v_reg,mem_3306_sv2v_reg,
  mem_3305_sv2v_reg,mem_3304_sv2v_reg,mem_3303_sv2v_reg,mem_3302_sv2v_reg,
  mem_3301_sv2v_reg,mem_3300_sv2v_reg,mem_3299_sv2v_reg,mem_3298_sv2v_reg,mem_3297_sv2v_reg,
  mem_3296_sv2v_reg,mem_3295_sv2v_reg,mem_3294_sv2v_reg,mem_3293_sv2v_reg,
  mem_3292_sv2v_reg,mem_3291_sv2v_reg,mem_3290_sv2v_reg,mem_3289_sv2v_reg,mem_3288_sv2v_reg,
  mem_3287_sv2v_reg,mem_3286_sv2v_reg,mem_3285_sv2v_reg,mem_3284_sv2v_reg,
  mem_3283_sv2v_reg,mem_3282_sv2v_reg,mem_3281_sv2v_reg,mem_3280_sv2v_reg,
  mem_3279_sv2v_reg,mem_3278_sv2v_reg,mem_3277_sv2v_reg,mem_3276_sv2v_reg,mem_3275_sv2v_reg,
  mem_3274_sv2v_reg,mem_3273_sv2v_reg,mem_3272_sv2v_reg,mem_3271_sv2v_reg,
  mem_3270_sv2v_reg,mem_3269_sv2v_reg,mem_3268_sv2v_reg,mem_3267_sv2v_reg,mem_3266_sv2v_reg,
  mem_3265_sv2v_reg,mem_3264_sv2v_reg,mem_3263_sv2v_reg,mem_3262_sv2v_reg,
  mem_3261_sv2v_reg,mem_3260_sv2v_reg,mem_3259_sv2v_reg,mem_3258_sv2v_reg,mem_3257_sv2v_reg,
  mem_3256_sv2v_reg,mem_3255_sv2v_reg,mem_3254_sv2v_reg,mem_3253_sv2v_reg,
  mem_3252_sv2v_reg,mem_3251_sv2v_reg,mem_3250_sv2v_reg,mem_3249_sv2v_reg,mem_3248_sv2v_reg,
  mem_3247_sv2v_reg,mem_3246_sv2v_reg,mem_3245_sv2v_reg,mem_3244_sv2v_reg,
  mem_3243_sv2v_reg,mem_3242_sv2v_reg,mem_3241_sv2v_reg,mem_3240_sv2v_reg,
  mem_3239_sv2v_reg,mem_3238_sv2v_reg,mem_3237_sv2v_reg,mem_3236_sv2v_reg,mem_3235_sv2v_reg,
  mem_3234_sv2v_reg,mem_3233_sv2v_reg,mem_3232_sv2v_reg,mem_3231_sv2v_reg,
  mem_3230_sv2v_reg,mem_3229_sv2v_reg,mem_3228_sv2v_reg,mem_3227_sv2v_reg,mem_3226_sv2v_reg,
  mem_3225_sv2v_reg,mem_3224_sv2v_reg,mem_3223_sv2v_reg,mem_3222_sv2v_reg,
  mem_3221_sv2v_reg,mem_3220_sv2v_reg,mem_3219_sv2v_reg,mem_3218_sv2v_reg,mem_3217_sv2v_reg,
  mem_3216_sv2v_reg,mem_3215_sv2v_reg,mem_3214_sv2v_reg,mem_3213_sv2v_reg,
  mem_3212_sv2v_reg,mem_3211_sv2v_reg,mem_3210_sv2v_reg,mem_3209_sv2v_reg,mem_3208_sv2v_reg,
  mem_3207_sv2v_reg,mem_3206_sv2v_reg,mem_3205_sv2v_reg,mem_3204_sv2v_reg,
  mem_3203_sv2v_reg,mem_3202_sv2v_reg,mem_3201_sv2v_reg,mem_3200_sv2v_reg,
  mem_3199_sv2v_reg,mem_3198_sv2v_reg,mem_3197_sv2v_reg,mem_3196_sv2v_reg,mem_3195_sv2v_reg,
  mem_3194_sv2v_reg,mem_3193_sv2v_reg,mem_3192_sv2v_reg,mem_3191_sv2v_reg,
  mem_3190_sv2v_reg,mem_3189_sv2v_reg,mem_3188_sv2v_reg,mem_3187_sv2v_reg,mem_3186_sv2v_reg,
  mem_3185_sv2v_reg,mem_3184_sv2v_reg,mem_3183_sv2v_reg,mem_3182_sv2v_reg,
  mem_3181_sv2v_reg,mem_3180_sv2v_reg,mem_3179_sv2v_reg,mem_3178_sv2v_reg,mem_3177_sv2v_reg,
  mem_3176_sv2v_reg,mem_3175_sv2v_reg,mem_3174_sv2v_reg,mem_3173_sv2v_reg,
  mem_3172_sv2v_reg,mem_3171_sv2v_reg,mem_3170_sv2v_reg,mem_3169_sv2v_reg,mem_3168_sv2v_reg,
  mem_3167_sv2v_reg,mem_3166_sv2v_reg,mem_3165_sv2v_reg,mem_3164_sv2v_reg,
  mem_3163_sv2v_reg,mem_3162_sv2v_reg,mem_3161_sv2v_reg,mem_3160_sv2v_reg,
  mem_3159_sv2v_reg,mem_3158_sv2v_reg,mem_3157_sv2v_reg,mem_3156_sv2v_reg,mem_3155_sv2v_reg,
  mem_3154_sv2v_reg,mem_3153_sv2v_reg,mem_3152_sv2v_reg,mem_3151_sv2v_reg,
  mem_3150_sv2v_reg,mem_3149_sv2v_reg,mem_3148_sv2v_reg,mem_3147_sv2v_reg,mem_3146_sv2v_reg,
  mem_3145_sv2v_reg,mem_3144_sv2v_reg,mem_3143_sv2v_reg,mem_3142_sv2v_reg,
  mem_3141_sv2v_reg,mem_3140_sv2v_reg,mem_3139_sv2v_reg,mem_3138_sv2v_reg,mem_3137_sv2v_reg,
  mem_3136_sv2v_reg,mem_3135_sv2v_reg,mem_3134_sv2v_reg,mem_3133_sv2v_reg,
  mem_3132_sv2v_reg,mem_3131_sv2v_reg,mem_3130_sv2v_reg,mem_3129_sv2v_reg,mem_3128_sv2v_reg,
  mem_3127_sv2v_reg,mem_3126_sv2v_reg,mem_3125_sv2v_reg,mem_3124_sv2v_reg,
  mem_3123_sv2v_reg,mem_3122_sv2v_reg,mem_3121_sv2v_reg,mem_3120_sv2v_reg,
  mem_3119_sv2v_reg,mem_3118_sv2v_reg,mem_3117_sv2v_reg,mem_3116_sv2v_reg,mem_3115_sv2v_reg,
  mem_3114_sv2v_reg,mem_3113_sv2v_reg,mem_3112_sv2v_reg,mem_3111_sv2v_reg,
  mem_3110_sv2v_reg,mem_3109_sv2v_reg,mem_3108_sv2v_reg,mem_3107_sv2v_reg,mem_3106_sv2v_reg,
  mem_3105_sv2v_reg,mem_3104_sv2v_reg,mem_3103_sv2v_reg,mem_3102_sv2v_reg,
  mem_3101_sv2v_reg,mem_3100_sv2v_reg,mem_3099_sv2v_reg,mem_3098_sv2v_reg,mem_3097_sv2v_reg,
  mem_3096_sv2v_reg,mem_3095_sv2v_reg,mem_3094_sv2v_reg,mem_3093_sv2v_reg,
  mem_3092_sv2v_reg,mem_3091_sv2v_reg,mem_3090_sv2v_reg,mem_3089_sv2v_reg,mem_3088_sv2v_reg,
  mem_3087_sv2v_reg,mem_3086_sv2v_reg,mem_3085_sv2v_reg,mem_3084_sv2v_reg,
  mem_3083_sv2v_reg,mem_3082_sv2v_reg,mem_3081_sv2v_reg,mem_3080_sv2v_reg,
  mem_3079_sv2v_reg,mem_3078_sv2v_reg,mem_3077_sv2v_reg,mem_3076_sv2v_reg,mem_3075_sv2v_reg,
  mem_3074_sv2v_reg,mem_3073_sv2v_reg,mem_3072_sv2v_reg,mem_3071_sv2v_reg,
  mem_3070_sv2v_reg,mem_3069_sv2v_reg,mem_3068_sv2v_reg,mem_3067_sv2v_reg,mem_3066_sv2v_reg,
  mem_3065_sv2v_reg,mem_3064_sv2v_reg,mem_3063_sv2v_reg,mem_3062_sv2v_reg,
  mem_3061_sv2v_reg,mem_3060_sv2v_reg,mem_3059_sv2v_reg,mem_3058_sv2v_reg,mem_3057_sv2v_reg,
  mem_3056_sv2v_reg,mem_3055_sv2v_reg,mem_3054_sv2v_reg,mem_3053_sv2v_reg,
  mem_3052_sv2v_reg,mem_3051_sv2v_reg,mem_3050_sv2v_reg,mem_3049_sv2v_reg,mem_3048_sv2v_reg,
  mem_3047_sv2v_reg,mem_3046_sv2v_reg,mem_3045_sv2v_reg,mem_3044_sv2v_reg,
  mem_3043_sv2v_reg,mem_3042_sv2v_reg,mem_3041_sv2v_reg,mem_3040_sv2v_reg,
  mem_3039_sv2v_reg,mem_3038_sv2v_reg,mem_3037_sv2v_reg,mem_3036_sv2v_reg,mem_3035_sv2v_reg,
  mem_3034_sv2v_reg,mem_3033_sv2v_reg,mem_3032_sv2v_reg,mem_3031_sv2v_reg,
  mem_3030_sv2v_reg,mem_3029_sv2v_reg,mem_3028_sv2v_reg,mem_3027_sv2v_reg,mem_3026_sv2v_reg,
  mem_3025_sv2v_reg,mem_3024_sv2v_reg,mem_3023_sv2v_reg,mem_3022_sv2v_reg,
  mem_3021_sv2v_reg,mem_3020_sv2v_reg,mem_3019_sv2v_reg,mem_3018_sv2v_reg,mem_3017_sv2v_reg,
  mem_3016_sv2v_reg,mem_3015_sv2v_reg,mem_3014_sv2v_reg,mem_3013_sv2v_reg,
  mem_3012_sv2v_reg,mem_3011_sv2v_reg,mem_3010_sv2v_reg,mem_3009_sv2v_reg,mem_3008_sv2v_reg,
  mem_3007_sv2v_reg,mem_3006_sv2v_reg,mem_3005_sv2v_reg,mem_3004_sv2v_reg,
  mem_3003_sv2v_reg,mem_3002_sv2v_reg,mem_3001_sv2v_reg,mem_3000_sv2v_reg,
  mem_2999_sv2v_reg,mem_2998_sv2v_reg,mem_2997_sv2v_reg,mem_2996_sv2v_reg,mem_2995_sv2v_reg,
  mem_2994_sv2v_reg,mem_2993_sv2v_reg,mem_2992_sv2v_reg,mem_2991_sv2v_reg,
  mem_2990_sv2v_reg,mem_2989_sv2v_reg,mem_2988_sv2v_reg,mem_2987_sv2v_reg,mem_2986_sv2v_reg,
  mem_2985_sv2v_reg,mem_2984_sv2v_reg,mem_2983_sv2v_reg,mem_2982_sv2v_reg,
  mem_2981_sv2v_reg,mem_2980_sv2v_reg,mem_2979_sv2v_reg,mem_2978_sv2v_reg,mem_2977_sv2v_reg,
  mem_2976_sv2v_reg,mem_2975_sv2v_reg,mem_2974_sv2v_reg,mem_2973_sv2v_reg,
  mem_2972_sv2v_reg,mem_2971_sv2v_reg,mem_2970_sv2v_reg,mem_2969_sv2v_reg,mem_2968_sv2v_reg,
  mem_2967_sv2v_reg,mem_2966_sv2v_reg,mem_2965_sv2v_reg,mem_2964_sv2v_reg,
  mem_2963_sv2v_reg,mem_2962_sv2v_reg,mem_2961_sv2v_reg,mem_2960_sv2v_reg,
  mem_2959_sv2v_reg,mem_2958_sv2v_reg,mem_2957_sv2v_reg,mem_2956_sv2v_reg,mem_2955_sv2v_reg,
  mem_2954_sv2v_reg,mem_2953_sv2v_reg,mem_2952_sv2v_reg,mem_2951_sv2v_reg,
  mem_2950_sv2v_reg,mem_2949_sv2v_reg,mem_2948_sv2v_reg,mem_2947_sv2v_reg,mem_2946_sv2v_reg,
  mem_2945_sv2v_reg,mem_2944_sv2v_reg,mem_2943_sv2v_reg,mem_2942_sv2v_reg,
  mem_2941_sv2v_reg,mem_2940_sv2v_reg,mem_2939_sv2v_reg,mem_2938_sv2v_reg,mem_2937_sv2v_reg,
  mem_2936_sv2v_reg,mem_2935_sv2v_reg,mem_2934_sv2v_reg,mem_2933_sv2v_reg,
  mem_2932_sv2v_reg,mem_2931_sv2v_reg,mem_2930_sv2v_reg,mem_2929_sv2v_reg,mem_2928_sv2v_reg,
  mem_2927_sv2v_reg,mem_2926_sv2v_reg,mem_2925_sv2v_reg,mem_2924_sv2v_reg,
  mem_2923_sv2v_reg,mem_2922_sv2v_reg,mem_2921_sv2v_reg,mem_2920_sv2v_reg,
  mem_2919_sv2v_reg,mem_2918_sv2v_reg,mem_2917_sv2v_reg,mem_2916_sv2v_reg,mem_2915_sv2v_reg,
  mem_2914_sv2v_reg,mem_2913_sv2v_reg,mem_2912_sv2v_reg,mem_2911_sv2v_reg,
  mem_2910_sv2v_reg,mem_2909_sv2v_reg,mem_2908_sv2v_reg,mem_2907_sv2v_reg,mem_2906_sv2v_reg,
  mem_2905_sv2v_reg,mem_2904_sv2v_reg,mem_2903_sv2v_reg,mem_2902_sv2v_reg,
  mem_2901_sv2v_reg,mem_2900_sv2v_reg,mem_2899_sv2v_reg,mem_2898_sv2v_reg,mem_2897_sv2v_reg,
  mem_2896_sv2v_reg,mem_2895_sv2v_reg,mem_2894_sv2v_reg,mem_2893_sv2v_reg,
  mem_2892_sv2v_reg,mem_2891_sv2v_reg,mem_2890_sv2v_reg,mem_2889_sv2v_reg,mem_2888_sv2v_reg,
  mem_2887_sv2v_reg,mem_2886_sv2v_reg,mem_2885_sv2v_reg,mem_2884_sv2v_reg,
  mem_2883_sv2v_reg,mem_2882_sv2v_reg,mem_2881_sv2v_reg,mem_2880_sv2v_reg,
  mem_2879_sv2v_reg,mem_2878_sv2v_reg,mem_2877_sv2v_reg,mem_2876_sv2v_reg,mem_2875_sv2v_reg,
  mem_2874_sv2v_reg,mem_2873_sv2v_reg,mem_2872_sv2v_reg,mem_2871_sv2v_reg,
  mem_2870_sv2v_reg,mem_2869_sv2v_reg,mem_2868_sv2v_reg,mem_2867_sv2v_reg,mem_2866_sv2v_reg,
  mem_2865_sv2v_reg,mem_2864_sv2v_reg,mem_2863_sv2v_reg,mem_2862_sv2v_reg,
  mem_2861_sv2v_reg,mem_2860_sv2v_reg,mem_2859_sv2v_reg,mem_2858_sv2v_reg,mem_2857_sv2v_reg,
  mem_2856_sv2v_reg,mem_2855_sv2v_reg,mem_2854_sv2v_reg,mem_2853_sv2v_reg,
  mem_2852_sv2v_reg,mem_2851_sv2v_reg,mem_2850_sv2v_reg,mem_2849_sv2v_reg,mem_2848_sv2v_reg,
  mem_2847_sv2v_reg,mem_2846_sv2v_reg,mem_2845_sv2v_reg,mem_2844_sv2v_reg,
  mem_2843_sv2v_reg,mem_2842_sv2v_reg,mem_2841_sv2v_reg,mem_2840_sv2v_reg,
  mem_2839_sv2v_reg,mem_2838_sv2v_reg,mem_2837_sv2v_reg,mem_2836_sv2v_reg,mem_2835_sv2v_reg,
  mem_2834_sv2v_reg,mem_2833_sv2v_reg,mem_2832_sv2v_reg,mem_2831_sv2v_reg,
  mem_2830_sv2v_reg,mem_2829_sv2v_reg,mem_2828_sv2v_reg,mem_2827_sv2v_reg,mem_2826_sv2v_reg,
  mem_2825_sv2v_reg,mem_2824_sv2v_reg,mem_2823_sv2v_reg,mem_2822_sv2v_reg,
  mem_2821_sv2v_reg,mem_2820_sv2v_reg,mem_2819_sv2v_reg,mem_2818_sv2v_reg,mem_2817_sv2v_reg,
  mem_2816_sv2v_reg,mem_2815_sv2v_reg,mem_2814_sv2v_reg,mem_2813_sv2v_reg,
  mem_2812_sv2v_reg,mem_2811_sv2v_reg,mem_2810_sv2v_reg,mem_2809_sv2v_reg,mem_2808_sv2v_reg,
  mem_2807_sv2v_reg,mem_2806_sv2v_reg,mem_2805_sv2v_reg,mem_2804_sv2v_reg,
  mem_2803_sv2v_reg,mem_2802_sv2v_reg,mem_2801_sv2v_reg,mem_2800_sv2v_reg,
  mem_2799_sv2v_reg,mem_2798_sv2v_reg,mem_2797_sv2v_reg,mem_2796_sv2v_reg,mem_2795_sv2v_reg,
  mem_2794_sv2v_reg,mem_2793_sv2v_reg,mem_2792_sv2v_reg,mem_2791_sv2v_reg,
  mem_2790_sv2v_reg,mem_2789_sv2v_reg,mem_2788_sv2v_reg,mem_2787_sv2v_reg,mem_2786_sv2v_reg,
  mem_2785_sv2v_reg,mem_2784_sv2v_reg,mem_2783_sv2v_reg,mem_2782_sv2v_reg,
  mem_2781_sv2v_reg,mem_2780_sv2v_reg,mem_2779_sv2v_reg,mem_2778_sv2v_reg,mem_2777_sv2v_reg,
  mem_2776_sv2v_reg,mem_2775_sv2v_reg,mem_2774_sv2v_reg,mem_2773_sv2v_reg,
  mem_2772_sv2v_reg,mem_2771_sv2v_reg,mem_2770_sv2v_reg,mem_2769_sv2v_reg,mem_2768_sv2v_reg,
  mem_2767_sv2v_reg,mem_2766_sv2v_reg,mem_2765_sv2v_reg,mem_2764_sv2v_reg,
  mem_2763_sv2v_reg,mem_2762_sv2v_reg,mem_2761_sv2v_reg,mem_2760_sv2v_reg,
  mem_2759_sv2v_reg,mem_2758_sv2v_reg,mem_2757_sv2v_reg,mem_2756_sv2v_reg,mem_2755_sv2v_reg,
  mem_2754_sv2v_reg,mem_2753_sv2v_reg,mem_2752_sv2v_reg,mem_2751_sv2v_reg,
  mem_2750_sv2v_reg,mem_2749_sv2v_reg,mem_2748_sv2v_reg,mem_2747_sv2v_reg,mem_2746_sv2v_reg,
  mem_2745_sv2v_reg,mem_2744_sv2v_reg,mem_2743_sv2v_reg,mem_2742_sv2v_reg,
  mem_2741_sv2v_reg,mem_2740_sv2v_reg,mem_2739_sv2v_reg,mem_2738_sv2v_reg,mem_2737_sv2v_reg,
  mem_2736_sv2v_reg,mem_2735_sv2v_reg,mem_2734_sv2v_reg,mem_2733_sv2v_reg,
  mem_2732_sv2v_reg,mem_2731_sv2v_reg,mem_2730_sv2v_reg,mem_2729_sv2v_reg,mem_2728_sv2v_reg,
  mem_2727_sv2v_reg,mem_2726_sv2v_reg,mem_2725_sv2v_reg,mem_2724_sv2v_reg,
  mem_2723_sv2v_reg,mem_2722_sv2v_reg,mem_2721_sv2v_reg,mem_2720_sv2v_reg,
  mem_2719_sv2v_reg,mem_2718_sv2v_reg,mem_2717_sv2v_reg,mem_2716_sv2v_reg,mem_2715_sv2v_reg,
  mem_2714_sv2v_reg,mem_2713_sv2v_reg,mem_2712_sv2v_reg,mem_2711_sv2v_reg,
  mem_2710_sv2v_reg,mem_2709_sv2v_reg,mem_2708_sv2v_reg,mem_2707_sv2v_reg,mem_2706_sv2v_reg,
  mem_2705_sv2v_reg,mem_2704_sv2v_reg,mem_2703_sv2v_reg,mem_2702_sv2v_reg,
  mem_2701_sv2v_reg,mem_2700_sv2v_reg,mem_2699_sv2v_reg,mem_2698_sv2v_reg,mem_2697_sv2v_reg,
  mem_2696_sv2v_reg,mem_2695_sv2v_reg,mem_2694_sv2v_reg,mem_2693_sv2v_reg,
  mem_2692_sv2v_reg,mem_2691_sv2v_reg,mem_2690_sv2v_reg,mem_2689_sv2v_reg,mem_2688_sv2v_reg,
  mem_2687_sv2v_reg,mem_2686_sv2v_reg,mem_2685_sv2v_reg,mem_2684_sv2v_reg,
  mem_2683_sv2v_reg,mem_2682_sv2v_reg,mem_2681_sv2v_reg,mem_2680_sv2v_reg,
  mem_2679_sv2v_reg,mem_2678_sv2v_reg,mem_2677_sv2v_reg,mem_2676_sv2v_reg,mem_2675_sv2v_reg,
  mem_2674_sv2v_reg,mem_2673_sv2v_reg,mem_2672_sv2v_reg,mem_2671_sv2v_reg,
  mem_2670_sv2v_reg,mem_2669_sv2v_reg,mem_2668_sv2v_reg,mem_2667_sv2v_reg,mem_2666_sv2v_reg,
  mem_2665_sv2v_reg,mem_2664_sv2v_reg,mem_2663_sv2v_reg,mem_2662_sv2v_reg,
  mem_2661_sv2v_reg,mem_2660_sv2v_reg,mem_2659_sv2v_reg,mem_2658_sv2v_reg,mem_2657_sv2v_reg,
  mem_2656_sv2v_reg,mem_2655_sv2v_reg,mem_2654_sv2v_reg,mem_2653_sv2v_reg,
  mem_2652_sv2v_reg,mem_2651_sv2v_reg,mem_2650_sv2v_reg,mem_2649_sv2v_reg,mem_2648_sv2v_reg,
  mem_2647_sv2v_reg,mem_2646_sv2v_reg,mem_2645_sv2v_reg,mem_2644_sv2v_reg,
  mem_2643_sv2v_reg,mem_2642_sv2v_reg,mem_2641_sv2v_reg,mem_2640_sv2v_reg,
  mem_2639_sv2v_reg,mem_2638_sv2v_reg,mem_2637_sv2v_reg,mem_2636_sv2v_reg,mem_2635_sv2v_reg,
  mem_2634_sv2v_reg,mem_2633_sv2v_reg,mem_2632_sv2v_reg,mem_2631_sv2v_reg,
  mem_2630_sv2v_reg,mem_2629_sv2v_reg,mem_2628_sv2v_reg,mem_2627_sv2v_reg,mem_2626_sv2v_reg,
  mem_2625_sv2v_reg,mem_2624_sv2v_reg,mem_2623_sv2v_reg,mem_2622_sv2v_reg,
  mem_2621_sv2v_reg,mem_2620_sv2v_reg,mem_2619_sv2v_reg,mem_2618_sv2v_reg,mem_2617_sv2v_reg,
  mem_2616_sv2v_reg,mem_2615_sv2v_reg,mem_2614_sv2v_reg,mem_2613_sv2v_reg,
  mem_2612_sv2v_reg,mem_2611_sv2v_reg,mem_2610_sv2v_reg,mem_2609_sv2v_reg,mem_2608_sv2v_reg,
  mem_2607_sv2v_reg,mem_2606_sv2v_reg,mem_2605_sv2v_reg,mem_2604_sv2v_reg,
  mem_2603_sv2v_reg,mem_2602_sv2v_reg,mem_2601_sv2v_reg,mem_2600_sv2v_reg,
  mem_2599_sv2v_reg,mem_2598_sv2v_reg,mem_2597_sv2v_reg,mem_2596_sv2v_reg,mem_2595_sv2v_reg,
  mem_2594_sv2v_reg,mem_2593_sv2v_reg,mem_2592_sv2v_reg,mem_2591_sv2v_reg,
  mem_2590_sv2v_reg,mem_2589_sv2v_reg,mem_2588_sv2v_reg,mem_2587_sv2v_reg,mem_2586_sv2v_reg,
  mem_2585_sv2v_reg,mem_2584_sv2v_reg,mem_2583_sv2v_reg,mem_2582_sv2v_reg,
  mem_2581_sv2v_reg,mem_2580_sv2v_reg,mem_2579_sv2v_reg,mem_2578_sv2v_reg,mem_2577_sv2v_reg,
  mem_2576_sv2v_reg,mem_2575_sv2v_reg,mem_2574_sv2v_reg,mem_2573_sv2v_reg,
  mem_2572_sv2v_reg,mem_2571_sv2v_reg,mem_2570_sv2v_reg,mem_2569_sv2v_reg,mem_2568_sv2v_reg,
  mem_2567_sv2v_reg,mem_2566_sv2v_reg,mem_2565_sv2v_reg,mem_2564_sv2v_reg,
  mem_2563_sv2v_reg,mem_2562_sv2v_reg,mem_2561_sv2v_reg,mem_2560_sv2v_reg,
  mem_2559_sv2v_reg,mem_2558_sv2v_reg,mem_2557_sv2v_reg,mem_2556_sv2v_reg,mem_2555_sv2v_reg,
  mem_2554_sv2v_reg,mem_2553_sv2v_reg,mem_2552_sv2v_reg,mem_2551_sv2v_reg,
  mem_2550_sv2v_reg,mem_2549_sv2v_reg,mem_2548_sv2v_reg,mem_2547_sv2v_reg,mem_2546_sv2v_reg,
  mem_2545_sv2v_reg,mem_2544_sv2v_reg,mem_2543_sv2v_reg,mem_2542_sv2v_reg,
  mem_2541_sv2v_reg,mem_2540_sv2v_reg,mem_2539_sv2v_reg,mem_2538_sv2v_reg,mem_2537_sv2v_reg,
  mem_2536_sv2v_reg,mem_2535_sv2v_reg,mem_2534_sv2v_reg,mem_2533_sv2v_reg,
  mem_2532_sv2v_reg,mem_2531_sv2v_reg,mem_2530_sv2v_reg,mem_2529_sv2v_reg,mem_2528_sv2v_reg,
  mem_2527_sv2v_reg,mem_2526_sv2v_reg,mem_2525_sv2v_reg,mem_2524_sv2v_reg,
  mem_2523_sv2v_reg,mem_2522_sv2v_reg,mem_2521_sv2v_reg,mem_2520_sv2v_reg,
  mem_2519_sv2v_reg,mem_2518_sv2v_reg,mem_2517_sv2v_reg,mem_2516_sv2v_reg,mem_2515_sv2v_reg,
  mem_2514_sv2v_reg,mem_2513_sv2v_reg,mem_2512_sv2v_reg,mem_2511_sv2v_reg,
  mem_2510_sv2v_reg,mem_2509_sv2v_reg,mem_2508_sv2v_reg,mem_2507_sv2v_reg,mem_2506_sv2v_reg,
  mem_2505_sv2v_reg,mem_2504_sv2v_reg,mem_2503_sv2v_reg,mem_2502_sv2v_reg,
  mem_2501_sv2v_reg,mem_2500_sv2v_reg,mem_2499_sv2v_reg,mem_2498_sv2v_reg,mem_2497_sv2v_reg,
  mem_2496_sv2v_reg,mem_2495_sv2v_reg,mem_2494_sv2v_reg,mem_2493_sv2v_reg,
  mem_2492_sv2v_reg,mem_2491_sv2v_reg,mem_2490_sv2v_reg,mem_2489_sv2v_reg,mem_2488_sv2v_reg,
  mem_2487_sv2v_reg,mem_2486_sv2v_reg,mem_2485_sv2v_reg,mem_2484_sv2v_reg,
  mem_2483_sv2v_reg,mem_2482_sv2v_reg,mem_2481_sv2v_reg,mem_2480_sv2v_reg,
  mem_2479_sv2v_reg,mem_2478_sv2v_reg,mem_2477_sv2v_reg,mem_2476_sv2v_reg,mem_2475_sv2v_reg,
  mem_2474_sv2v_reg,mem_2473_sv2v_reg,mem_2472_sv2v_reg,mem_2471_sv2v_reg,
  mem_2470_sv2v_reg,mem_2469_sv2v_reg,mem_2468_sv2v_reg,mem_2467_sv2v_reg,mem_2466_sv2v_reg,
  mem_2465_sv2v_reg,mem_2464_sv2v_reg,mem_2463_sv2v_reg,mem_2462_sv2v_reg,
  mem_2461_sv2v_reg,mem_2460_sv2v_reg,mem_2459_sv2v_reg,mem_2458_sv2v_reg,mem_2457_sv2v_reg,
  mem_2456_sv2v_reg,mem_2455_sv2v_reg,mem_2454_sv2v_reg,mem_2453_sv2v_reg,
  mem_2452_sv2v_reg,mem_2451_sv2v_reg,mem_2450_sv2v_reg,mem_2449_sv2v_reg,mem_2448_sv2v_reg,
  mem_2447_sv2v_reg,mem_2446_sv2v_reg,mem_2445_sv2v_reg,mem_2444_sv2v_reg,
  mem_2443_sv2v_reg,mem_2442_sv2v_reg,mem_2441_sv2v_reg,mem_2440_sv2v_reg,
  mem_2439_sv2v_reg,mem_2438_sv2v_reg,mem_2437_sv2v_reg,mem_2436_sv2v_reg,mem_2435_sv2v_reg,
  mem_2434_sv2v_reg,mem_2433_sv2v_reg,mem_2432_sv2v_reg,mem_2431_sv2v_reg,
  mem_2430_sv2v_reg,mem_2429_sv2v_reg,mem_2428_sv2v_reg,mem_2427_sv2v_reg,mem_2426_sv2v_reg,
  mem_2425_sv2v_reg,mem_2424_sv2v_reg,mem_2423_sv2v_reg,mem_2422_sv2v_reg,
  mem_2421_sv2v_reg,mem_2420_sv2v_reg,mem_2419_sv2v_reg,mem_2418_sv2v_reg,mem_2417_sv2v_reg,
  mem_2416_sv2v_reg,mem_2415_sv2v_reg,mem_2414_sv2v_reg,mem_2413_sv2v_reg,
  mem_2412_sv2v_reg,mem_2411_sv2v_reg,mem_2410_sv2v_reg,mem_2409_sv2v_reg,mem_2408_sv2v_reg,
  mem_2407_sv2v_reg,mem_2406_sv2v_reg,mem_2405_sv2v_reg,mem_2404_sv2v_reg,
  mem_2403_sv2v_reg,mem_2402_sv2v_reg,mem_2401_sv2v_reg,mem_2400_sv2v_reg,
  mem_2399_sv2v_reg,mem_2398_sv2v_reg,mem_2397_sv2v_reg,mem_2396_sv2v_reg,mem_2395_sv2v_reg,
  mem_2394_sv2v_reg,mem_2393_sv2v_reg,mem_2392_sv2v_reg,mem_2391_sv2v_reg,
  mem_2390_sv2v_reg,mem_2389_sv2v_reg,mem_2388_sv2v_reg,mem_2387_sv2v_reg,mem_2386_sv2v_reg,
  mem_2385_sv2v_reg,mem_2384_sv2v_reg,mem_2383_sv2v_reg,mem_2382_sv2v_reg,
  mem_2381_sv2v_reg,mem_2380_sv2v_reg,mem_2379_sv2v_reg,mem_2378_sv2v_reg,mem_2377_sv2v_reg,
  mem_2376_sv2v_reg,mem_2375_sv2v_reg,mem_2374_sv2v_reg,mem_2373_sv2v_reg,
  mem_2372_sv2v_reg,mem_2371_sv2v_reg,mem_2370_sv2v_reg,mem_2369_sv2v_reg,mem_2368_sv2v_reg,
  mem_2367_sv2v_reg,mem_2366_sv2v_reg,mem_2365_sv2v_reg,mem_2364_sv2v_reg,
  mem_2363_sv2v_reg,mem_2362_sv2v_reg,mem_2361_sv2v_reg,mem_2360_sv2v_reg,
  mem_2359_sv2v_reg,mem_2358_sv2v_reg,mem_2357_sv2v_reg,mem_2356_sv2v_reg,mem_2355_sv2v_reg,
  mem_2354_sv2v_reg,mem_2353_sv2v_reg,mem_2352_sv2v_reg,mem_2351_sv2v_reg,
  mem_2350_sv2v_reg,mem_2349_sv2v_reg,mem_2348_sv2v_reg,mem_2347_sv2v_reg,mem_2346_sv2v_reg,
  mem_2345_sv2v_reg,mem_2344_sv2v_reg,mem_2343_sv2v_reg,mem_2342_sv2v_reg,
  mem_2341_sv2v_reg,mem_2340_sv2v_reg,mem_2339_sv2v_reg,mem_2338_sv2v_reg,mem_2337_sv2v_reg,
  mem_2336_sv2v_reg,mem_2335_sv2v_reg,mem_2334_sv2v_reg,mem_2333_sv2v_reg,
  mem_2332_sv2v_reg,mem_2331_sv2v_reg,mem_2330_sv2v_reg,mem_2329_sv2v_reg,mem_2328_sv2v_reg,
  mem_2327_sv2v_reg,mem_2326_sv2v_reg,mem_2325_sv2v_reg,mem_2324_sv2v_reg,
  mem_2323_sv2v_reg,mem_2322_sv2v_reg,mem_2321_sv2v_reg,mem_2320_sv2v_reg,
  mem_2319_sv2v_reg,mem_2318_sv2v_reg,mem_2317_sv2v_reg,mem_2316_sv2v_reg,mem_2315_sv2v_reg,
  mem_2314_sv2v_reg,mem_2313_sv2v_reg,mem_2312_sv2v_reg,mem_2311_sv2v_reg,
  mem_2310_sv2v_reg,mem_2309_sv2v_reg,mem_2308_sv2v_reg,mem_2307_sv2v_reg,mem_2306_sv2v_reg,
  mem_2305_sv2v_reg,mem_2304_sv2v_reg,mem_2303_sv2v_reg,mem_2302_sv2v_reg,
  mem_2301_sv2v_reg,mem_2300_sv2v_reg,mem_2299_sv2v_reg,mem_2298_sv2v_reg,mem_2297_sv2v_reg,
  mem_2296_sv2v_reg,mem_2295_sv2v_reg,mem_2294_sv2v_reg,mem_2293_sv2v_reg,
  mem_2292_sv2v_reg,mem_2291_sv2v_reg,mem_2290_sv2v_reg,mem_2289_sv2v_reg,mem_2288_sv2v_reg,
  mem_2287_sv2v_reg,mem_2286_sv2v_reg,mem_2285_sv2v_reg,mem_2284_sv2v_reg,
  mem_2283_sv2v_reg,mem_2282_sv2v_reg,mem_2281_sv2v_reg,mem_2280_sv2v_reg,
  mem_2279_sv2v_reg,mem_2278_sv2v_reg,mem_2277_sv2v_reg,mem_2276_sv2v_reg,mem_2275_sv2v_reg,
  mem_2274_sv2v_reg,mem_2273_sv2v_reg,mem_2272_sv2v_reg,mem_2271_sv2v_reg,
  mem_2270_sv2v_reg,mem_2269_sv2v_reg,mem_2268_sv2v_reg,mem_2267_sv2v_reg,mem_2266_sv2v_reg,
  mem_2265_sv2v_reg,mem_2264_sv2v_reg,mem_2263_sv2v_reg,mem_2262_sv2v_reg,
  mem_2261_sv2v_reg,mem_2260_sv2v_reg,mem_2259_sv2v_reg,mem_2258_sv2v_reg,mem_2257_sv2v_reg,
  mem_2256_sv2v_reg,mem_2255_sv2v_reg,mem_2254_sv2v_reg,mem_2253_sv2v_reg,
  mem_2252_sv2v_reg,mem_2251_sv2v_reg,mem_2250_sv2v_reg,mem_2249_sv2v_reg,mem_2248_sv2v_reg,
  mem_2247_sv2v_reg,mem_2246_sv2v_reg,mem_2245_sv2v_reg,mem_2244_sv2v_reg,
  mem_2243_sv2v_reg,mem_2242_sv2v_reg,mem_2241_sv2v_reg,mem_2240_sv2v_reg,
  mem_2239_sv2v_reg,mem_2238_sv2v_reg,mem_2237_sv2v_reg,mem_2236_sv2v_reg,mem_2235_sv2v_reg,
  mem_2234_sv2v_reg,mem_2233_sv2v_reg,mem_2232_sv2v_reg,mem_2231_sv2v_reg,
  mem_2230_sv2v_reg,mem_2229_sv2v_reg,mem_2228_sv2v_reg,mem_2227_sv2v_reg,mem_2226_sv2v_reg,
  mem_2225_sv2v_reg,mem_2224_sv2v_reg,mem_2223_sv2v_reg,mem_2222_sv2v_reg,
  mem_2221_sv2v_reg,mem_2220_sv2v_reg,mem_2219_sv2v_reg,mem_2218_sv2v_reg,mem_2217_sv2v_reg,
  mem_2216_sv2v_reg,mem_2215_sv2v_reg,mem_2214_sv2v_reg,mem_2213_sv2v_reg,
  mem_2212_sv2v_reg,mem_2211_sv2v_reg,mem_2210_sv2v_reg,mem_2209_sv2v_reg,mem_2208_sv2v_reg,
  mem_2207_sv2v_reg,mem_2206_sv2v_reg,mem_2205_sv2v_reg,mem_2204_sv2v_reg,
  mem_2203_sv2v_reg,mem_2202_sv2v_reg,mem_2201_sv2v_reg,mem_2200_sv2v_reg,
  mem_2199_sv2v_reg,mem_2198_sv2v_reg,mem_2197_sv2v_reg,mem_2196_sv2v_reg,mem_2195_sv2v_reg,
  mem_2194_sv2v_reg,mem_2193_sv2v_reg,mem_2192_sv2v_reg,mem_2191_sv2v_reg,
  mem_2190_sv2v_reg,mem_2189_sv2v_reg,mem_2188_sv2v_reg,mem_2187_sv2v_reg,mem_2186_sv2v_reg,
  mem_2185_sv2v_reg,mem_2184_sv2v_reg,mem_2183_sv2v_reg,mem_2182_sv2v_reg,
  mem_2181_sv2v_reg,mem_2180_sv2v_reg,mem_2179_sv2v_reg,mem_2178_sv2v_reg,mem_2177_sv2v_reg,
  mem_2176_sv2v_reg,mem_2175_sv2v_reg,mem_2174_sv2v_reg,mem_2173_sv2v_reg,
  mem_2172_sv2v_reg,mem_2171_sv2v_reg,mem_2170_sv2v_reg,mem_2169_sv2v_reg,mem_2168_sv2v_reg,
  mem_2167_sv2v_reg,mem_2166_sv2v_reg,mem_2165_sv2v_reg,mem_2164_sv2v_reg,
  mem_2163_sv2v_reg,mem_2162_sv2v_reg,mem_2161_sv2v_reg,mem_2160_sv2v_reg,
  mem_2159_sv2v_reg,mem_2158_sv2v_reg,mem_2157_sv2v_reg,mem_2156_sv2v_reg,mem_2155_sv2v_reg,
  mem_2154_sv2v_reg,mem_2153_sv2v_reg,mem_2152_sv2v_reg,mem_2151_sv2v_reg,
  mem_2150_sv2v_reg,mem_2149_sv2v_reg,mem_2148_sv2v_reg,mem_2147_sv2v_reg,mem_2146_sv2v_reg,
  mem_2145_sv2v_reg,mem_2144_sv2v_reg,mem_2143_sv2v_reg,mem_2142_sv2v_reg,
  mem_2141_sv2v_reg,mem_2140_sv2v_reg,mem_2139_sv2v_reg,mem_2138_sv2v_reg,mem_2137_sv2v_reg,
  mem_2136_sv2v_reg,mem_2135_sv2v_reg,mem_2134_sv2v_reg,mem_2133_sv2v_reg,
  mem_2132_sv2v_reg,mem_2131_sv2v_reg,mem_2130_sv2v_reg,mem_2129_sv2v_reg,mem_2128_sv2v_reg,
  mem_2127_sv2v_reg,mem_2126_sv2v_reg,mem_2125_sv2v_reg,mem_2124_sv2v_reg,
  mem_2123_sv2v_reg,mem_2122_sv2v_reg,mem_2121_sv2v_reg,mem_2120_sv2v_reg,
  mem_2119_sv2v_reg,mem_2118_sv2v_reg,mem_2117_sv2v_reg,mem_2116_sv2v_reg,mem_2115_sv2v_reg,
  mem_2114_sv2v_reg,mem_2113_sv2v_reg,mem_2112_sv2v_reg,mem_2111_sv2v_reg,
  mem_2110_sv2v_reg,mem_2109_sv2v_reg,mem_2108_sv2v_reg,mem_2107_sv2v_reg,mem_2106_sv2v_reg,
  mem_2105_sv2v_reg,mem_2104_sv2v_reg,mem_2103_sv2v_reg,mem_2102_sv2v_reg,
  mem_2101_sv2v_reg,mem_2100_sv2v_reg,mem_2099_sv2v_reg,mem_2098_sv2v_reg,mem_2097_sv2v_reg,
  mem_2096_sv2v_reg,mem_2095_sv2v_reg,mem_2094_sv2v_reg,mem_2093_sv2v_reg,
  mem_2092_sv2v_reg,mem_2091_sv2v_reg,mem_2090_sv2v_reg,mem_2089_sv2v_reg,mem_2088_sv2v_reg,
  mem_2087_sv2v_reg,mem_2086_sv2v_reg,mem_2085_sv2v_reg,mem_2084_sv2v_reg,
  mem_2083_sv2v_reg,mem_2082_sv2v_reg,mem_2081_sv2v_reg,mem_2080_sv2v_reg,
  mem_2079_sv2v_reg,mem_2078_sv2v_reg,mem_2077_sv2v_reg,mem_2076_sv2v_reg,mem_2075_sv2v_reg,
  mem_2074_sv2v_reg,mem_2073_sv2v_reg,mem_2072_sv2v_reg,mem_2071_sv2v_reg,
  mem_2070_sv2v_reg,mem_2069_sv2v_reg,mem_2068_sv2v_reg,mem_2067_sv2v_reg,mem_2066_sv2v_reg,
  mem_2065_sv2v_reg,mem_2064_sv2v_reg,mem_2063_sv2v_reg,mem_2062_sv2v_reg,
  mem_2061_sv2v_reg,mem_2060_sv2v_reg,mem_2059_sv2v_reg,mem_2058_sv2v_reg,mem_2057_sv2v_reg,
  mem_2056_sv2v_reg,mem_2055_sv2v_reg,mem_2054_sv2v_reg,mem_2053_sv2v_reg,
  mem_2052_sv2v_reg,mem_2051_sv2v_reg,mem_2050_sv2v_reg,mem_2049_sv2v_reg,mem_2048_sv2v_reg,
  mem_2047_sv2v_reg,mem_2046_sv2v_reg,mem_2045_sv2v_reg,mem_2044_sv2v_reg,
  mem_2043_sv2v_reg,mem_2042_sv2v_reg,mem_2041_sv2v_reg,mem_2040_sv2v_reg,
  mem_2039_sv2v_reg,mem_2038_sv2v_reg,mem_2037_sv2v_reg,mem_2036_sv2v_reg,mem_2035_sv2v_reg,
  mem_2034_sv2v_reg,mem_2033_sv2v_reg,mem_2032_sv2v_reg,mem_2031_sv2v_reg,
  mem_2030_sv2v_reg,mem_2029_sv2v_reg,mem_2028_sv2v_reg,mem_2027_sv2v_reg,mem_2026_sv2v_reg,
  mem_2025_sv2v_reg,mem_2024_sv2v_reg,mem_2023_sv2v_reg,mem_2022_sv2v_reg,
  mem_2021_sv2v_reg,mem_2020_sv2v_reg,mem_2019_sv2v_reg,mem_2018_sv2v_reg,mem_2017_sv2v_reg,
  mem_2016_sv2v_reg,mem_2015_sv2v_reg,mem_2014_sv2v_reg,mem_2013_sv2v_reg,
  mem_2012_sv2v_reg,mem_2011_sv2v_reg,mem_2010_sv2v_reg,mem_2009_sv2v_reg,mem_2008_sv2v_reg,
  mem_2007_sv2v_reg,mem_2006_sv2v_reg,mem_2005_sv2v_reg,mem_2004_sv2v_reg,
  mem_2003_sv2v_reg,mem_2002_sv2v_reg,mem_2001_sv2v_reg,mem_2000_sv2v_reg,
  mem_1999_sv2v_reg,mem_1998_sv2v_reg,mem_1997_sv2v_reg,mem_1996_sv2v_reg,mem_1995_sv2v_reg,
  mem_1994_sv2v_reg,mem_1993_sv2v_reg,mem_1992_sv2v_reg,mem_1991_sv2v_reg,
  mem_1990_sv2v_reg,mem_1989_sv2v_reg,mem_1988_sv2v_reg,mem_1987_sv2v_reg,mem_1986_sv2v_reg,
  mem_1985_sv2v_reg,mem_1984_sv2v_reg,mem_1983_sv2v_reg,mem_1982_sv2v_reg,
  mem_1981_sv2v_reg,mem_1980_sv2v_reg,mem_1979_sv2v_reg,mem_1978_sv2v_reg,mem_1977_sv2v_reg,
  mem_1976_sv2v_reg,mem_1975_sv2v_reg,mem_1974_sv2v_reg,mem_1973_sv2v_reg,
  mem_1972_sv2v_reg,mem_1971_sv2v_reg,mem_1970_sv2v_reg,mem_1969_sv2v_reg,mem_1968_sv2v_reg,
  mem_1967_sv2v_reg,mem_1966_sv2v_reg,mem_1965_sv2v_reg,mem_1964_sv2v_reg,
  mem_1963_sv2v_reg,mem_1962_sv2v_reg,mem_1961_sv2v_reg,mem_1960_sv2v_reg,
  mem_1959_sv2v_reg,mem_1958_sv2v_reg,mem_1957_sv2v_reg,mem_1956_sv2v_reg,mem_1955_sv2v_reg,
  mem_1954_sv2v_reg,mem_1953_sv2v_reg,mem_1952_sv2v_reg,mem_1951_sv2v_reg,
  mem_1950_sv2v_reg,mem_1949_sv2v_reg,mem_1948_sv2v_reg,mem_1947_sv2v_reg,mem_1946_sv2v_reg,
  mem_1945_sv2v_reg,mem_1944_sv2v_reg,mem_1943_sv2v_reg,mem_1942_sv2v_reg,
  mem_1941_sv2v_reg,mem_1940_sv2v_reg,mem_1939_sv2v_reg,mem_1938_sv2v_reg,mem_1937_sv2v_reg,
  mem_1936_sv2v_reg,mem_1935_sv2v_reg,mem_1934_sv2v_reg,mem_1933_sv2v_reg,
  mem_1932_sv2v_reg,mem_1931_sv2v_reg,mem_1930_sv2v_reg,mem_1929_sv2v_reg,mem_1928_sv2v_reg,
  mem_1927_sv2v_reg,mem_1926_sv2v_reg,mem_1925_sv2v_reg,mem_1924_sv2v_reg,
  mem_1923_sv2v_reg,mem_1922_sv2v_reg,mem_1921_sv2v_reg,mem_1920_sv2v_reg,
  mem_1919_sv2v_reg,mem_1918_sv2v_reg,mem_1917_sv2v_reg,mem_1916_sv2v_reg,mem_1915_sv2v_reg,
  mem_1914_sv2v_reg,mem_1913_sv2v_reg,mem_1912_sv2v_reg,mem_1911_sv2v_reg,
  mem_1910_sv2v_reg,mem_1909_sv2v_reg,mem_1908_sv2v_reg,mem_1907_sv2v_reg,mem_1906_sv2v_reg,
  mem_1905_sv2v_reg,mem_1904_sv2v_reg,mem_1903_sv2v_reg,mem_1902_sv2v_reg,
  mem_1901_sv2v_reg,mem_1900_sv2v_reg,mem_1899_sv2v_reg,mem_1898_sv2v_reg,mem_1897_sv2v_reg,
  mem_1896_sv2v_reg,mem_1895_sv2v_reg,mem_1894_sv2v_reg,mem_1893_sv2v_reg,
  mem_1892_sv2v_reg,mem_1891_sv2v_reg,mem_1890_sv2v_reg,mem_1889_sv2v_reg,mem_1888_sv2v_reg,
  mem_1887_sv2v_reg,mem_1886_sv2v_reg,mem_1885_sv2v_reg,mem_1884_sv2v_reg,
  mem_1883_sv2v_reg,mem_1882_sv2v_reg,mem_1881_sv2v_reg,mem_1880_sv2v_reg,
  mem_1879_sv2v_reg,mem_1878_sv2v_reg,mem_1877_sv2v_reg,mem_1876_sv2v_reg,mem_1875_sv2v_reg,
  mem_1874_sv2v_reg,mem_1873_sv2v_reg,mem_1872_sv2v_reg,mem_1871_sv2v_reg,
  mem_1870_sv2v_reg,mem_1869_sv2v_reg,mem_1868_sv2v_reg,mem_1867_sv2v_reg,mem_1866_sv2v_reg,
  mem_1865_sv2v_reg,mem_1864_sv2v_reg,mem_1863_sv2v_reg,mem_1862_sv2v_reg,
  mem_1861_sv2v_reg,mem_1860_sv2v_reg,mem_1859_sv2v_reg,mem_1858_sv2v_reg,mem_1857_sv2v_reg,
  mem_1856_sv2v_reg,mem_1855_sv2v_reg,mem_1854_sv2v_reg,mem_1853_sv2v_reg,
  mem_1852_sv2v_reg,mem_1851_sv2v_reg,mem_1850_sv2v_reg,mem_1849_sv2v_reg,mem_1848_sv2v_reg,
  mem_1847_sv2v_reg,mem_1846_sv2v_reg,mem_1845_sv2v_reg,mem_1844_sv2v_reg,
  mem_1843_sv2v_reg,mem_1842_sv2v_reg,mem_1841_sv2v_reg,mem_1840_sv2v_reg,
  mem_1839_sv2v_reg,mem_1838_sv2v_reg,mem_1837_sv2v_reg,mem_1836_sv2v_reg,mem_1835_sv2v_reg,
  mem_1834_sv2v_reg,mem_1833_sv2v_reg,mem_1832_sv2v_reg,mem_1831_sv2v_reg,
  mem_1830_sv2v_reg,mem_1829_sv2v_reg,mem_1828_sv2v_reg,mem_1827_sv2v_reg,mem_1826_sv2v_reg,
  mem_1825_sv2v_reg,mem_1824_sv2v_reg,mem_1823_sv2v_reg,mem_1822_sv2v_reg,
  mem_1821_sv2v_reg,mem_1820_sv2v_reg,mem_1819_sv2v_reg,mem_1818_sv2v_reg,mem_1817_sv2v_reg,
  mem_1816_sv2v_reg,mem_1815_sv2v_reg,mem_1814_sv2v_reg,mem_1813_sv2v_reg,
  mem_1812_sv2v_reg,mem_1811_sv2v_reg,mem_1810_sv2v_reg,mem_1809_sv2v_reg,mem_1808_sv2v_reg,
  mem_1807_sv2v_reg,mem_1806_sv2v_reg,mem_1805_sv2v_reg,mem_1804_sv2v_reg,
  mem_1803_sv2v_reg,mem_1802_sv2v_reg,mem_1801_sv2v_reg,mem_1800_sv2v_reg,
  mem_1799_sv2v_reg,mem_1798_sv2v_reg,mem_1797_sv2v_reg,mem_1796_sv2v_reg,mem_1795_sv2v_reg,
  mem_1794_sv2v_reg,mem_1793_sv2v_reg,mem_1792_sv2v_reg,mem_1791_sv2v_reg,
  mem_1790_sv2v_reg,mem_1789_sv2v_reg,mem_1788_sv2v_reg,mem_1787_sv2v_reg,mem_1786_sv2v_reg,
  mem_1785_sv2v_reg,mem_1784_sv2v_reg,mem_1783_sv2v_reg,mem_1782_sv2v_reg,
  mem_1781_sv2v_reg,mem_1780_sv2v_reg,mem_1779_sv2v_reg,mem_1778_sv2v_reg,mem_1777_sv2v_reg,
  mem_1776_sv2v_reg,mem_1775_sv2v_reg,mem_1774_sv2v_reg,mem_1773_sv2v_reg,
  mem_1772_sv2v_reg,mem_1771_sv2v_reg,mem_1770_sv2v_reg,mem_1769_sv2v_reg,mem_1768_sv2v_reg,
  mem_1767_sv2v_reg,mem_1766_sv2v_reg,mem_1765_sv2v_reg,mem_1764_sv2v_reg,
  mem_1763_sv2v_reg,mem_1762_sv2v_reg,mem_1761_sv2v_reg,mem_1760_sv2v_reg,
  mem_1759_sv2v_reg,mem_1758_sv2v_reg,mem_1757_sv2v_reg,mem_1756_sv2v_reg,mem_1755_sv2v_reg,
  mem_1754_sv2v_reg,mem_1753_sv2v_reg,mem_1752_sv2v_reg,mem_1751_sv2v_reg,
  mem_1750_sv2v_reg,mem_1749_sv2v_reg,mem_1748_sv2v_reg,mem_1747_sv2v_reg,mem_1746_sv2v_reg,
  mem_1745_sv2v_reg,mem_1744_sv2v_reg,mem_1743_sv2v_reg,mem_1742_sv2v_reg,
  mem_1741_sv2v_reg,mem_1740_sv2v_reg,mem_1739_sv2v_reg,mem_1738_sv2v_reg,mem_1737_sv2v_reg,
  mem_1736_sv2v_reg,mem_1735_sv2v_reg,mem_1734_sv2v_reg,mem_1733_sv2v_reg,
  mem_1732_sv2v_reg,mem_1731_sv2v_reg,mem_1730_sv2v_reg,mem_1729_sv2v_reg,mem_1728_sv2v_reg,
  mem_1727_sv2v_reg,mem_1726_sv2v_reg,mem_1725_sv2v_reg,mem_1724_sv2v_reg,
  mem_1723_sv2v_reg,mem_1722_sv2v_reg,mem_1721_sv2v_reg,mem_1720_sv2v_reg,
  mem_1719_sv2v_reg,mem_1718_sv2v_reg,mem_1717_sv2v_reg,mem_1716_sv2v_reg,mem_1715_sv2v_reg,
  mem_1714_sv2v_reg,mem_1713_sv2v_reg,mem_1712_sv2v_reg,mem_1711_sv2v_reg,
  mem_1710_sv2v_reg,mem_1709_sv2v_reg,mem_1708_sv2v_reg,mem_1707_sv2v_reg,mem_1706_sv2v_reg,
  mem_1705_sv2v_reg,mem_1704_sv2v_reg,mem_1703_sv2v_reg,mem_1702_sv2v_reg,
  mem_1701_sv2v_reg,mem_1700_sv2v_reg,mem_1699_sv2v_reg,mem_1698_sv2v_reg,mem_1697_sv2v_reg,
  mem_1696_sv2v_reg,mem_1695_sv2v_reg,mem_1694_sv2v_reg,mem_1693_sv2v_reg,
  mem_1692_sv2v_reg,mem_1691_sv2v_reg,mem_1690_sv2v_reg,mem_1689_sv2v_reg,mem_1688_sv2v_reg,
  mem_1687_sv2v_reg,mem_1686_sv2v_reg,mem_1685_sv2v_reg,mem_1684_sv2v_reg,
  mem_1683_sv2v_reg,mem_1682_sv2v_reg,mem_1681_sv2v_reg,mem_1680_sv2v_reg,
  mem_1679_sv2v_reg,mem_1678_sv2v_reg,mem_1677_sv2v_reg,mem_1676_sv2v_reg,mem_1675_sv2v_reg,
  mem_1674_sv2v_reg,mem_1673_sv2v_reg,mem_1672_sv2v_reg,mem_1671_sv2v_reg,
  mem_1670_sv2v_reg,mem_1669_sv2v_reg,mem_1668_sv2v_reg,mem_1667_sv2v_reg,mem_1666_sv2v_reg,
  mem_1665_sv2v_reg,mem_1664_sv2v_reg,mem_1663_sv2v_reg,mem_1662_sv2v_reg,
  mem_1661_sv2v_reg,mem_1660_sv2v_reg,mem_1659_sv2v_reg,mem_1658_sv2v_reg,mem_1657_sv2v_reg,
  mem_1656_sv2v_reg,mem_1655_sv2v_reg,mem_1654_sv2v_reg,mem_1653_sv2v_reg,
  mem_1652_sv2v_reg,mem_1651_sv2v_reg,mem_1650_sv2v_reg,mem_1649_sv2v_reg,mem_1648_sv2v_reg,
  mem_1647_sv2v_reg,mem_1646_sv2v_reg,mem_1645_sv2v_reg,mem_1644_sv2v_reg,
  mem_1643_sv2v_reg,mem_1642_sv2v_reg,mem_1641_sv2v_reg,mem_1640_sv2v_reg,
  mem_1639_sv2v_reg,mem_1638_sv2v_reg,mem_1637_sv2v_reg,mem_1636_sv2v_reg,mem_1635_sv2v_reg,
  mem_1634_sv2v_reg,mem_1633_sv2v_reg,mem_1632_sv2v_reg,mem_1631_sv2v_reg,
  mem_1630_sv2v_reg,mem_1629_sv2v_reg,mem_1628_sv2v_reg,mem_1627_sv2v_reg,mem_1626_sv2v_reg,
  mem_1625_sv2v_reg,mem_1624_sv2v_reg,mem_1623_sv2v_reg,mem_1622_sv2v_reg,
  mem_1621_sv2v_reg,mem_1620_sv2v_reg,mem_1619_sv2v_reg,mem_1618_sv2v_reg,mem_1617_sv2v_reg,
  mem_1616_sv2v_reg,mem_1615_sv2v_reg,mem_1614_sv2v_reg,mem_1613_sv2v_reg,
  mem_1612_sv2v_reg,mem_1611_sv2v_reg,mem_1610_sv2v_reg,mem_1609_sv2v_reg,mem_1608_sv2v_reg,
  mem_1607_sv2v_reg,mem_1606_sv2v_reg,mem_1605_sv2v_reg,mem_1604_sv2v_reg,
  mem_1603_sv2v_reg,mem_1602_sv2v_reg,mem_1601_sv2v_reg,mem_1600_sv2v_reg,
  mem_1599_sv2v_reg,mem_1598_sv2v_reg,mem_1597_sv2v_reg,mem_1596_sv2v_reg,mem_1595_sv2v_reg,
  mem_1594_sv2v_reg,mem_1593_sv2v_reg,mem_1592_sv2v_reg,mem_1591_sv2v_reg,
  mem_1590_sv2v_reg,mem_1589_sv2v_reg,mem_1588_sv2v_reg,mem_1587_sv2v_reg,mem_1586_sv2v_reg,
  mem_1585_sv2v_reg,mem_1584_sv2v_reg,mem_1583_sv2v_reg,mem_1582_sv2v_reg,
  mem_1581_sv2v_reg,mem_1580_sv2v_reg,mem_1579_sv2v_reg,mem_1578_sv2v_reg,mem_1577_sv2v_reg,
  mem_1576_sv2v_reg,mem_1575_sv2v_reg,mem_1574_sv2v_reg,mem_1573_sv2v_reg,
  mem_1572_sv2v_reg,mem_1571_sv2v_reg,mem_1570_sv2v_reg,mem_1569_sv2v_reg,mem_1568_sv2v_reg,
  mem_1567_sv2v_reg,mem_1566_sv2v_reg,mem_1565_sv2v_reg,mem_1564_sv2v_reg,
  mem_1563_sv2v_reg,mem_1562_sv2v_reg,mem_1561_sv2v_reg,mem_1560_sv2v_reg,
  mem_1559_sv2v_reg,mem_1558_sv2v_reg,mem_1557_sv2v_reg,mem_1556_sv2v_reg,mem_1555_sv2v_reg,
  mem_1554_sv2v_reg,mem_1553_sv2v_reg,mem_1552_sv2v_reg,mem_1551_sv2v_reg,
  mem_1550_sv2v_reg,mem_1549_sv2v_reg,mem_1548_sv2v_reg,mem_1547_sv2v_reg,mem_1546_sv2v_reg,
  mem_1545_sv2v_reg,mem_1544_sv2v_reg,mem_1543_sv2v_reg,mem_1542_sv2v_reg,
  mem_1541_sv2v_reg,mem_1540_sv2v_reg,mem_1539_sv2v_reg,mem_1538_sv2v_reg,mem_1537_sv2v_reg,
  mem_1536_sv2v_reg,mem_1535_sv2v_reg,mem_1534_sv2v_reg,mem_1533_sv2v_reg,
  mem_1532_sv2v_reg,mem_1531_sv2v_reg,mem_1530_sv2v_reg,mem_1529_sv2v_reg,mem_1528_sv2v_reg,
  mem_1527_sv2v_reg,mem_1526_sv2v_reg,mem_1525_sv2v_reg,mem_1524_sv2v_reg,
  mem_1523_sv2v_reg,mem_1522_sv2v_reg,mem_1521_sv2v_reg,mem_1520_sv2v_reg,
  mem_1519_sv2v_reg,mem_1518_sv2v_reg,mem_1517_sv2v_reg,mem_1516_sv2v_reg,mem_1515_sv2v_reg,
  mem_1514_sv2v_reg,mem_1513_sv2v_reg,mem_1512_sv2v_reg,mem_1511_sv2v_reg,
  mem_1510_sv2v_reg,mem_1509_sv2v_reg,mem_1508_sv2v_reg,mem_1507_sv2v_reg,mem_1506_sv2v_reg,
  mem_1505_sv2v_reg,mem_1504_sv2v_reg,mem_1503_sv2v_reg,mem_1502_sv2v_reg,
  mem_1501_sv2v_reg,mem_1500_sv2v_reg,mem_1499_sv2v_reg,mem_1498_sv2v_reg,mem_1497_sv2v_reg,
  mem_1496_sv2v_reg,mem_1495_sv2v_reg,mem_1494_sv2v_reg,mem_1493_sv2v_reg,
  mem_1492_sv2v_reg,mem_1491_sv2v_reg,mem_1490_sv2v_reg,mem_1489_sv2v_reg,mem_1488_sv2v_reg,
  mem_1487_sv2v_reg,mem_1486_sv2v_reg,mem_1485_sv2v_reg,mem_1484_sv2v_reg,
  mem_1483_sv2v_reg,mem_1482_sv2v_reg,mem_1481_sv2v_reg,mem_1480_sv2v_reg,
  mem_1479_sv2v_reg,mem_1478_sv2v_reg,mem_1477_sv2v_reg,mem_1476_sv2v_reg,mem_1475_sv2v_reg,
  mem_1474_sv2v_reg,mem_1473_sv2v_reg,mem_1472_sv2v_reg,mem_1471_sv2v_reg,
  mem_1470_sv2v_reg,mem_1469_sv2v_reg,mem_1468_sv2v_reg,mem_1467_sv2v_reg,mem_1466_sv2v_reg,
  mem_1465_sv2v_reg,mem_1464_sv2v_reg,mem_1463_sv2v_reg,mem_1462_sv2v_reg,
  mem_1461_sv2v_reg,mem_1460_sv2v_reg,mem_1459_sv2v_reg,mem_1458_sv2v_reg,mem_1457_sv2v_reg,
  mem_1456_sv2v_reg,mem_1455_sv2v_reg,mem_1454_sv2v_reg,mem_1453_sv2v_reg,
  mem_1452_sv2v_reg,mem_1451_sv2v_reg,mem_1450_sv2v_reg,mem_1449_sv2v_reg,mem_1448_sv2v_reg,
  mem_1447_sv2v_reg,mem_1446_sv2v_reg,mem_1445_sv2v_reg,mem_1444_sv2v_reg,
  mem_1443_sv2v_reg,mem_1442_sv2v_reg,mem_1441_sv2v_reg,mem_1440_sv2v_reg,
  mem_1439_sv2v_reg,mem_1438_sv2v_reg,mem_1437_sv2v_reg,mem_1436_sv2v_reg,mem_1435_sv2v_reg,
  mem_1434_sv2v_reg,mem_1433_sv2v_reg,mem_1432_sv2v_reg,mem_1431_sv2v_reg,
  mem_1430_sv2v_reg,mem_1429_sv2v_reg,mem_1428_sv2v_reg,mem_1427_sv2v_reg,mem_1426_sv2v_reg,
  mem_1425_sv2v_reg,mem_1424_sv2v_reg,mem_1423_sv2v_reg,mem_1422_sv2v_reg,
  mem_1421_sv2v_reg,mem_1420_sv2v_reg,mem_1419_sv2v_reg,mem_1418_sv2v_reg,mem_1417_sv2v_reg,
  mem_1416_sv2v_reg,mem_1415_sv2v_reg,mem_1414_sv2v_reg,mem_1413_sv2v_reg,
  mem_1412_sv2v_reg,mem_1411_sv2v_reg,mem_1410_sv2v_reg,mem_1409_sv2v_reg,mem_1408_sv2v_reg,
  mem_1407_sv2v_reg,mem_1406_sv2v_reg,mem_1405_sv2v_reg,mem_1404_sv2v_reg,
  mem_1403_sv2v_reg,mem_1402_sv2v_reg,mem_1401_sv2v_reg,mem_1400_sv2v_reg,
  mem_1399_sv2v_reg,mem_1398_sv2v_reg,mem_1397_sv2v_reg,mem_1396_sv2v_reg,mem_1395_sv2v_reg,
  mem_1394_sv2v_reg,mem_1393_sv2v_reg,mem_1392_sv2v_reg,mem_1391_sv2v_reg,
  mem_1390_sv2v_reg,mem_1389_sv2v_reg,mem_1388_sv2v_reg,mem_1387_sv2v_reg,mem_1386_sv2v_reg,
  mem_1385_sv2v_reg,mem_1384_sv2v_reg,mem_1383_sv2v_reg,mem_1382_sv2v_reg,
  mem_1381_sv2v_reg,mem_1380_sv2v_reg,mem_1379_sv2v_reg,mem_1378_sv2v_reg,mem_1377_sv2v_reg,
  mem_1376_sv2v_reg,mem_1375_sv2v_reg,mem_1374_sv2v_reg,mem_1373_sv2v_reg,
  mem_1372_sv2v_reg,mem_1371_sv2v_reg,mem_1370_sv2v_reg,mem_1369_sv2v_reg,mem_1368_sv2v_reg,
  mem_1367_sv2v_reg,mem_1366_sv2v_reg,mem_1365_sv2v_reg,mem_1364_sv2v_reg,
  mem_1363_sv2v_reg,mem_1362_sv2v_reg,mem_1361_sv2v_reg,mem_1360_sv2v_reg,
  mem_1359_sv2v_reg,mem_1358_sv2v_reg,mem_1357_sv2v_reg,mem_1356_sv2v_reg,mem_1355_sv2v_reg,
  mem_1354_sv2v_reg,mem_1353_sv2v_reg,mem_1352_sv2v_reg,mem_1351_sv2v_reg,
  mem_1350_sv2v_reg,mem_1349_sv2v_reg,mem_1348_sv2v_reg,mem_1347_sv2v_reg,mem_1346_sv2v_reg,
  mem_1345_sv2v_reg,mem_1344_sv2v_reg,mem_1343_sv2v_reg,mem_1342_sv2v_reg,
  mem_1341_sv2v_reg,mem_1340_sv2v_reg,mem_1339_sv2v_reg,mem_1338_sv2v_reg,mem_1337_sv2v_reg,
  mem_1336_sv2v_reg,mem_1335_sv2v_reg,mem_1334_sv2v_reg,mem_1333_sv2v_reg,
  mem_1332_sv2v_reg,mem_1331_sv2v_reg,mem_1330_sv2v_reg,mem_1329_sv2v_reg,mem_1328_sv2v_reg,
  mem_1327_sv2v_reg,mem_1326_sv2v_reg,mem_1325_sv2v_reg,mem_1324_sv2v_reg,
  mem_1323_sv2v_reg,mem_1322_sv2v_reg,mem_1321_sv2v_reg,mem_1320_sv2v_reg,
  mem_1319_sv2v_reg,mem_1318_sv2v_reg,mem_1317_sv2v_reg,mem_1316_sv2v_reg,mem_1315_sv2v_reg,
  mem_1314_sv2v_reg,mem_1313_sv2v_reg,mem_1312_sv2v_reg,mem_1311_sv2v_reg,
  mem_1310_sv2v_reg,mem_1309_sv2v_reg,mem_1308_sv2v_reg,mem_1307_sv2v_reg,mem_1306_sv2v_reg,
  mem_1305_sv2v_reg,mem_1304_sv2v_reg,mem_1303_sv2v_reg,mem_1302_sv2v_reg,
  mem_1301_sv2v_reg,mem_1300_sv2v_reg,mem_1299_sv2v_reg,mem_1298_sv2v_reg,mem_1297_sv2v_reg,
  mem_1296_sv2v_reg,mem_1295_sv2v_reg,mem_1294_sv2v_reg,mem_1293_sv2v_reg,
  mem_1292_sv2v_reg,mem_1291_sv2v_reg,mem_1290_sv2v_reg,mem_1289_sv2v_reg,mem_1288_sv2v_reg,
  mem_1287_sv2v_reg,mem_1286_sv2v_reg,mem_1285_sv2v_reg,mem_1284_sv2v_reg,
  mem_1283_sv2v_reg,mem_1282_sv2v_reg,mem_1281_sv2v_reg,mem_1280_sv2v_reg,
  mem_1279_sv2v_reg,mem_1278_sv2v_reg,mem_1277_sv2v_reg,mem_1276_sv2v_reg,mem_1275_sv2v_reg,
  mem_1274_sv2v_reg,mem_1273_sv2v_reg,mem_1272_sv2v_reg,mem_1271_sv2v_reg,
  mem_1270_sv2v_reg,mem_1269_sv2v_reg,mem_1268_sv2v_reg,mem_1267_sv2v_reg,mem_1266_sv2v_reg,
  mem_1265_sv2v_reg,mem_1264_sv2v_reg,mem_1263_sv2v_reg,mem_1262_sv2v_reg,
  mem_1261_sv2v_reg,mem_1260_sv2v_reg,mem_1259_sv2v_reg,mem_1258_sv2v_reg,mem_1257_sv2v_reg,
  mem_1256_sv2v_reg,mem_1255_sv2v_reg,mem_1254_sv2v_reg,mem_1253_sv2v_reg,
  mem_1252_sv2v_reg,mem_1251_sv2v_reg,mem_1250_sv2v_reg,mem_1249_sv2v_reg,mem_1248_sv2v_reg,
  mem_1247_sv2v_reg,mem_1246_sv2v_reg,mem_1245_sv2v_reg,mem_1244_sv2v_reg,
  mem_1243_sv2v_reg,mem_1242_sv2v_reg,mem_1241_sv2v_reg,mem_1240_sv2v_reg,
  mem_1239_sv2v_reg,mem_1238_sv2v_reg,mem_1237_sv2v_reg,mem_1236_sv2v_reg,mem_1235_sv2v_reg,
  mem_1234_sv2v_reg,mem_1233_sv2v_reg,mem_1232_sv2v_reg,mem_1231_sv2v_reg,
  mem_1230_sv2v_reg,mem_1229_sv2v_reg,mem_1228_sv2v_reg,mem_1227_sv2v_reg,mem_1226_sv2v_reg,
  mem_1225_sv2v_reg,mem_1224_sv2v_reg,mem_1223_sv2v_reg,mem_1222_sv2v_reg,
  mem_1221_sv2v_reg,mem_1220_sv2v_reg,mem_1219_sv2v_reg,mem_1218_sv2v_reg,mem_1217_sv2v_reg,
  mem_1216_sv2v_reg,mem_1215_sv2v_reg,mem_1214_sv2v_reg,mem_1213_sv2v_reg,
  mem_1212_sv2v_reg,mem_1211_sv2v_reg,mem_1210_sv2v_reg,mem_1209_sv2v_reg,mem_1208_sv2v_reg,
  mem_1207_sv2v_reg,mem_1206_sv2v_reg,mem_1205_sv2v_reg,mem_1204_sv2v_reg,
  mem_1203_sv2v_reg,mem_1202_sv2v_reg,mem_1201_sv2v_reg,mem_1200_sv2v_reg,
  mem_1199_sv2v_reg,mem_1198_sv2v_reg,mem_1197_sv2v_reg,mem_1196_sv2v_reg,mem_1195_sv2v_reg,
  mem_1194_sv2v_reg,mem_1193_sv2v_reg,mem_1192_sv2v_reg,mem_1191_sv2v_reg,
  mem_1190_sv2v_reg,mem_1189_sv2v_reg,mem_1188_sv2v_reg,mem_1187_sv2v_reg,mem_1186_sv2v_reg,
  mem_1185_sv2v_reg,mem_1184_sv2v_reg,mem_1183_sv2v_reg,mem_1182_sv2v_reg,
  mem_1181_sv2v_reg,mem_1180_sv2v_reg,mem_1179_sv2v_reg,mem_1178_sv2v_reg,mem_1177_sv2v_reg,
  mem_1176_sv2v_reg,mem_1175_sv2v_reg,mem_1174_sv2v_reg,mem_1173_sv2v_reg,
  mem_1172_sv2v_reg,mem_1171_sv2v_reg,mem_1170_sv2v_reg,mem_1169_sv2v_reg,mem_1168_sv2v_reg,
  mem_1167_sv2v_reg,mem_1166_sv2v_reg,mem_1165_sv2v_reg,mem_1164_sv2v_reg,
  mem_1163_sv2v_reg,mem_1162_sv2v_reg,mem_1161_sv2v_reg,mem_1160_sv2v_reg,
  mem_1159_sv2v_reg,mem_1158_sv2v_reg,mem_1157_sv2v_reg,mem_1156_sv2v_reg,mem_1155_sv2v_reg,
  mem_1154_sv2v_reg,mem_1153_sv2v_reg,mem_1152_sv2v_reg,mem_1151_sv2v_reg,
  mem_1150_sv2v_reg,mem_1149_sv2v_reg,mem_1148_sv2v_reg,mem_1147_sv2v_reg,mem_1146_sv2v_reg,
  mem_1145_sv2v_reg,mem_1144_sv2v_reg,mem_1143_sv2v_reg,mem_1142_sv2v_reg,
  mem_1141_sv2v_reg,mem_1140_sv2v_reg,mem_1139_sv2v_reg,mem_1138_sv2v_reg,mem_1137_sv2v_reg,
  mem_1136_sv2v_reg,mem_1135_sv2v_reg,mem_1134_sv2v_reg,mem_1133_sv2v_reg,
  mem_1132_sv2v_reg,mem_1131_sv2v_reg,mem_1130_sv2v_reg,mem_1129_sv2v_reg,mem_1128_sv2v_reg,
  mem_1127_sv2v_reg,mem_1126_sv2v_reg,mem_1125_sv2v_reg,mem_1124_sv2v_reg,
  mem_1123_sv2v_reg,mem_1122_sv2v_reg,mem_1121_sv2v_reg,mem_1120_sv2v_reg,
  mem_1119_sv2v_reg,mem_1118_sv2v_reg,mem_1117_sv2v_reg,mem_1116_sv2v_reg,mem_1115_sv2v_reg,
  mem_1114_sv2v_reg,mem_1113_sv2v_reg,mem_1112_sv2v_reg,mem_1111_sv2v_reg,
  mem_1110_sv2v_reg,mem_1109_sv2v_reg,mem_1108_sv2v_reg,mem_1107_sv2v_reg,mem_1106_sv2v_reg,
  mem_1105_sv2v_reg,mem_1104_sv2v_reg,mem_1103_sv2v_reg,mem_1102_sv2v_reg,
  mem_1101_sv2v_reg,mem_1100_sv2v_reg,mem_1099_sv2v_reg,mem_1098_sv2v_reg,mem_1097_sv2v_reg,
  mem_1096_sv2v_reg,mem_1095_sv2v_reg,mem_1094_sv2v_reg,mem_1093_sv2v_reg,
  mem_1092_sv2v_reg,mem_1091_sv2v_reg,mem_1090_sv2v_reg,mem_1089_sv2v_reg,mem_1088_sv2v_reg,
  mem_1087_sv2v_reg,mem_1086_sv2v_reg,mem_1085_sv2v_reg,mem_1084_sv2v_reg,
  mem_1083_sv2v_reg,mem_1082_sv2v_reg,mem_1081_sv2v_reg,mem_1080_sv2v_reg,
  mem_1079_sv2v_reg,mem_1078_sv2v_reg,mem_1077_sv2v_reg,mem_1076_sv2v_reg,mem_1075_sv2v_reg,
  mem_1074_sv2v_reg,mem_1073_sv2v_reg,mem_1072_sv2v_reg,mem_1071_sv2v_reg,
  mem_1070_sv2v_reg,mem_1069_sv2v_reg,mem_1068_sv2v_reg,mem_1067_sv2v_reg,mem_1066_sv2v_reg,
  mem_1065_sv2v_reg,mem_1064_sv2v_reg,mem_1063_sv2v_reg,mem_1062_sv2v_reg,
  mem_1061_sv2v_reg,mem_1060_sv2v_reg,mem_1059_sv2v_reg,mem_1058_sv2v_reg,mem_1057_sv2v_reg,
  mem_1056_sv2v_reg,mem_1055_sv2v_reg,mem_1054_sv2v_reg,mem_1053_sv2v_reg,
  mem_1052_sv2v_reg,mem_1051_sv2v_reg,mem_1050_sv2v_reg,mem_1049_sv2v_reg,mem_1048_sv2v_reg,
  mem_1047_sv2v_reg,mem_1046_sv2v_reg,mem_1045_sv2v_reg,mem_1044_sv2v_reg,
  mem_1043_sv2v_reg,mem_1042_sv2v_reg,mem_1041_sv2v_reg,mem_1040_sv2v_reg,
  mem_1039_sv2v_reg,mem_1038_sv2v_reg,mem_1037_sv2v_reg,mem_1036_sv2v_reg,mem_1035_sv2v_reg,
  mem_1034_sv2v_reg,mem_1033_sv2v_reg,mem_1032_sv2v_reg,mem_1031_sv2v_reg,
  mem_1030_sv2v_reg,mem_1029_sv2v_reg,mem_1028_sv2v_reg,mem_1027_sv2v_reg,mem_1026_sv2v_reg,
  mem_1025_sv2v_reg,mem_1024_sv2v_reg,mem_1023_sv2v_reg,mem_1022_sv2v_reg,
  mem_1021_sv2v_reg,mem_1020_sv2v_reg,mem_1019_sv2v_reg,mem_1018_sv2v_reg,mem_1017_sv2v_reg,
  mem_1016_sv2v_reg,mem_1015_sv2v_reg,mem_1014_sv2v_reg,mem_1013_sv2v_reg,
  mem_1012_sv2v_reg,mem_1011_sv2v_reg,mem_1010_sv2v_reg,mem_1009_sv2v_reg,mem_1008_sv2v_reg,
  mem_1007_sv2v_reg,mem_1006_sv2v_reg,mem_1005_sv2v_reg,mem_1004_sv2v_reg,
  mem_1003_sv2v_reg,mem_1002_sv2v_reg,mem_1001_sv2v_reg,mem_1000_sv2v_reg,
  mem_999_sv2v_reg,mem_998_sv2v_reg,mem_997_sv2v_reg,mem_996_sv2v_reg,mem_995_sv2v_reg,
  mem_994_sv2v_reg,mem_993_sv2v_reg,mem_992_sv2v_reg,mem_991_sv2v_reg,mem_990_sv2v_reg,
  mem_989_sv2v_reg,mem_988_sv2v_reg,mem_987_sv2v_reg,mem_986_sv2v_reg,mem_985_sv2v_reg,
  mem_984_sv2v_reg,mem_983_sv2v_reg,mem_982_sv2v_reg,mem_981_sv2v_reg,
  mem_980_sv2v_reg,mem_979_sv2v_reg,mem_978_sv2v_reg,mem_977_sv2v_reg,mem_976_sv2v_reg,
  mem_975_sv2v_reg,mem_974_sv2v_reg,mem_973_sv2v_reg,mem_972_sv2v_reg,mem_971_sv2v_reg,
  mem_970_sv2v_reg,mem_969_sv2v_reg,mem_968_sv2v_reg,mem_967_sv2v_reg,
  mem_966_sv2v_reg,mem_965_sv2v_reg,mem_964_sv2v_reg,mem_963_sv2v_reg,mem_962_sv2v_reg,
  mem_961_sv2v_reg,mem_960_sv2v_reg,mem_959_sv2v_reg,mem_958_sv2v_reg,mem_957_sv2v_reg,
  mem_956_sv2v_reg,mem_955_sv2v_reg,mem_954_sv2v_reg,mem_953_sv2v_reg,mem_952_sv2v_reg,
  mem_951_sv2v_reg,mem_950_sv2v_reg,mem_949_sv2v_reg,mem_948_sv2v_reg,
  mem_947_sv2v_reg,mem_946_sv2v_reg,mem_945_sv2v_reg,mem_944_sv2v_reg,mem_943_sv2v_reg,
  mem_942_sv2v_reg,mem_941_sv2v_reg,mem_940_sv2v_reg,mem_939_sv2v_reg,mem_938_sv2v_reg,
  mem_937_sv2v_reg,mem_936_sv2v_reg,mem_935_sv2v_reg,mem_934_sv2v_reg,
  mem_933_sv2v_reg,mem_932_sv2v_reg,mem_931_sv2v_reg,mem_930_sv2v_reg,mem_929_sv2v_reg,
  mem_928_sv2v_reg,mem_927_sv2v_reg,mem_926_sv2v_reg,mem_925_sv2v_reg,mem_924_sv2v_reg,
  mem_923_sv2v_reg,mem_922_sv2v_reg,mem_921_sv2v_reg,mem_920_sv2v_reg,
  mem_919_sv2v_reg,mem_918_sv2v_reg,mem_917_sv2v_reg,mem_916_sv2v_reg,mem_915_sv2v_reg,
  mem_914_sv2v_reg,mem_913_sv2v_reg,mem_912_sv2v_reg,mem_911_sv2v_reg,mem_910_sv2v_reg,
  mem_909_sv2v_reg,mem_908_sv2v_reg,mem_907_sv2v_reg,mem_906_sv2v_reg,mem_905_sv2v_reg,
  mem_904_sv2v_reg,mem_903_sv2v_reg,mem_902_sv2v_reg,mem_901_sv2v_reg,
  mem_900_sv2v_reg,mem_899_sv2v_reg,mem_898_sv2v_reg,mem_897_sv2v_reg,mem_896_sv2v_reg,
  mem_895_sv2v_reg,mem_894_sv2v_reg,mem_893_sv2v_reg,mem_892_sv2v_reg,mem_891_sv2v_reg,
  mem_890_sv2v_reg,mem_889_sv2v_reg,mem_888_sv2v_reg,mem_887_sv2v_reg,
  mem_886_sv2v_reg,mem_885_sv2v_reg,mem_884_sv2v_reg,mem_883_sv2v_reg,mem_882_sv2v_reg,
  mem_881_sv2v_reg,mem_880_sv2v_reg,mem_879_sv2v_reg,mem_878_sv2v_reg,mem_877_sv2v_reg,
  mem_876_sv2v_reg,mem_875_sv2v_reg,mem_874_sv2v_reg,mem_873_sv2v_reg,mem_872_sv2v_reg,
  mem_871_sv2v_reg,mem_870_sv2v_reg,mem_869_sv2v_reg,mem_868_sv2v_reg,
  mem_867_sv2v_reg,mem_866_sv2v_reg,mem_865_sv2v_reg,mem_864_sv2v_reg,mem_863_sv2v_reg,
  mem_862_sv2v_reg,mem_861_sv2v_reg,mem_860_sv2v_reg,mem_859_sv2v_reg,mem_858_sv2v_reg,
  mem_857_sv2v_reg,mem_856_sv2v_reg,mem_855_sv2v_reg,mem_854_sv2v_reg,
  mem_853_sv2v_reg,mem_852_sv2v_reg,mem_851_sv2v_reg,mem_850_sv2v_reg,mem_849_sv2v_reg,
  mem_848_sv2v_reg,mem_847_sv2v_reg,mem_846_sv2v_reg,mem_845_sv2v_reg,mem_844_sv2v_reg,
  mem_843_sv2v_reg,mem_842_sv2v_reg,mem_841_sv2v_reg,mem_840_sv2v_reg,
  mem_839_sv2v_reg,mem_838_sv2v_reg,mem_837_sv2v_reg,mem_836_sv2v_reg,mem_835_sv2v_reg,
  mem_834_sv2v_reg,mem_833_sv2v_reg,mem_832_sv2v_reg,mem_831_sv2v_reg,mem_830_sv2v_reg,
  mem_829_sv2v_reg,mem_828_sv2v_reg,mem_827_sv2v_reg,mem_826_sv2v_reg,mem_825_sv2v_reg,
  mem_824_sv2v_reg,mem_823_sv2v_reg,mem_822_sv2v_reg,mem_821_sv2v_reg,
  mem_820_sv2v_reg,mem_819_sv2v_reg,mem_818_sv2v_reg,mem_817_sv2v_reg,mem_816_sv2v_reg,
  mem_815_sv2v_reg,mem_814_sv2v_reg,mem_813_sv2v_reg,mem_812_sv2v_reg,mem_811_sv2v_reg,
  mem_810_sv2v_reg,mem_809_sv2v_reg,mem_808_sv2v_reg,mem_807_sv2v_reg,
  mem_806_sv2v_reg,mem_805_sv2v_reg,mem_804_sv2v_reg,mem_803_sv2v_reg,mem_802_sv2v_reg,
  mem_801_sv2v_reg,mem_800_sv2v_reg,mem_799_sv2v_reg,mem_798_sv2v_reg,mem_797_sv2v_reg,
  mem_796_sv2v_reg,mem_795_sv2v_reg,mem_794_sv2v_reg,mem_793_sv2v_reg,mem_792_sv2v_reg,
  mem_791_sv2v_reg,mem_790_sv2v_reg,mem_789_sv2v_reg,mem_788_sv2v_reg,
  mem_787_sv2v_reg,mem_786_sv2v_reg,mem_785_sv2v_reg,mem_784_sv2v_reg,mem_783_sv2v_reg,
  mem_782_sv2v_reg,mem_781_sv2v_reg,mem_780_sv2v_reg,mem_779_sv2v_reg,mem_778_sv2v_reg,
  mem_777_sv2v_reg,mem_776_sv2v_reg,mem_775_sv2v_reg,mem_774_sv2v_reg,
  mem_773_sv2v_reg,mem_772_sv2v_reg,mem_771_sv2v_reg,mem_770_sv2v_reg,mem_769_sv2v_reg,
  mem_768_sv2v_reg,mem_767_sv2v_reg,mem_766_sv2v_reg,mem_765_sv2v_reg,mem_764_sv2v_reg,
  mem_763_sv2v_reg,mem_762_sv2v_reg,mem_761_sv2v_reg,mem_760_sv2v_reg,
  mem_759_sv2v_reg,mem_758_sv2v_reg,mem_757_sv2v_reg,mem_756_sv2v_reg,mem_755_sv2v_reg,
  mem_754_sv2v_reg,mem_753_sv2v_reg,mem_752_sv2v_reg,mem_751_sv2v_reg,mem_750_sv2v_reg,
  mem_749_sv2v_reg,mem_748_sv2v_reg,mem_747_sv2v_reg,mem_746_sv2v_reg,mem_745_sv2v_reg,
  mem_744_sv2v_reg,mem_743_sv2v_reg,mem_742_sv2v_reg,mem_741_sv2v_reg,
  mem_740_sv2v_reg,mem_739_sv2v_reg,mem_738_sv2v_reg,mem_737_sv2v_reg,mem_736_sv2v_reg,
  mem_735_sv2v_reg,mem_734_sv2v_reg,mem_733_sv2v_reg,mem_732_sv2v_reg,mem_731_sv2v_reg,
  mem_730_sv2v_reg,mem_729_sv2v_reg,mem_728_sv2v_reg,mem_727_sv2v_reg,
  mem_726_sv2v_reg,mem_725_sv2v_reg,mem_724_sv2v_reg,mem_723_sv2v_reg,mem_722_sv2v_reg,
  mem_721_sv2v_reg,mem_720_sv2v_reg,mem_719_sv2v_reg,mem_718_sv2v_reg,mem_717_sv2v_reg,
  mem_716_sv2v_reg,mem_715_sv2v_reg,mem_714_sv2v_reg,mem_713_sv2v_reg,mem_712_sv2v_reg,
  mem_711_sv2v_reg,mem_710_sv2v_reg,mem_709_sv2v_reg,mem_708_sv2v_reg,
  mem_707_sv2v_reg,mem_706_sv2v_reg,mem_705_sv2v_reg,mem_704_sv2v_reg,mem_703_sv2v_reg,
  mem_702_sv2v_reg,mem_701_sv2v_reg,mem_700_sv2v_reg,mem_699_sv2v_reg,mem_698_sv2v_reg,
  mem_697_sv2v_reg,mem_696_sv2v_reg,mem_695_sv2v_reg,mem_694_sv2v_reg,
  mem_693_sv2v_reg,mem_692_sv2v_reg,mem_691_sv2v_reg,mem_690_sv2v_reg,mem_689_sv2v_reg,
  mem_688_sv2v_reg,mem_687_sv2v_reg,mem_686_sv2v_reg,mem_685_sv2v_reg,mem_684_sv2v_reg,
  mem_683_sv2v_reg,mem_682_sv2v_reg,mem_681_sv2v_reg,mem_680_sv2v_reg,
  mem_679_sv2v_reg,mem_678_sv2v_reg,mem_677_sv2v_reg,mem_676_sv2v_reg,mem_675_sv2v_reg,
  mem_674_sv2v_reg,mem_673_sv2v_reg,mem_672_sv2v_reg,mem_671_sv2v_reg,mem_670_sv2v_reg,
  mem_669_sv2v_reg,mem_668_sv2v_reg,mem_667_sv2v_reg,mem_666_sv2v_reg,mem_665_sv2v_reg,
  mem_664_sv2v_reg,mem_663_sv2v_reg,mem_662_sv2v_reg,mem_661_sv2v_reg,
  mem_660_sv2v_reg,mem_659_sv2v_reg,mem_658_sv2v_reg,mem_657_sv2v_reg,mem_656_sv2v_reg,
  mem_655_sv2v_reg,mem_654_sv2v_reg,mem_653_sv2v_reg,mem_652_sv2v_reg,mem_651_sv2v_reg,
  mem_650_sv2v_reg,mem_649_sv2v_reg,mem_648_sv2v_reg,mem_647_sv2v_reg,
  mem_646_sv2v_reg,mem_645_sv2v_reg,mem_644_sv2v_reg,mem_643_sv2v_reg,mem_642_sv2v_reg,
  mem_641_sv2v_reg,mem_640_sv2v_reg,mem_639_sv2v_reg,mem_638_sv2v_reg,mem_637_sv2v_reg,
  mem_636_sv2v_reg,mem_635_sv2v_reg,mem_634_sv2v_reg,mem_633_sv2v_reg,mem_632_sv2v_reg,
  mem_631_sv2v_reg,mem_630_sv2v_reg,mem_629_sv2v_reg,mem_628_sv2v_reg,
  mem_627_sv2v_reg,mem_626_sv2v_reg,mem_625_sv2v_reg,mem_624_sv2v_reg,mem_623_sv2v_reg,
  mem_622_sv2v_reg,mem_621_sv2v_reg,mem_620_sv2v_reg,mem_619_sv2v_reg,mem_618_sv2v_reg,
  mem_617_sv2v_reg,mem_616_sv2v_reg,mem_615_sv2v_reg,mem_614_sv2v_reg,
  mem_613_sv2v_reg,mem_612_sv2v_reg,mem_611_sv2v_reg,mem_610_sv2v_reg,mem_609_sv2v_reg,
  mem_608_sv2v_reg,mem_607_sv2v_reg,mem_606_sv2v_reg,mem_605_sv2v_reg,mem_604_sv2v_reg,
  mem_603_sv2v_reg,mem_602_sv2v_reg,mem_601_sv2v_reg,mem_600_sv2v_reg,
  mem_599_sv2v_reg,mem_598_sv2v_reg,mem_597_sv2v_reg,mem_596_sv2v_reg,mem_595_sv2v_reg,
  mem_594_sv2v_reg,mem_593_sv2v_reg,mem_592_sv2v_reg,mem_591_sv2v_reg,mem_590_sv2v_reg,
  mem_589_sv2v_reg,mem_588_sv2v_reg,mem_587_sv2v_reg,mem_586_sv2v_reg,mem_585_sv2v_reg,
  mem_584_sv2v_reg,mem_583_sv2v_reg,mem_582_sv2v_reg,mem_581_sv2v_reg,
  mem_580_sv2v_reg,mem_579_sv2v_reg,mem_578_sv2v_reg,mem_577_sv2v_reg,mem_576_sv2v_reg,
  mem_575_sv2v_reg,mem_574_sv2v_reg,mem_573_sv2v_reg,mem_572_sv2v_reg,mem_571_sv2v_reg,
  mem_570_sv2v_reg,mem_569_sv2v_reg,mem_568_sv2v_reg,mem_567_sv2v_reg,
  mem_566_sv2v_reg,mem_565_sv2v_reg,mem_564_sv2v_reg,mem_563_sv2v_reg,mem_562_sv2v_reg,
  mem_561_sv2v_reg,mem_560_sv2v_reg,mem_559_sv2v_reg,mem_558_sv2v_reg,mem_557_sv2v_reg,
  mem_556_sv2v_reg,mem_555_sv2v_reg,mem_554_sv2v_reg,mem_553_sv2v_reg,mem_552_sv2v_reg,
  mem_551_sv2v_reg,mem_550_sv2v_reg,mem_549_sv2v_reg,mem_548_sv2v_reg,
  mem_547_sv2v_reg,mem_546_sv2v_reg,mem_545_sv2v_reg,mem_544_sv2v_reg,mem_543_sv2v_reg,
  mem_542_sv2v_reg,mem_541_sv2v_reg,mem_540_sv2v_reg,mem_539_sv2v_reg,mem_538_sv2v_reg,
  mem_537_sv2v_reg,mem_536_sv2v_reg,mem_535_sv2v_reg,mem_534_sv2v_reg,
  mem_533_sv2v_reg,mem_532_sv2v_reg,mem_531_sv2v_reg,mem_530_sv2v_reg,mem_529_sv2v_reg,
  mem_528_sv2v_reg,mem_527_sv2v_reg,mem_526_sv2v_reg,mem_525_sv2v_reg,mem_524_sv2v_reg,
  mem_523_sv2v_reg,mem_522_sv2v_reg,mem_521_sv2v_reg,mem_520_sv2v_reg,
  mem_519_sv2v_reg,mem_518_sv2v_reg,mem_517_sv2v_reg,mem_516_sv2v_reg,mem_515_sv2v_reg,
  mem_514_sv2v_reg,mem_513_sv2v_reg,mem_512_sv2v_reg,mem_511_sv2v_reg,mem_510_sv2v_reg,
  mem_509_sv2v_reg,mem_508_sv2v_reg,mem_507_sv2v_reg,mem_506_sv2v_reg,mem_505_sv2v_reg,
  mem_504_sv2v_reg,mem_503_sv2v_reg,mem_502_sv2v_reg,mem_501_sv2v_reg,
  mem_500_sv2v_reg,mem_499_sv2v_reg,mem_498_sv2v_reg,mem_497_sv2v_reg,mem_496_sv2v_reg,
  mem_495_sv2v_reg,mem_494_sv2v_reg,mem_493_sv2v_reg,mem_492_sv2v_reg,mem_491_sv2v_reg,
  mem_490_sv2v_reg,mem_489_sv2v_reg,mem_488_sv2v_reg,mem_487_sv2v_reg,
  mem_486_sv2v_reg,mem_485_sv2v_reg,mem_484_sv2v_reg,mem_483_sv2v_reg,mem_482_sv2v_reg,
  mem_481_sv2v_reg,mem_480_sv2v_reg,mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,
  mem_476_sv2v_reg,mem_475_sv2v_reg,mem_474_sv2v_reg,mem_473_sv2v_reg,mem_472_sv2v_reg,
  mem_471_sv2v_reg,mem_470_sv2v_reg,mem_469_sv2v_reg,mem_468_sv2v_reg,
  mem_467_sv2v_reg,mem_466_sv2v_reg,mem_465_sv2v_reg,mem_464_sv2v_reg,mem_463_sv2v_reg,
  mem_462_sv2v_reg,mem_461_sv2v_reg,mem_460_sv2v_reg,mem_459_sv2v_reg,mem_458_sv2v_reg,
  mem_457_sv2v_reg,mem_456_sv2v_reg,mem_455_sv2v_reg,mem_454_sv2v_reg,
  mem_453_sv2v_reg,mem_452_sv2v_reg,mem_451_sv2v_reg,mem_450_sv2v_reg,mem_449_sv2v_reg,
  mem_448_sv2v_reg,mem_447_sv2v_reg,mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,
  mem_443_sv2v_reg,mem_442_sv2v_reg,mem_441_sv2v_reg,mem_440_sv2v_reg,
  mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,mem_436_sv2v_reg,mem_435_sv2v_reg,
  mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,mem_431_sv2v_reg,mem_430_sv2v_reg,
  mem_429_sv2v_reg,mem_428_sv2v_reg,mem_427_sv2v_reg,mem_426_sv2v_reg,mem_425_sv2v_reg,
  mem_424_sv2v_reg,mem_423_sv2v_reg,mem_422_sv2v_reg,mem_421_sv2v_reg,
  mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,mem_417_sv2v_reg,mem_416_sv2v_reg,
  mem_415_sv2v_reg,mem_414_sv2v_reg,mem_413_sv2v_reg,mem_412_sv2v_reg,mem_411_sv2v_reg,
  mem_410_sv2v_reg,mem_409_sv2v_reg,mem_408_sv2v_reg,mem_407_sv2v_reg,
  mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,mem_403_sv2v_reg,mem_402_sv2v_reg,
  mem_401_sv2v_reg,mem_400_sv2v_reg,mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,
  mem_396_sv2v_reg,mem_395_sv2v_reg,mem_394_sv2v_reg,mem_393_sv2v_reg,mem_392_sv2v_reg,
  mem_391_sv2v_reg,mem_390_sv2v_reg,mem_389_sv2v_reg,mem_388_sv2v_reg,
  mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,mem_384_sv2v_reg,mem_383_sv2v_reg,
  mem_382_sv2v_reg,mem_381_sv2v_reg,mem_380_sv2v_reg,mem_379_sv2v_reg,mem_378_sv2v_reg,
  mem_377_sv2v_reg,mem_376_sv2v_reg,mem_375_sv2v_reg,mem_374_sv2v_reg,
  mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,mem_370_sv2v_reg,mem_369_sv2v_reg,
  mem_368_sv2v_reg,mem_367_sv2v_reg,mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,
  mem_363_sv2v_reg,mem_362_sv2v_reg,mem_361_sv2v_reg,mem_360_sv2v_reg,
  mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,mem_356_sv2v_reg,mem_355_sv2v_reg,
  mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,mem_351_sv2v_reg,mem_350_sv2v_reg,
  mem_349_sv2v_reg,mem_348_sv2v_reg,mem_347_sv2v_reg,mem_346_sv2v_reg,mem_345_sv2v_reg,
  mem_344_sv2v_reg,mem_343_sv2v_reg,mem_342_sv2v_reg,mem_341_sv2v_reg,
  mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,mem_337_sv2v_reg,mem_336_sv2v_reg,
  mem_335_sv2v_reg,mem_334_sv2v_reg,mem_333_sv2v_reg,mem_332_sv2v_reg,mem_331_sv2v_reg,
  mem_330_sv2v_reg,mem_329_sv2v_reg,mem_328_sv2v_reg,mem_327_sv2v_reg,
  mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,mem_323_sv2v_reg,mem_322_sv2v_reg,
  mem_321_sv2v_reg,mem_320_sv2v_reg,mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,
  mem_316_sv2v_reg,mem_315_sv2v_reg,mem_314_sv2v_reg,mem_313_sv2v_reg,mem_312_sv2v_reg,
  mem_311_sv2v_reg,mem_310_sv2v_reg,mem_309_sv2v_reg,mem_308_sv2v_reg,
  mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,mem_304_sv2v_reg,mem_303_sv2v_reg,
  mem_302_sv2v_reg,mem_301_sv2v_reg,mem_300_sv2v_reg,mem_299_sv2v_reg,mem_298_sv2v_reg,
  mem_297_sv2v_reg,mem_296_sv2v_reg,mem_295_sv2v_reg,mem_294_sv2v_reg,
  mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,mem_290_sv2v_reg,mem_289_sv2v_reg,
  mem_288_sv2v_reg,mem_287_sv2v_reg,mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,
  mem_283_sv2v_reg,mem_282_sv2v_reg,mem_281_sv2v_reg,mem_280_sv2v_reg,
  mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,mem_276_sv2v_reg,mem_275_sv2v_reg,
  mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,mem_271_sv2v_reg,mem_270_sv2v_reg,
  mem_269_sv2v_reg,mem_268_sv2v_reg,mem_267_sv2v_reg,mem_266_sv2v_reg,mem_265_sv2v_reg,
  mem_264_sv2v_reg,mem_263_sv2v_reg,mem_262_sv2v_reg,mem_261_sv2v_reg,
  mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,mem_257_sv2v_reg,mem_256_sv2v_reg,
  mem_255_sv2v_reg,mem_254_sv2v_reg,mem_253_sv2v_reg,mem_252_sv2v_reg,mem_251_sv2v_reg,
  mem_250_sv2v_reg,mem_249_sv2v_reg,mem_248_sv2v_reg,mem_247_sv2v_reg,
  mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,mem_243_sv2v_reg,mem_242_sv2v_reg,
  mem_241_sv2v_reg,mem_240_sv2v_reg,mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,
  mem_236_sv2v_reg,mem_235_sv2v_reg,mem_234_sv2v_reg,mem_233_sv2v_reg,mem_232_sv2v_reg,
  mem_231_sv2v_reg,mem_230_sv2v_reg,mem_229_sv2v_reg,mem_228_sv2v_reg,
  mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,mem_224_sv2v_reg,mem_223_sv2v_reg,
  mem_222_sv2v_reg,mem_221_sv2v_reg,mem_220_sv2v_reg,mem_219_sv2v_reg,mem_218_sv2v_reg,
  mem_217_sv2v_reg,mem_216_sv2v_reg,mem_215_sv2v_reg,mem_214_sv2v_reg,
  mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,mem_210_sv2v_reg,mem_209_sv2v_reg,
  mem_208_sv2v_reg,mem_207_sv2v_reg,mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,
  mem_203_sv2v_reg,mem_202_sv2v_reg,mem_201_sv2v_reg,mem_200_sv2v_reg,
  mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,mem_196_sv2v_reg,mem_195_sv2v_reg,
  mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,mem_191_sv2v_reg,mem_190_sv2v_reg,
  mem_189_sv2v_reg,mem_188_sv2v_reg,mem_187_sv2v_reg,mem_186_sv2v_reg,mem_185_sv2v_reg,
  mem_184_sv2v_reg,mem_183_sv2v_reg,mem_182_sv2v_reg,mem_181_sv2v_reg,
  mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,mem_177_sv2v_reg,mem_176_sv2v_reg,
  mem_175_sv2v_reg,mem_174_sv2v_reg,mem_173_sv2v_reg,mem_172_sv2v_reg,mem_171_sv2v_reg,
  mem_170_sv2v_reg,mem_169_sv2v_reg,mem_168_sv2v_reg,mem_167_sv2v_reg,
  mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,mem_163_sv2v_reg,mem_162_sv2v_reg,
  mem_161_sv2v_reg,mem_160_sv2v_reg,mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,
  mem_156_sv2v_reg,mem_155_sv2v_reg,mem_154_sv2v_reg,mem_153_sv2v_reg,mem_152_sv2v_reg,
  mem_151_sv2v_reg,mem_150_sv2v_reg,mem_149_sv2v_reg,mem_148_sv2v_reg,
  mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,mem_144_sv2v_reg,mem_143_sv2v_reg,
  mem_142_sv2v_reg,mem_141_sv2v_reg,mem_140_sv2v_reg,mem_139_sv2v_reg,mem_138_sv2v_reg,
  mem_137_sv2v_reg,mem_136_sv2v_reg,mem_135_sv2v_reg,mem_134_sv2v_reg,
  mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,mem_130_sv2v_reg,mem_129_sv2v_reg,
  mem_128_sv2v_reg,mem_127_sv2v_reg,mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,
  mem_123_sv2v_reg,mem_122_sv2v_reg,mem_121_sv2v_reg,mem_120_sv2v_reg,
  mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,mem_116_sv2v_reg,mem_115_sv2v_reg,
  mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,mem_111_sv2v_reg,mem_110_sv2v_reg,
  mem_109_sv2v_reg,mem_108_sv2v_reg,mem_107_sv2v_reg,mem_106_sv2v_reg,mem_105_sv2v_reg,
  mem_104_sv2v_reg,mem_103_sv2v_reg,mem_102_sv2v_reg,mem_101_sv2v_reg,
  mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,mem_97_sv2v_reg,mem_96_sv2v_reg,
  mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,mem_92_sv2v_reg,mem_91_sv2v_reg,
  mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,mem_87_sv2v_reg,mem_86_sv2v_reg,
  mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,mem_82_sv2v_reg,mem_81_sv2v_reg,
  mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,mem_77_sv2v_reg,mem_76_sv2v_reg,
  mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,mem_72_sv2v_reg,mem_71_sv2v_reg,
  mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,mem_67_sv2v_reg,mem_66_sv2v_reg,
  mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,
  mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,
  mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,
  mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,
  mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,
  mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,
  mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,
  mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,
  mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,
  mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,
  mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,
  mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,
  mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[3967] = mem_3967_sv2v_reg;
  assign mem[3966] = mem_3966_sv2v_reg;
  assign mem[3965] = mem_3965_sv2v_reg;
  assign mem[3964] = mem_3964_sv2v_reg;
  assign mem[3963] = mem_3963_sv2v_reg;
  assign mem[3962] = mem_3962_sv2v_reg;
  assign mem[3961] = mem_3961_sv2v_reg;
  assign mem[3960] = mem_3960_sv2v_reg;
  assign mem[3959] = mem_3959_sv2v_reg;
  assign mem[3958] = mem_3958_sv2v_reg;
  assign mem[3957] = mem_3957_sv2v_reg;
  assign mem[3956] = mem_3956_sv2v_reg;
  assign mem[3955] = mem_3955_sv2v_reg;
  assign mem[3954] = mem_3954_sv2v_reg;
  assign mem[3953] = mem_3953_sv2v_reg;
  assign mem[3952] = mem_3952_sv2v_reg;
  assign mem[3951] = mem_3951_sv2v_reg;
  assign mem[3950] = mem_3950_sv2v_reg;
  assign mem[3949] = mem_3949_sv2v_reg;
  assign mem[3948] = mem_3948_sv2v_reg;
  assign mem[3947] = mem_3947_sv2v_reg;
  assign mem[3946] = mem_3946_sv2v_reg;
  assign mem[3945] = mem_3945_sv2v_reg;
  assign mem[3944] = mem_3944_sv2v_reg;
  assign mem[3943] = mem_3943_sv2v_reg;
  assign mem[3942] = mem_3942_sv2v_reg;
  assign mem[3941] = mem_3941_sv2v_reg;
  assign mem[3940] = mem_3940_sv2v_reg;
  assign mem[3939] = mem_3939_sv2v_reg;
  assign mem[3938] = mem_3938_sv2v_reg;
  assign mem[3937] = mem_3937_sv2v_reg;
  assign mem[3936] = mem_3936_sv2v_reg;
  assign mem[3935] = mem_3935_sv2v_reg;
  assign mem[3934] = mem_3934_sv2v_reg;
  assign mem[3933] = mem_3933_sv2v_reg;
  assign mem[3932] = mem_3932_sv2v_reg;
  assign mem[3931] = mem_3931_sv2v_reg;
  assign mem[3930] = mem_3930_sv2v_reg;
  assign mem[3929] = mem_3929_sv2v_reg;
  assign mem[3928] = mem_3928_sv2v_reg;
  assign mem[3927] = mem_3927_sv2v_reg;
  assign mem[3926] = mem_3926_sv2v_reg;
  assign mem[3925] = mem_3925_sv2v_reg;
  assign mem[3924] = mem_3924_sv2v_reg;
  assign mem[3923] = mem_3923_sv2v_reg;
  assign mem[3922] = mem_3922_sv2v_reg;
  assign mem[3921] = mem_3921_sv2v_reg;
  assign mem[3920] = mem_3920_sv2v_reg;
  assign mem[3919] = mem_3919_sv2v_reg;
  assign mem[3918] = mem_3918_sv2v_reg;
  assign mem[3917] = mem_3917_sv2v_reg;
  assign mem[3916] = mem_3916_sv2v_reg;
  assign mem[3915] = mem_3915_sv2v_reg;
  assign mem[3914] = mem_3914_sv2v_reg;
  assign mem[3913] = mem_3913_sv2v_reg;
  assign mem[3912] = mem_3912_sv2v_reg;
  assign mem[3911] = mem_3911_sv2v_reg;
  assign mem[3910] = mem_3910_sv2v_reg;
  assign mem[3909] = mem_3909_sv2v_reg;
  assign mem[3908] = mem_3908_sv2v_reg;
  assign mem[3907] = mem_3907_sv2v_reg;
  assign mem[3906] = mem_3906_sv2v_reg;
  assign mem[3905] = mem_3905_sv2v_reg;
  assign mem[3904] = mem_3904_sv2v_reg;
  assign mem[3903] = mem_3903_sv2v_reg;
  assign mem[3902] = mem_3902_sv2v_reg;
  assign mem[3901] = mem_3901_sv2v_reg;
  assign mem[3900] = mem_3900_sv2v_reg;
  assign mem[3899] = mem_3899_sv2v_reg;
  assign mem[3898] = mem_3898_sv2v_reg;
  assign mem[3897] = mem_3897_sv2v_reg;
  assign mem[3896] = mem_3896_sv2v_reg;
  assign mem[3895] = mem_3895_sv2v_reg;
  assign mem[3894] = mem_3894_sv2v_reg;
  assign mem[3893] = mem_3893_sv2v_reg;
  assign mem[3892] = mem_3892_sv2v_reg;
  assign mem[3891] = mem_3891_sv2v_reg;
  assign mem[3890] = mem_3890_sv2v_reg;
  assign mem[3889] = mem_3889_sv2v_reg;
  assign mem[3888] = mem_3888_sv2v_reg;
  assign mem[3887] = mem_3887_sv2v_reg;
  assign mem[3886] = mem_3886_sv2v_reg;
  assign mem[3885] = mem_3885_sv2v_reg;
  assign mem[3884] = mem_3884_sv2v_reg;
  assign mem[3883] = mem_3883_sv2v_reg;
  assign mem[3882] = mem_3882_sv2v_reg;
  assign mem[3881] = mem_3881_sv2v_reg;
  assign mem[3880] = mem_3880_sv2v_reg;
  assign mem[3879] = mem_3879_sv2v_reg;
  assign mem[3878] = mem_3878_sv2v_reg;
  assign mem[3877] = mem_3877_sv2v_reg;
  assign mem[3876] = mem_3876_sv2v_reg;
  assign mem[3875] = mem_3875_sv2v_reg;
  assign mem[3874] = mem_3874_sv2v_reg;
  assign mem[3873] = mem_3873_sv2v_reg;
  assign mem[3872] = mem_3872_sv2v_reg;
  assign mem[3871] = mem_3871_sv2v_reg;
  assign mem[3870] = mem_3870_sv2v_reg;
  assign mem[3869] = mem_3869_sv2v_reg;
  assign mem[3868] = mem_3868_sv2v_reg;
  assign mem[3867] = mem_3867_sv2v_reg;
  assign mem[3866] = mem_3866_sv2v_reg;
  assign mem[3865] = mem_3865_sv2v_reg;
  assign mem[3864] = mem_3864_sv2v_reg;
  assign mem[3863] = mem_3863_sv2v_reg;
  assign mem[3862] = mem_3862_sv2v_reg;
  assign mem[3861] = mem_3861_sv2v_reg;
  assign mem[3860] = mem_3860_sv2v_reg;
  assign mem[3859] = mem_3859_sv2v_reg;
  assign mem[3858] = mem_3858_sv2v_reg;
  assign mem[3857] = mem_3857_sv2v_reg;
  assign mem[3856] = mem_3856_sv2v_reg;
  assign mem[3855] = mem_3855_sv2v_reg;
  assign mem[3854] = mem_3854_sv2v_reg;
  assign mem[3853] = mem_3853_sv2v_reg;
  assign mem[3852] = mem_3852_sv2v_reg;
  assign mem[3851] = mem_3851_sv2v_reg;
  assign mem[3850] = mem_3850_sv2v_reg;
  assign mem[3849] = mem_3849_sv2v_reg;
  assign mem[3848] = mem_3848_sv2v_reg;
  assign mem[3847] = mem_3847_sv2v_reg;
  assign mem[3846] = mem_3846_sv2v_reg;
  assign mem[3845] = mem_3845_sv2v_reg;
  assign mem[3844] = mem_3844_sv2v_reg;
  assign mem[3843] = mem_3843_sv2v_reg;
  assign mem[3842] = mem_3842_sv2v_reg;
  assign mem[3841] = mem_3841_sv2v_reg;
  assign mem[3840] = mem_3840_sv2v_reg;
  assign mem[3839] = mem_3839_sv2v_reg;
  assign mem[3838] = mem_3838_sv2v_reg;
  assign mem[3837] = mem_3837_sv2v_reg;
  assign mem[3836] = mem_3836_sv2v_reg;
  assign mem[3835] = mem_3835_sv2v_reg;
  assign mem[3834] = mem_3834_sv2v_reg;
  assign mem[3833] = mem_3833_sv2v_reg;
  assign mem[3832] = mem_3832_sv2v_reg;
  assign mem[3831] = mem_3831_sv2v_reg;
  assign mem[3830] = mem_3830_sv2v_reg;
  assign mem[3829] = mem_3829_sv2v_reg;
  assign mem[3828] = mem_3828_sv2v_reg;
  assign mem[3827] = mem_3827_sv2v_reg;
  assign mem[3826] = mem_3826_sv2v_reg;
  assign mem[3825] = mem_3825_sv2v_reg;
  assign mem[3824] = mem_3824_sv2v_reg;
  assign mem[3823] = mem_3823_sv2v_reg;
  assign mem[3822] = mem_3822_sv2v_reg;
  assign mem[3821] = mem_3821_sv2v_reg;
  assign mem[3820] = mem_3820_sv2v_reg;
  assign mem[3819] = mem_3819_sv2v_reg;
  assign mem[3818] = mem_3818_sv2v_reg;
  assign mem[3817] = mem_3817_sv2v_reg;
  assign mem[3816] = mem_3816_sv2v_reg;
  assign mem[3815] = mem_3815_sv2v_reg;
  assign mem[3814] = mem_3814_sv2v_reg;
  assign mem[3813] = mem_3813_sv2v_reg;
  assign mem[3812] = mem_3812_sv2v_reg;
  assign mem[3811] = mem_3811_sv2v_reg;
  assign mem[3810] = mem_3810_sv2v_reg;
  assign mem[3809] = mem_3809_sv2v_reg;
  assign mem[3808] = mem_3808_sv2v_reg;
  assign mem[3807] = mem_3807_sv2v_reg;
  assign mem[3806] = mem_3806_sv2v_reg;
  assign mem[3805] = mem_3805_sv2v_reg;
  assign mem[3804] = mem_3804_sv2v_reg;
  assign mem[3803] = mem_3803_sv2v_reg;
  assign mem[3802] = mem_3802_sv2v_reg;
  assign mem[3801] = mem_3801_sv2v_reg;
  assign mem[3800] = mem_3800_sv2v_reg;
  assign mem[3799] = mem_3799_sv2v_reg;
  assign mem[3798] = mem_3798_sv2v_reg;
  assign mem[3797] = mem_3797_sv2v_reg;
  assign mem[3796] = mem_3796_sv2v_reg;
  assign mem[3795] = mem_3795_sv2v_reg;
  assign mem[3794] = mem_3794_sv2v_reg;
  assign mem[3793] = mem_3793_sv2v_reg;
  assign mem[3792] = mem_3792_sv2v_reg;
  assign mem[3791] = mem_3791_sv2v_reg;
  assign mem[3790] = mem_3790_sv2v_reg;
  assign mem[3789] = mem_3789_sv2v_reg;
  assign mem[3788] = mem_3788_sv2v_reg;
  assign mem[3787] = mem_3787_sv2v_reg;
  assign mem[3786] = mem_3786_sv2v_reg;
  assign mem[3785] = mem_3785_sv2v_reg;
  assign mem[3784] = mem_3784_sv2v_reg;
  assign mem[3783] = mem_3783_sv2v_reg;
  assign mem[3782] = mem_3782_sv2v_reg;
  assign mem[3781] = mem_3781_sv2v_reg;
  assign mem[3780] = mem_3780_sv2v_reg;
  assign mem[3779] = mem_3779_sv2v_reg;
  assign mem[3778] = mem_3778_sv2v_reg;
  assign mem[3777] = mem_3777_sv2v_reg;
  assign mem[3776] = mem_3776_sv2v_reg;
  assign mem[3775] = mem_3775_sv2v_reg;
  assign mem[3774] = mem_3774_sv2v_reg;
  assign mem[3773] = mem_3773_sv2v_reg;
  assign mem[3772] = mem_3772_sv2v_reg;
  assign mem[3771] = mem_3771_sv2v_reg;
  assign mem[3770] = mem_3770_sv2v_reg;
  assign mem[3769] = mem_3769_sv2v_reg;
  assign mem[3768] = mem_3768_sv2v_reg;
  assign mem[3767] = mem_3767_sv2v_reg;
  assign mem[3766] = mem_3766_sv2v_reg;
  assign mem[3765] = mem_3765_sv2v_reg;
  assign mem[3764] = mem_3764_sv2v_reg;
  assign mem[3763] = mem_3763_sv2v_reg;
  assign mem[3762] = mem_3762_sv2v_reg;
  assign mem[3761] = mem_3761_sv2v_reg;
  assign mem[3760] = mem_3760_sv2v_reg;
  assign mem[3759] = mem_3759_sv2v_reg;
  assign mem[3758] = mem_3758_sv2v_reg;
  assign mem[3757] = mem_3757_sv2v_reg;
  assign mem[3756] = mem_3756_sv2v_reg;
  assign mem[3755] = mem_3755_sv2v_reg;
  assign mem[3754] = mem_3754_sv2v_reg;
  assign mem[3753] = mem_3753_sv2v_reg;
  assign mem[3752] = mem_3752_sv2v_reg;
  assign mem[3751] = mem_3751_sv2v_reg;
  assign mem[3750] = mem_3750_sv2v_reg;
  assign mem[3749] = mem_3749_sv2v_reg;
  assign mem[3748] = mem_3748_sv2v_reg;
  assign mem[3747] = mem_3747_sv2v_reg;
  assign mem[3746] = mem_3746_sv2v_reg;
  assign mem[3745] = mem_3745_sv2v_reg;
  assign mem[3744] = mem_3744_sv2v_reg;
  assign mem[3743] = mem_3743_sv2v_reg;
  assign mem[3742] = mem_3742_sv2v_reg;
  assign mem[3741] = mem_3741_sv2v_reg;
  assign mem[3740] = mem_3740_sv2v_reg;
  assign mem[3739] = mem_3739_sv2v_reg;
  assign mem[3738] = mem_3738_sv2v_reg;
  assign mem[3737] = mem_3737_sv2v_reg;
  assign mem[3736] = mem_3736_sv2v_reg;
  assign mem[3735] = mem_3735_sv2v_reg;
  assign mem[3734] = mem_3734_sv2v_reg;
  assign mem[3733] = mem_3733_sv2v_reg;
  assign mem[3732] = mem_3732_sv2v_reg;
  assign mem[3731] = mem_3731_sv2v_reg;
  assign mem[3730] = mem_3730_sv2v_reg;
  assign mem[3729] = mem_3729_sv2v_reg;
  assign mem[3728] = mem_3728_sv2v_reg;
  assign mem[3727] = mem_3727_sv2v_reg;
  assign mem[3726] = mem_3726_sv2v_reg;
  assign mem[3725] = mem_3725_sv2v_reg;
  assign mem[3724] = mem_3724_sv2v_reg;
  assign mem[3723] = mem_3723_sv2v_reg;
  assign mem[3722] = mem_3722_sv2v_reg;
  assign mem[3721] = mem_3721_sv2v_reg;
  assign mem[3720] = mem_3720_sv2v_reg;
  assign mem[3719] = mem_3719_sv2v_reg;
  assign mem[3718] = mem_3718_sv2v_reg;
  assign mem[3717] = mem_3717_sv2v_reg;
  assign mem[3716] = mem_3716_sv2v_reg;
  assign mem[3715] = mem_3715_sv2v_reg;
  assign mem[3714] = mem_3714_sv2v_reg;
  assign mem[3713] = mem_3713_sv2v_reg;
  assign mem[3712] = mem_3712_sv2v_reg;
  assign mem[3711] = mem_3711_sv2v_reg;
  assign mem[3710] = mem_3710_sv2v_reg;
  assign mem[3709] = mem_3709_sv2v_reg;
  assign mem[3708] = mem_3708_sv2v_reg;
  assign mem[3707] = mem_3707_sv2v_reg;
  assign mem[3706] = mem_3706_sv2v_reg;
  assign mem[3705] = mem_3705_sv2v_reg;
  assign mem[3704] = mem_3704_sv2v_reg;
  assign mem[3703] = mem_3703_sv2v_reg;
  assign mem[3702] = mem_3702_sv2v_reg;
  assign mem[3701] = mem_3701_sv2v_reg;
  assign mem[3700] = mem_3700_sv2v_reg;
  assign mem[3699] = mem_3699_sv2v_reg;
  assign mem[3698] = mem_3698_sv2v_reg;
  assign mem[3697] = mem_3697_sv2v_reg;
  assign mem[3696] = mem_3696_sv2v_reg;
  assign mem[3695] = mem_3695_sv2v_reg;
  assign mem[3694] = mem_3694_sv2v_reg;
  assign mem[3693] = mem_3693_sv2v_reg;
  assign mem[3692] = mem_3692_sv2v_reg;
  assign mem[3691] = mem_3691_sv2v_reg;
  assign mem[3690] = mem_3690_sv2v_reg;
  assign mem[3689] = mem_3689_sv2v_reg;
  assign mem[3688] = mem_3688_sv2v_reg;
  assign mem[3687] = mem_3687_sv2v_reg;
  assign mem[3686] = mem_3686_sv2v_reg;
  assign mem[3685] = mem_3685_sv2v_reg;
  assign mem[3684] = mem_3684_sv2v_reg;
  assign mem[3683] = mem_3683_sv2v_reg;
  assign mem[3682] = mem_3682_sv2v_reg;
  assign mem[3681] = mem_3681_sv2v_reg;
  assign mem[3680] = mem_3680_sv2v_reg;
  assign mem[3679] = mem_3679_sv2v_reg;
  assign mem[3678] = mem_3678_sv2v_reg;
  assign mem[3677] = mem_3677_sv2v_reg;
  assign mem[3676] = mem_3676_sv2v_reg;
  assign mem[3675] = mem_3675_sv2v_reg;
  assign mem[3674] = mem_3674_sv2v_reg;
  assign mem[3673] = mem_3673_sv2v_reg;
  assign mem[3672] = mem_3672_sv2v_reg;
  assign mem[3671] = mem_3671_sv2v_reg;
  assign mem[3670] = mem_3670_sv2v_reg;
  assign mem[3669] = mem_3669_sv2v_reg;
  assign mem[3668] = mem_3668_sv2v_reg;
  assign mem[3667] = mem_3667_sv2v_reg;
  assign mem[3666] = mem_3666_sv2v_reg;
  assign mem[3665] = mem_3665_sv2v_reg;
  assign mem[3664] = mem_3664_sv2v_reg;
  assign mem[3663] = mem_3663_sv2v_reg;
  assign mem[3662] = mem_3662_sv2v_reg;
  assign mem[3661] = mem_3661_sv2v_reg;
  assign mem[3660] = mem_3660_sv2v_reg;
  assign mem[3659] = mem_3659_sv2v_reg;
  assign mem[3658] = mem_3658_sv2v_reg;
  assign mem[3657] = mem_3657_sv2v_reg;
  assign mem[3656] = mem_3656_sv2v_reg;
  assign mem[3655] = mem_3655_sv2v_reg;
  assign mem[3654] = mem_3654_sv2v_reg;
  assign mem[3653] = mem_3653_sv2v_reg;
  assign mem[3652] = mem_3652_sv2v_reg;
  assign mem[3651] = mem_3651_sv2v_reg;
  assign mem[3650] = mem_3650_sv2v_reg;
  assign mem[3649] = mem_3649_sv2v_reg;
  assign mem[3648] = mem_3648_sv2v_reg;
  assign mem[3647] = mem_3647_sv2v_reg;
  assign mem[3646] = mem_3646_sv2v_reg;
  assign mem[3645] = mem_3645_sv2v_reg;
  assign mem[3644] = mem_3644_sv2v_reg;
  assign mem[3643] = mem_3643_sv2v_reg;
  assign mem[3642] = mem_3642_sv2v_reg;
  assign mem[3641] = mem_3641_sv2v_reg;
  assign mem[3640] = mem_3640_sv2v_reg;
  assign mem[3639] = mem_3639_sv2v_reg;
  assign mem[3638] = mem_3638_sv2v_reg;
  assign mem[3637] = mem_3637_sv2v_reg;
  assign mem[3636] = mem_3636_sv2v_reg;
  assign mem[3635] = mem_3635_sv2v_reg;
  assign mem[3634] = mem_3634_sv2v_reg;
  assign mem[3633] = mem_3633_sv2v_reg;
  assign mem[3632] = mem_3632_sv2v_reg;
  assign mem[3631] = mem_3631_sv2v_reg;
  assign mem[3630] = mem_3630_sv2v_reg;
  assign mem[3629] = mem_3629_sv2v_reg;
  assign mem[3628] = mem_3628_sv2v_reg;
  assign mem[3627] = mem_3627_sv2v_reg;
  assign mem[3626] = mem_3626_sv2v_reg;
  assign mem[3625] = mem_3625_sv2v_reg;
  assign mem[3624] = mem_3624_sv2v_reg;
  assign mem[3623] = mem_3623_sv2v_reg;
  assign mem[3622] = mem_3622_sv2v_reg;
  assign mem[3621] = mem_3621_sv2v_reg;
  assign mem[3620] = mem_3620_sv2v_reg;
  assign mem[3619] = mem_3619_sv2v_reg;
  assign mem[3618] = mem_3618_sv2v_reg;
  assign mem[3617] = mem_3617_sv2v_reg;
  assign mem[3616] = mem_3616_sv2v_reg;
  assign mem[3615] = mem_3615_sv2v_reg;
  assign mem[3614] = mem_3614_sv2v_reg;
  assign mem[3613] = mem_3613_sv2v_reg;
  assign mem[3612] = mem_3612_sv2v_reg;
  assign mem[3611] = mem_3611_sv2v_reg;
  assign mem[3610] = mem_3610_sv2v_reg;
  assign mem[3609] = mem_3609_sv2v_reg;
  assign mem[3608] = mem_3608_sv2v_reg;
  assign mem[3607] = mem_3607_sv2v_reg;
  assign mem[3606] = mem_3606_sv2v_reg;
  assign mem[3605] = mem_3605_sv2v_reg;
  assign mem[3604] = mem_3604_sv2v_reg;
  assign mem[3603] = mem_3603_sv2v_reg;
  assign mem[3602] = mem_3602_sv2v_reg;
  assign mem[3601] = mem_3601_sv2v_reg;
  assign mem[3600] = mem_3600_sv2v_reg;
  assign mem[3599] = mem_3599_sv2v_reg;
  assign mem[3598] = mem_3598_sv2v_reg;
  assign mem[3597] = mem_3597_sv2v_reg;
  assign mem[3596] = mem_3596_sv2v_reg;
  assign mem[3595] = mem_3595_sv2v_reg;
  assign mem[3594] = mem_3594_sv2v_reg;
  assign mem[3593] = mem_3593_sv2v_reg;
  assign mem[3592] = mem_3592_sv2v_reg;
  assign mem[3591] = mem_3591_sv2v_reg;
  assign mem[3590] = mem_3590_sv2v_reg;
  assign mem[3589] = mem_3589_sv2v_reg;
  assign mem[3588] = mem_3588_sv2v_reg;
  assign mem[3587] = mem_3587_sv2v_reg;
  assign mem[3586] = mem_3586_sv2v_reg;
  assign mem[3585] = mem_3585_sv2v_reg;
  assign mem[3584] = mem_3584_sv2v_reg;
  assign mem[3583] = mem_3583_sv2v_reg;
  assign mem[3582] = mem_3582_sv2v_reg;
  assign mem[3581] = mem_3581_sv2v_reg;
  assign mem[3580] = mem_3580_sv2v_reg;
  assign mem[3579] = mem_3579_sv2v_reg;
  assign mem[3578] = mem_3578_sv2v_reg;
  assign mem[3577] = mem_3577_sv2v_reg;
  assign mem[3576] = mem_3576_sv2v_reg;
  assign mem[3575] = mem_3575_sv2v_reg;
  assign mem[3574] = mem_3574_sv2v_reg;
  assign mem[3573] = mem_3573_sv2v_reg;
  assign mem[3572] = mem_3572_sv2v_reg;
  assign mem[3571] = mem_3571_sv2v_reg;
  assign mem[3570] = mem_3570_sv2v_reg;
  assign mem[3569] = mem_3569_sv2v_reg;
  assign mem[3568] = mem_3568_sv2v_reg;
  assign mem[3567] = mem_3567_sv2v_reg;
  assign mem[3566] = mem_3566_sv2v_reg;
  assign mem[3565] = mem_3565_sv2v_reg;
  assign mem[3564] = mem_3564_sv2v_reg;
  assign mem[3563] = mem_3563_sv2v_reg;
  assign mem[3562] = mem_3562_sv2v_reg;
  assign mem[3561] = mem_3561_sv2v_reg;
  assign mem[3560] = mem_3560_sv2v_reg;
  assign mem[3559] = mem_3559_sv2v_reg;
  assign mem[3558] = mem_3558_sv2v_reg;
  assign mem[3557] = mem_3557_sv2v_reg;
  assign mem[3556] = mem_3556_sv2v_reg;
  assign mem[3555] = mem_3555_sv2v_reg;
  assign mem[3554] = mem_3554_sv2v_reg;
  assign mem[3553] = mem_3553_sv2v_reg;
  assign mem[3552] = mem_3552_sv2v_reg;
  assign mem[3551] = mem_3551_sv2v_reg;
  assign mem[3550] = mem_3550_sv2v_reg;
  assign mem[3549] = mem_3549_sv2v_reg;
  assign mem[3548] = mem_3548_sv2v_reg;
  assign mem[3547] = mem_3547_sv2v_reg;
  assign mem[3546] = mem_3546_sv2v_reg;
  assign mem[3545] = mem_3545_sv2v_reg;
  assign mem[3544] = mem_3544_sv2v_reg;
  assign mem[3543] = mem_3543_sv2v_reg;
  assign mem[3542] = mem_3542_sv2v_reg;
  assign mem[3541] = mem_3541_sv2v_reg;
  assign mem[3540] = mem_3540_sv2v_reg;
  assign mem[3539] = mem_3539_sv2v_reg;
  assign mem[3538] = mem_3538_sv2v_reg;
  assign mem[3537] = mem_3537_sv2v_reg;
  assign mem[3536] = mem_3536_sv2v_reg;
  assign mem[3535] = mem_3535_sv2v_reg;
  assign mem[3534] = mem_3534_sv2v_reg;
  assign mem[3533] = mem_3533_sv2v_reg;
  assign mem[3532] = mem_3532_sv2v_reg;
  assign mem[3531] = mem_3531_sv2v_reg;
  assign mem[3530] = mem_3530_sv2v_reg;
  assign mem[3529] = mem_3529_sv2v_reg;
  assign mem[3528] = mem_3528_sv2v_reg;
  assign mem[3527] = mem_3527_sv2v_reg;
  assign mem[3526] = mem_3526_sv2v_reg;
  assign mem[3525] = mem_3525_sv2v_reg;
  assign mem[3524] = mem_3524_sv2v_reg;
  assign mem[3523] = mem_3523_sv2v_reg;
  assign mem[3522] = mem_3522_sv2v_reg;
  assign mem[3521] = mem_3521_sv2v_reg;
  assign mem[3520] = mem_3520_sv2v_reg;
  assign mem[3519] = mem_3519_sv2v_reg;
  assign mem[3518] = mem_3518_sv2v_reg;
  assign mem[3517] = mem_3517_sv2v_reg;
  assign mem[3516] = mem_3516_sv2v_reg;
  assign mem[3515] = mem_3515_sv2v_reg;
  assign mem[3514] = mem_3514_sv2v_reg;
  assign mem[3513] = mem_3513_sv2v_reg;
  assign mem[3512] = mem_3512_sv2v_reg;
  assign mem[3511] = mem_3511_sv2v_reg;
  assign mem[3510] = mem_3510_sv2v_reg;
  assign mem[3509] = mem_3509_sv2v_reg;
  assign mem[3508] = mem_3508_sv2v_reg;
  assign mem[3507] = mem_3507_sv2v_reg;
  assign mem[3506] = mem_3506_sv2v_reg;
  assign mem[3505] = mem_3505_sv2v_reg;
  assign mem[3504] = mem_3504_sv2v_reg;
  assign mem[3503] = mem_3503_sv2v_reg;
  assign mem[3502] = mem_3502_sv2v_reg;
  assign mem[3501] = mem_3501_sv2v_reg;
  assign mem[3500] = mem_3500_sv2v_reg;
  assign mem[3499] = mem_3499_sv2v_reg;
  assign mem[3498] = mem_3498_sv2v_reg;
  assign mem[3497] = mem_3497_sv2v_reg;
  assign mem[3496] = mem_3496_sv2v_reg;
  assign mem[3495] = mem_3495_sv2v_reg;
  assign mem[3494] = mem_3494_sv2v_reg;
  assign mem[3493] = mem_3493_sv2v_reg;
  assign mem[3492] = mem_3492_sv2v_reg;
  assign mem[3491] = mem_3491_sv2v_reg;
  assign mem[3490] = mem_3490_sv2v_reg;
  assign mem[3489] = mem_3489_sv2v_reg;
  assign mem[3488] = mem_3488_sv2v_reg;
  assign mem[3487] = mem_3487_sv2v_reg;
  assign mem[3486] = mem_3486_sv2v_reg;
  assign mem[3485] = mem_3485_sv2v_reg;
  assign mem[3484] = mem_3484_sv2v_reg;
  assign mem[3483] = mem_3483_sv2v_reg;
  assign mem[3482] = mem_3482_sv2v_reg;
  assign mem[3481] = mem_3481_sv2v_reg;
  assign mem[3480] = mem_3480_sv2v_reg;
  assign mem[3479] = mem_3479_sv2v_reg;
  assign mem[3478] = mem_3478_sv2v_reg;
  assign mem[3477] = mem_3477_sv2v_reg;
  assign mem[3476] = mem_3476_sv2v_reg;
  assign mem[3475] = mem_3475_sv2v_reg;
  assign mem[3474] = mem_3474_sv2v_reg;
  assign mem[3473] = mem_3473_sv2v_reg;
  assign mem[3472] = mem_3472_sv2v_reg;
  assign mem[3471] = mem_3471_sv2v_reg;
  assign mem[3470] = mem_3470_sv2v_reg;
  assign mem[3469] = mem_3469_sv2v_reg;
  assign mem[3468] = mem_3468_sv2v_reg;
  assign mem[3467] = mem_3467_sv2v_reg;
  assign mem[3466] = mem_3466_sv2v_reg;
  assign mem[3465] = mem_3465_sv2v_reg;
  assign mem[3464] = mem_3464_sv2v_reg;
  assign mem[3463] = mem_3463_sv2v_reg;
  assign mem[3462] = mem_3462_sv2v_reg;
  assign mem[3461] = mem_3461_sv2v_reg;
  assign mem[3460] = mem_3460_sv2v_reg;
  assign mem[3459] = mem_3459_sv2v_reg;
  assign mem[3458] = mem_3458_sv2v_reg;
  assign mem[3457] = mem_3457_sv2v_reg;
  assign mem[3456] = mem_3456_sv2v_reg;
  assign mem[3455] = mem_3455_sv2v_reg;
  assign mem[3454] = mem_3454_sv2v_reg;
  assign mem[3453] = mem_3453_sv2v_reg;
  assign mem[3452] = mem_3452_sv2v_reg;
  assign mem[3451] = mem_3451_sv2v_reg;
  assign mem[3450] = mem_3450_sv2v_reg;
  assign mem[3449] = mem_3449_sv2v_reg;
  assign mem[3448] = mem_3448_sv2v_reg;
  assign mem[3447] = mem_3447_sv2v_reg;
  assign mem[3446] = mem_3446_sv2v_reg;
  assign mem[3445] = mem_3445_sv2v_reg;
  assign mem[3444] = mem_3444_sv2v_reg;
  assign mem[3443] = mem_3443_sv2v_reg;
  assign mem[3442] = mem_3442_sv2v_reg;
  assign mem[3441] = mem_3441_sv2v_reg;
  assign mem[3440] = mem_3440_sv2v_reg;
  assign mem[3439] = mem_3439_sv2v_reg;
  assign mem[3438] = mem_3438_sv2v_reg;
  assign mem[3437] = mem_3437_sv2v_reg;
  assign mem[3436] = mem_3436_sv2v_reg;
  assign mem[3435] = mem_3435_sv2v_reg;
  assign mem[3434] = mem_3434_sv2v_reg;
  assign mem[3433] = mem_3433_sv2v_reg;
  assign mem[3432] = mem_3432_sv2v_reg;
  assign mem[3431] = mem_3431_sv2v_reg;
  assign mem[3430] = mem_3430_sv2v_reg;
  assign mem[3429] = mem_3429_sv2v_reg;
  assign mem[3428] = mem_3428_sv2v_reg;
  assign mem[3427] = mem_3427_sv2v_reg;
  assign mem[3426] = mem_3426_sv2v_reg;
  assign mem[3425] = mem_3425_sv2v_reg;
  assign mem[3424] = mem_3424_sv2v_reg;
  assign mem[3423] = mem_3423_sv2v_reg;
  assign mem[3422] = mem_3422_sv2v_reg;
  assign mem[3421] = mem_3421_sv2v_reg;
  assign mem[3420] = mem_3420_sv2v_reg;
  assign mem[3419] = mem_3419_sv2v_reg;
  assign mem[3418] = mem_3418_sv2v_reg;
  assign mem[3417] = mem_3417_sv2v_reg;
  assign mem[3416] = mem_3416_sv2v_reg;
  assign mem[3415] = mem_3415_sv2v_reg;
  assign mem[3414] = mem_3414_sv2v_reg;
  assign mem[3413] = mem_3413_sv2v_reg;
  assign mem[3412] = mem_3412_sv2v_reg;
  assign mem[3411] = mem_3411_sv2v_reg;
  assign mem[3410] = mem_3410_sv2v_reg;
  assign mem[3409] = mem_3409_sv2v_reg;
  assign mem[3408] = mem_3408_sv2v_reg;
  assign mem[3407] = mem_3407_sv2v_reg;
  assign mem[3406] = mem_3406_sv2v_reg;
  assign mem[3405] = mem_3405_sv2v_reg;
  assign mem[3404] = mem_3404_sv2v_reg;
  assign mem[3403] = mem_3403_sv2v_reg;
  assign mem[3402] = mem_3402_sv2v_reg;
  assign mem[3401] = mem_3401_sv2v_reg;
  assign mem[3400] = mem_3400_sv2v_reg;
  assign mem[3399] = mem_3399_sv2v_reg;
  assign mem[3398] = mem_3398_sv2v_reg;
  assign mem[3397] = mem_3397_sv2v_reg;
  assign mem[3396] = mem_3396_sv2v_reg;
  assign mem[3395] = mem_3395_sv2v_reg;
  assign mem[3394] = mem_3394_sv2v_reg;
  assign mem[3393] = mem_3393_sv2v_reg;
  assign mem[3392] = mem_3392_sv2v_reg;
  assign mem[3391] = mem_3391_sv2v_reg;
  assign mem[3390] = mem_3390_sv2v_reg;
  assign mem[3389] = mem_3389_sv2v_reg;
  assign mem[3388] = mem_3388_sv2v_reg;
  assign mem[3387] = mem_3387_sv2v_reg;
  assign mem[3386] = mem_3386_sv2v_reg;
  assign mem[3385] = mem_3385_sv2v_reg;
  assign mem[3384] = mem_3384_sv2v_reg;
  assign mem[3383] = mem_3383_sv2v_reg;
  assign mem[3382] = mem_3382_sv2v_reg;
  assign mem[3381] = mem_3381_sv2v_reg;
  assign mem[3380] = mem_3380_sv2v_reg;
  assign mem[3379] = mem_3379_sv2v_reg;
  assign mem[3378] = mem_3378_sv2v_reg;
  assign mem[3377] = mem_3377_sv2v_reg;
  assign mem[3376] = mem_3376_sv2v_reg;
  assign mem[3375] = mem_3375_sv2v_reg;
  assign mem[3374] = mem_3374_sv2v_reg;
  assign mem[3373] = mem_3373_sv2v_reg;
  assign mem[3372] = mem_3372_sv2v_reg;
  assign mem[3371] = mem_3371_sv2v_reg;
  assign mem[3370] = mem_3370_sv2v_reg;
  assign mem[3369] = mem_3369_sv2v_reg;
  assign mem[3368] = mem_3368_sv2v_reg;
  assign mem[3367] = mem_3367_sv2v_reg;
  assign mem[3366] = mem_3366_sv2v_reg;
  assign mem[3365] = mem_3365_sv2v_reg;
  assign mem[3364] = mem_3364_sv2v_reg;
  assign mem[3363] = mem_3363_sv2v_reg;
  assign mem[3362] = mem_3362_sv2v_reg;
  assign mem[3361] = mem_3361_sv2v_reg;
  assign mem[3360] = mem_3360_sv2v_reg;
  assign mem[3359] = mem_3359_sv2v_reg;
  assign mem[3358] = mem_3358_sv2v_reg;
  assign mem[3357] = mem_3357_sv2v_reg;
  assign mem[3356] = mem_3356_sv2v_reg;
  assign mem[3355] = mem_3355_sv2v_reg;
  assign mem[3354] = mem_3354_sv2v_reg;
  assign mem[3353] = mem_3353_sv2v_reg;
  assign mem[3352] = mem_3352_sv2v_reg;
  assign mem[3351] = mem_3351_sv2v_reg;
  assign mem[3350] = mem_3350_sv2v_reg;
  assign mem[3349] = mem_3349_sv2v_reg;
  assign mem[3348] = mem_3348_sv2v_reg;
  assign mem[3347] = mem_3347_sv2v_reg;
  assign mem[3346] = mem_3346_sv2v_reg;
  assign mem[3345] = mem_3345_sv2v_reg;
  assign mem[3344] = mem_3344_sv2v_reg;
  assign mem[3343] = mem_3343_sv2v_reg;
  assign mem[3342] = mem_3342_sv2v_reg;
  assign mem[3341] = mem_3341_sv2v_reg;
  assign mem[3340] = mem_3340_sv2v_reg;
  assign mem[3339] = mem_3339_sv2v_reg;
  assign mem[3338] = mem_3338_sv2v_reg;
  assign mem[3337] = mem_3337_sv2v_reg;
  assign mem[3336] = mem_3336_sv2v_reg;
  assign mem[3335] = mem_3335_sv2v_reg;
  assign mem[3334] = mem_3334_sv2v_reg;
  assign mem[3333] = mem_3333_sv2v_reg;
  assign mem[3332] = mem_3332_sv2v_reg;
  assign mem[3331] = mem_3331_sv2v_reg;
  assign mem[3330] = mem_3330_sv2v_reg;
  assign mem[3329] = mem_3329_sv2v_reg;
  assign mem[3328] = mem_3328_sv2v_reg;
  assign mem[3327] = mem_3327_sv2v_reg;
  assign mem[3326] = mem_3326_sv2v_reg;
  assign mem[3325] = mem_3325_sv2v_reg;
  assign mem[3324] = mem_3324_sv2v_reg;
  assign mem[3323] = mem_3323_sv2v_reg;
  assign mem[3322] = mem_3322_sv2v_reg;
  assign mem[3321] = mem_3321_sv2v_reg;
  assign mem[3320] = mem_3320_sv2v_reg;
  assign mem[3319] = mem_3319_sv2v_reg;
  assign mem[3318] = mem_3318_sv2v_reg;
  assign mem[3317] = mem_3317_sv2v_reg;
  assign mem[3316] = mem_3316_sv2v_reg;
  assign mem[3315] = mem_3315_sv2v_reg;
  assign mem[3314] = mem_3314_sv2v_reg;
  assign mem[3313] = mem_3313_sv2v_reg;
  assign mem[3312] = mem_3312_sv2v_reg;
  assign mem[3311] = mem_3311_sv2v_reg;
  assign mem[3310] = mem_3310_sv2v_reg;
  assign mem[3309] = mem_3309_sv2v_reg;
  assign mem[3308] = mem_3308_sv2v_reg;
  assign mem[3307] = mem_3307_sv2v_reg;
  assign mem[3306] = mem_3306_sv2v_reg;
  assign mem[3305] = mem_3305_sv2v_reg;
  assign mem[3304] = mem_3304_sv2v_reg;
  assign mem[3303] = mem_3303_sv2v_reg;
  assign mem[3302] = mem_3302_sv2v_reg;
  assign mem[3301] = mem_3301_sv2v_reg;
  assign mem[3300] = mem_3300_sv2v_reg;
  assign mem[3299] = mem_3299_sv2v_reg;
  assign mem[3298] = mem_3298_sv2v_reg;
  assign mem[3297] = mem_3297_sv2v_reg;
  assign mem[3296] = mem_3296_sv2v_reg;
  assign mem[3295] = mem_3295_sv2v_reg;
  assign mem[3294] = mem_3294_sv2v_reg;
  assign mem[3293] = mem_3293_sv2v_reg;
  assign mem[3292] = mem_3292_sv2v_reg;
  assign mem[3291] = mem_3291_sv2v_reg;
  assign mem[3290] = mem_3290_sv2v_reg;
  assign mem[3289] = mem_3289_sv2v_reg;
  assign mem[3288] = mem_3288_sv2v_reg;
  assign mem[3287] = mem_3287_sv2v_reg;
  assign mem[3286] = mem_3286_sv2v_reg;
  assign mem[3285] = mem_3285_sv2v_reg;
  assign mem[3284] = mem_3284_sv2v_reg;
  assign mem[3283] = mem_3283_sv2v_reg;
  assign mem[3282] = mem_3282_sv2v_reg;
  assign mem[3281] = mem_3281_sv2v_reg;
  assign mem[3280] = mem_3280_sv2v_reg;
  assign mem[3279] = mem_3279_sv2v_reg;
  assign mem[3278] = mem_3278_sv2v_reg;
  assign mem[3277] = mem_3277_sv2v_reg;
  assign mem[3276] = mem_3276_sv2v_reg;
  assign mem[3275] = mem_3275_sv2v_reg;
  assign mem[3274] = mem_3274_sv2v_reg;
  assign mem[3273] = mem_3273_sv2v_reg;
  assign mem[3272] = mem_3272_sv2v_reg;
  assign mem[3271] = mem_3271_sv2v_reg;
  assign mem[3270] = mem_3270_sv2v_reg;
  assign mem[3269] = mem_3269_sv2v_reg;
  assign mem[3268] = mem_3268_sv2v_reg;
  assign mem[3267] = mem_3267_sv2v_reg;
  assign mem[3266] = mem_3266_sv2v_reg;
  assign mem[3265] = mem_3265_sv2v_reg;
  assign mem[3264] = mem_3264_sv2v_reg;
  assign mem[3263] = mem_3263_sv2v_reg;
  assign mem[3262] = mem_3262_sv2v_reg;
  assign mem[3261] = mem_3261_sv2v_reg;
  assign mem[3260] = mem_3260_sv2v_reg;
  assign mem[3259] = mem_3259_sv2v_reg;
  assign mem[3258] = mem_3258_sv2v_reg;
  assign mem[3257] = mem_3257_sv2v_reg;
  assign mem[3256] = mem_3256_sv2v_reg;
  assign mem[3255] = mem_3255_sv2v_reg;
  assign mem[3254] = mem_3254_sv2v_reg;
  assign mem[3253] = mem_3253_sv2v_reg;
  assign mem[3252] = mem_3252_sv2v_reg;
  assign mem[3251] = mem_3251_sv2v_reg;
  assign mem[3250] = mem_3250_sv2v_reg;
  assign mem[3249] = mem_3249_sv2v_reg;
  assign mem[3248] = mem_3248_sv2v_reg;
  assign mem[3247] = mem_3247_sv2v_reg;
  assign mem[3246] = mem_3246_sv2v_reg;
  assign mem[3245] = mem_3245_sv2v_reg;
  assign mem[3244] = mem_3244_sv2v_reg;
  assign mem[3243] = mem_3243_sv2v_reg;
  assign mem[3242] = mem_3242_sv2v_reg;
  assign mem[3241] = mem_3241_sv2v_reg;
  assign mem[3240] = mem_3240_sv2v_reg;
  assign mem[3239] = mem_3239_sv2v_reg;
  assign mem[3238] = mem_3238_sv2v_reg;
  assign mem[3237] = mem_3237_sv2v_reg;
  assign mem[3236] = mem_3236_sv2v_reg;
  assign mem[3235] = mem_3235_sv2v_reg;
  assign mem[3234] = mem_3234_sv2v_reg;
  assign mem[3233] = mem_3233_sv2v_reg;
  assign mem[3232] = mem_3232_sv2v_reg;
  assign mem[3231] = mem_3231_sv2v_reg;
  assign mem[3230] = mem_3230_sv2v_reg;
  assign mem[3229] = mem_3229_sv2v_reg;
  assign mem[3228] = mem_3228_sv2v_reg;
  assign mem[3227] = mem_3227_sv2v_reg;
  assign mem[3226] = mem_3226_sv2v_reg;
  assign mem[3225] = mem_3225_sv2v_reg;
  assign mem[3224] = mem_3224_sv2v_reg;
  assign mem[3223] = mem_3223_sv2v_reg;
  assign mem[3222] = mem_3222_sv2v_reg;
  assign mem[3221] = mem_3221_sv2v_reg;
  assign mem[3220] = mem_3220_sv2v_reg;
  assign mem[3219] = mem_3219_sv2v_reg;
  assign mem[3218] = mem_3218_sv2v_reg;
  assign mem[3217] = mem_3217_sv2v_reg;
  assign mem[3216] = mem_3216_sv2v_reg;
  assign mem[3215] = mem_3215_sv2v_reg;
  assign mem[3214] = mem_3214_sv2v_reg;
  assign mem[3213] = mem_3213_sv2v_reg;
  assign mem[3212] = mem_3212_sv2v_reg;
  assign mem[3211] = mem_3211_sv2v_reg;
  assign mem[3210] = mem_3210_sv2v_reg;
  assign mem[3209] = mem_3209_sv2v_reg;
  assign mem[3208] = mem_3208_sv2v_reg;
  assign mem[3207] = mem_3207_sv2v_reg;
  assign mem[3206] = mem_3206_sv2v_reg;
  assign mem[3205] = mem_3205_sv2v_reg;
  assign mem[3204] = mem_3204_sv2v_reg;
  assign mem[3203] = mem_3203_sv2v_reg;
  assign mem[3202] = mem_3202_sv2v_reg;
  assign mem[3201] = mem_3201_sv2v_reg;
  assign mem[3200] = mem_3200_sv2v_reg;
  assign mem[3199] = mem_3199_sv2v_reg;
  assign mem[3198] = mem_3198_sv2v_reg;
  assign mem[3197] = mem_3197_sv2v_reg;
  assign mem[3196] = mem_3196_sv2v_reg;
  assign mem[3195] = mem_3195_sv2v_reg;
  assign mem[3194] = mem_3194_sv2v_reg;
  assign mem[3193] = mem_3193_sv2v_reg;
  assign mem[3192] = mem_3192_sv2v_reg;
  assign mem[3191] = mem_3191_sv2v_reg;
  assign mem[3190] = mem_3190_sv2v_reg;
  assign mem[3189] = mem_3189_sv2v_reg;
  assign mem[3188] = mem_3188_sv2v_reg;
  assign mem[3187] = mem_3187_sv2v_reg;
  assign mem[3186] = mem_3186_sv2v_reg;
  assign mem[3185] = mem_3185_sv2v_reg;
  assign mem[3184] = mem_3184_sv2v_reg;
  assign mem[3183] = mem_3183_sv2v_reg;
  assign mem[3182] = mem_3182_sv2v_reg;
  assign mem[3181] = mem_3181_sv2v_reg;
  assign mem[3180] = mem_3180_sv2v_reg;
  assign mem[3179] = mem_3179_sv2v_reg;
  assign mem[3178] = mem_3178_sv2v_reg;
  assign mem[3177] = mem_3177_sv2v_reg;
  assign mem[3176] = mem_3176_sv2v_reg;
  assign mem[3175] = mem_3175_sv2v_reg;
  assign mem[3174] = mem_3174_sv2v_reg;
  assign mem[3173] = mem_3173_sv2v_reg;
  assign mem[3172] = mem_3172_sv2v_reg;
  assign mem[3171] = mem_3171_sv2v_reg;
  assign mem[3170] = mem_3170_sv2v_reg;
  assign mem[3169] = mem_3169_sv2v_reg;
  assign mem[3168] = mem_3168_sv2v_reg;
  assign mem[3167] = mem_3167_sv2v_reg;
  assign mem[3166] = mem_3166_sv2v_reg;
  assign mem[3165] = mem_3165_sv2v_reg;
  assign mem[3164] = mem_3164_sv2v_reg;
  assign mem[3163] = mem_3163_sv2v_reg;
  assign mem[3162] = mem_3162_sv2v_reg;
  assign mem[3161] = mem_3161_sv2v_reg;
  assign mem[3160] = mem_3160_sv2v_reg;
  assign mem[3159] = mem_3159_sv2v_reg;
  assign mem[3158] = mem_3158_sv2v_reg;
  assign mem[3157] = mem_3157_sv2v_reg;
  assign mem[3156] = mem_3156_sv2v_reg;
  assign mem[3155] = mem_3155_sv2v_reg;
  assign mem[3154] = mem_3154_sv2v_reg;
  assign mem[3153] = mem_3153_sv2v_reg;
  assign mem[3152] = mem_3152_sv2v_reg;
  assign mem[3151] = mem_3151_sv2v_reg;
  assign mem[3150] = mem_3150_sv2v_reg;
  assign mem[3149] = mem_3149_sv2v_reg;
  assign mem[3148] = mem_3148_sv2v_reg;
  assign mem[3147] = mem_3147_sv2v_reg;
  assign mem[3146] = mem_3146_sv2v_reg;
  assign mem[3145] = mem_3145_sv2v_reg;
  assign mem[3144] = mem_3144_sv2v_reg;
  assign mem[3143] = mem_3143_sv2v_reg;
  assign mem[3142] = mem_3142_sv2v_reg;
  assign mem[3141] = mem_3141_sv2v_reg;
  assign mem[3140] = mem_3140_sv2v_reg;
  assign mem[3139] = mem_3139_sv2v_reg;
  assign mem[3138] = mem_3138_sv2v_reg;
  assign mem[3137] = mem_3137_sv2v_reg;
  assign mem[3136] = mem_3136_sv2v_reg;
  assign mem[3135] = mem_3135_sv2v_reg;
  assign mem[3134] = mem_3134_sv2v_reg;
  assign mem[3133] = mem_3133_sv2v_reg;
  assign mem[3132] = mem_3132_sv2v_reg;
  assign mem[3131] = mem_3131_sv2v_reg;
  assign mem[3130] = mem_3130_sv2v_reg;
  assign mem[3129] = mem_3129_sv2v_reg;
  assign mem[3128] = mem_3128_sv2v_reg;
  assign mem[3127] = mem_3127_sv2v_reg;
  assign mem[3126] = mem_3126_sv2v_reg;
  assign mem[3125] = mem_3125_sv2v_reg;
  assign mem[3124] = mem_3124_sv2v_reg;
  assign mem[3123] = mem_3123_sv2v_reg;
  assign mem[3122] = mem_3122_sv2v_reg;
  assign mem[3121] = mem_3121_sv2v_reg;
  assign mem[3120] = mem_3120_sv2v_reg;
  assign mem[3119] = mem_3119_sv2v_reg;
  assign mem[3118] = mem_3118_sv2v_reg;
  assign mem[3117] = mem_3117_sv2v_reg;
  assign mem[3116] = mem_3116_sv2v_reg;
  assign mem[3115] = mem_3115_sv2v_reg;
  assign mem[3114] = mem_3114_sv2v_reg;
  assign mem[3113] = mem_3113_sv2v_reg;
  assign mem[3112] = mem_3112_sv2v_reg;
  assign mem[3111] = mem_3111_sv2v_reg;
  assign mem[3110] = mem_3110_sv2v_reg;
  assign mem[3109] = mem_3109_sv2v_reg;
  assign mem[3108] = mem_3108_sv2v_reg;
  assign mem[3107] = mem_3107_sv2v_reg;
  assign mem[3106] = mem_3106_sv2v_reg;
  assign mem[3105] = mem_3105_sv2v_reg;
  assign mem[3104] = mem_3104_sv2v_reg;
  assign mem[3103] = mem_3103_sv2v_reg;
  assign mem[3102] = mem_3102_sv2v_reg;
  assign mem[3101] = mem_3101_sv2v_reg;
  assign mem[3100] = mem_3100_sv2v_reg;
  assign mem[3099] = mem_3099_sv2v_reg;
  assign mem[3098] = mem_3098_sv2v_reg;
  assign mem[3097] = mem_3097_sv2v_reg;
  assign mem[3096] = mem_3096_sv2v_reg;
  assign mem[3095] = mem_3095_sv2v_reg;
  assign mem[3094] = mem_3094_sv2v_reg;
  assign mem[3093] = mem_3093_sv2v_reg;
  assign mem[3092] = mem_3092_sv2v_reg;
  assign mem[3091] = mem_3091_sv2v_reg;
  assign mem[3090] = mem_3090_sv2v_reg;
  assign mem[3089] = mem_3089_sv2v_reg;
  assign mem[3088] = mem_3088_sv2v_reg;
  assign mem[3087] = mem_3087_sv2v_reg;
  assign mem[3086] = mem_3086_sv2v_reg;
  assign mem[3085] = mem_3085_sv2v_reg;
  assign mem[3084] = mem_3084_sv2v_reg;
  assign mem[3083] = mem_3083_sv2v_reg;
  assign mem[3082] = mem_3082_sv2v_reg;
  assign mem[3081] = mem_3081_sv2v_reg;
  assign mem[3080] = mem_3080_sv2v_reg;
  assign mem[3079] = mem_3079_sv2v_reg;
  assign mem[3078] = mem_3078_sv2v_reg;
  assign mem[3077] = mem_3077_sv2v_reg;
  assign mem[3076] = mem_3076_sv2v_reg;
  assign mem[3075] = mem_3075_sv2v_reg;
  assign mem[3074] = mem_3074_sv2v_reg;
  assign mem[3073] = mem_3073_sv2v_reg;
  assign mem[3072] = mem_3072_sv2v_reg;
  assign mem[3071] = mem_3071_sv2v_reg;
  assign mem[3070] = mem_3070_sv2v_reg;
  assign mem[3069] = mem_3069_sv2v_reg;
  assign mem[3068] = mem_3068_sv2v_reg;
  assign mem[3067] = mem_3067_sv2v_reg;
  assign mem[3066] = mem_3066_sv2v_reg;
  assign mem[3065] = mem_3065_sv2v_reg;
  assign mem[3064] = mem_3064_sv2v_reg;
  assign mem[3063] = mem_3063_sv2v_reg;
  assign mem[3062] = mem_3062_sv2v_reg;
  assign mem[3061] = mem_3061_sv2v_reg;
  assign mem[3060] = mem_3060_sv2v_reg;
  assign mem[3059] = mem_3059_sv2v_reg;
  assign mem[3058] = mem_3058_sv2v_reg;
  assign mem[3057] = mem_3057_sv2v_reg;
  assign mem[3056] = mem_3056_sv2v_reg;
  assign mem[3055] = mem_3055_sv2v_reg;
  assign mem[3054] = mem_3054_sv2v_reg;
  assign mem[3053] = mem_3053_sv2v_reg;
  assign mem[3052] = mem_3052_sv2v_reg;
  assign mem[3051] = mem_3051_sv2v_reg;
  assign mem[3050] = mem_3050_sv2v_reg;
  assign mem[3049] = mem_3049_sv2v_reg;
  assign mem[3048] = mem_3048_sv2v_reg;
  assign mem[3047] = mem_3047_sv2v_reg;
  assign mem[3046] = mem_3046_sv2v_reg;
  assign mem[3045] = mem_3045_sv2v_reg;
  assign mem[3044] = mem_3044_sv2v_reg;
  assign mem[3043] = mem_3043_sv2v_reg;
  assign mem[3042] = mem_3042_sv2v_reg;
  assign mem[3041] = mem_3041_sv2v_reg;
  assign mem[3040] = mem_3040_sv2v_reg;
  assign mem[3039] = mem_3039_sv2v_reg;
  assign mem[3038] = mem_3038_sv2v_reg;
  assign mem[3037] = mem_3037_sv2v_reg;
  assign mem[3036] = mem_3036_sv2v_reg;
  assign mem[3035] = mem_3035_sv2v_reg;
  assign mem[3034] = mem_3034_sv2v_reg;
  assign mem[3033] = mem_3033_sv2v_reg;
  assign mem[3032] = mem_3032_sv2v_reg;
  assign mem[3031] = mem_3031_sv2v_reg;
  assign mem[3030] = mem_3030_sv2v_reg;
  assign mem[3029] = mem_3029_sv2v_reg;
  assign mem[3028] = mem_3028_sv2v_reg;
  assign mem[3027] = mem_3027_sv2v_reg;
  assign mem[3026] = mem_3026_sv2v_reg;
  assign mem[3025] = mem_3025_sv2v_reg;
  assign mem[3024] = mem_3024_sv2v_reg;
  assign mem[3023] = mem_3023_sv2v_reg;
  assign mem[3022] = mem_3022_sv2v_reg;
  assign mem[3021] = mem_3021_sv2v_reg;
  assign mem[3020] = mem_3020_sv2v_reg;
  assign mem[3019] = mem_3019_sv2v_reg;
  assign mem[3018] = mem_3018_sv2v_reg;
  assign mem[3017] = mem_3017_sv2v_reg;
  assign mem[3016] = mem_3016_sv2v_reg;
  assign mem[3015] = mem_3015_sv2v_reg;
  assign mem[3014] = mem_3014_sv2v_reg;
  assign mem[3013] = mem_3013_sv2v_reg;
  assign mem[3012] = mem_3012_sv2v_reg;
  assign mem[3011] = mem_3011_sv2v_reg;
  assign mem[3010] = mem_3010_sv2v_reg;
  assign mem[3009] = mem_3009_sv2v_reg;
  assign mem[3008] = mem_3008_sv2v_reg;
  assign mem[3007] = mem_3007_sv2v_reg;
  assign mem[3006] = mem_3006_sv2v_reg;
  assign mem[3005] = mem_3005_sv2v_reg;
  assign mem[3004] = mem_3004_sv2v_reg;
  assign mem[3003] = mem_3003_sv2v_reg;
  assign mem[3002] = mem_3002_sv2v_reg;
  assign mem[3001] = mem_3001_sv2v_reg;
  assign mem[3000] = mem_3000_sv2v_reg;
  assign mem[2999] = mem_2999_sv2v_reg;
  assign mem[2998] = mem_2998_sv2v_reg;
  assign mem[2997] = mem_2997_sv2v_reg;
  assign mem[2996] = mem_2996_sv2v_reg;
  assign mem[2995] = mem_2995_sv2v_reg;
  assign mem[2994] = mem_2994_sv2v_reg;
  assign mem[2993] = mem_2993_sv2v_reg;
  assign mem[2992] = mem_2992_sv2v_reg;
  assign mem[2991] = mem_2991_sv2v_reg;
  assign mem[2990] = mem_2990_sv2v_reg;
  assign mem[2989] = mem_2989_sv2v_reg;
  assign mem[2988] = mem_2988_sv2v_reg;
  assign mem[2987] = mem_2987_sv2v_reg;
  assign mem[2986] = mem_2986_sv2v_reg;
  assign mem[2985] = mem_2985_sv2v_reg;
  assign mem[2984] = mem_2984_sv2v_reg;
  assign mem[2983] = mem_2983_sv2v_reg;
  assign mem[2982] = mem_2982_sv2v_reg;
  assign mem[2981] = mem_2981_sv2v_reg;
  assign mem[2980] = mem_2980_sv2v_reg;
  assign mem[2979] = mem_2979_sv2v_reg;
  assign mem[2978] = mem_2978_sv2v_reg;
  assign mem[2977] = mem_2977_sv2v_reg;
  assign mem[2976] = mem_2976_sv2v_reg;
  assign mem[2975] = mem_2975_sv2v_reg;
  assign mem[2974] = mem_2974_sv2v_reg;
  assign mem[2973] = mem_2973_sv2v_reg;
  assign mem[2972] = mem_2972_sv2v_reg;
  assign mem[2971] = mem_2971_sv2v_reg;
  assign mem[2970] = mem_2970_sv2v_reg;
  assign mem[2969] = mem_2969_sv2v_reg;
  assign mem[2968] = mem_2968_sv2v_reg;
  assign mem[2967] = mem_2967_sv2v_reg;
  assign mem[2966] = mem_2966_sv2v_reg;
  assign mem[2965] = mem_2965_sv2v_reg;
  assign mem[2964] = mem_2964_sv2v_reg;
  assign mem[2963] = mem_2963_sv2v_reg;
  assign mem[2962] = mem_2962_sv2v_reg;
  assign mem[2961] = mem_2961_sv2v_reg;
  assign mem[2960] = mem_2960_sv2v_reg;
  assign mem[2959] = mem_2959_sv2v_reg;
  assign mem[2958] = mem_2958_sv2v_reg;
  assign mem[2957] = mem_2957_sv2v_reg;
  assign mem[2956] = mem_2956_sv2v_reg;
  assign mem[2955] = mem_2955_sv2v_reg;
  assign mem[2954] = mem_2954_sv2v_reg;
  assign mem[2953] = mem_2953_sv2v_reg;
  assign mem[2952] = mem_2952_sv2v_reg;
  assign mem[2951] = mem_2951_sv2v_reg;
  assign mem[2950] = mem_2950_sv2v_reg;
  assign mem[2949] = mem_2949_sv2v_reg;
  assign mem[2948] = mem_2948_sv2v_reg;
  assign mem[2947] = mem_2947_sv2v_reg;
  assign mem[2946] = mem_2946_sv2v_reg;
  assign mem[2945] = mem_2945_sv2v_reg;
  assign mem[2944] = mem_2944_sv2v_reg;
  assign mem[2943] = mem_2943_sv2v_reg;
  assign mem[2942] = mem_2942_sv2v_reg;
  assign mem[2941] = mem_2941_sv2v_reg;
  assign mem[2940] = mem_2940_sv2v_reg;
  assign mem[2939] = mem_2939_sv2v_reg;
  assign mem[2938] = mem_2938_sv2v_reg;
  assign mem[2937] = mem_2937_sv2v_reg;
  assign mem[2936] = mem_2936_sv2v_reg;
  assign mem[2935] = mem_2935_sv2v_reg;
  assign mem[2934] = mem_2934_sv2v_reg;
  assign mem[2933] = mem_2933_sv2v_reg;
  assign mem[2932] = mem_2932_sv2v_reg;
  assign mem[2931] = mem_2931_sv2v_reg;
  assign mem[2930] = mem_2930_sv2v_reg;
  assign mem[2929] = mem_2929_sv2v_reg;
  assign mem[2928] = mem_2928_sv2v_reg;
  assign mem[2927] = mem_2927_sv2v_reg;
  assign mem[2926] = mem_2926_sv2v_reg;
  assign mem[2925] = mem_2925_sv2v_reg;
  assign mem[2924] = mem_2924_sv2v_reg;
  assign mem[2923] = mem_2923_sv2v_reg;
  assign mem[2922] = mem_2922_sv2v_reg;
  assign mem[2921] = mem_2921_sv2v_reg;
  assign mem[2920] = mem_2920_sv2v_reg;
  assign mem[2919] = mem_2919_sv2v_reg;
  assign mem[2918] = mem_2918_sv2v_reg;
  assign mem[2917] = mem_2917_sv2v_reg;
  assign mem[2916] = mem_2916_sv2v_reg;
  assign mem[2915] = mem_2915_sv2v_reg;
  assign mem[2914] = mem_2914_sv2v_reg;
  assign mem[2913] = mem_2913_sv2v_reg;
  assign mem[2912] = mem_2912_sv2v_reg;
  assign mem[2911] = mem_2911_sv2v_reg;
  assign mem[2910] = mem_2910_sv2v_reg;
  assign mem[2909] = mem_2909_sv2v_reg;
  assign mem[2908] = mem_2908_sv2v_reg;
  assign mem[2907] = mem_2907_sv2v_reg;
  assign mem[2906] = mem_2906_sv2v_reg;
  assign mem[2905] = mem_2905_sv2v_reg;
  assign mem[2904] = mem_2904_sv2v_reg;
  assign mem[2903] = mem_2903_sv2v_reg;
  assign mem[2902] = mem_2902_sv2v_reg;
  assign mem[2901] = mem_2901_sv2v_reg;
  assign mem[2900] = mem_2900_sv2v_reg;
  assign mem[2899] = mem_2899_sv2v_reg;
  assign mem[2898] = mem_2898_sv2v_reg;
  assign mem[2897] = mem_2897_sv2v_reg;
  assign mem[2896] = mem_2896_sv2v_reg;
  assign mem[2895] = mem_2895_sv2v_reg;
  assign mem[2894] = mem_2894_sv2v_reg;
  assign mem[2893] = mem_2893_sv2v_reg;
  assign mem[2892] = mem_2892_sv2v_reg;
  assign mem[2891] = mem_2891_sv2v_reg;
  assign mem[2890] = mem_2890_sv2v_reg;
  assign mem[2889] = mem_2889_sv2v_reg;
  assign mem[2888] = mem_2888_sv2v_reg;
  assign mem[2887] = mem_2887_sv2v_reg;
  assign mem[2886] = mem_2886_sv2v_reg;
  assign mem[2885] = mem_2885_sv2v_reg;
  assign mem[2884] = mem_2884_sv2v_reg;
  assign mem[2883] = mem_2883_sv2v_reg;
  assign mem[2882] = mem_2882_sv2v_reg;
  assign mem[2881] = mem_2881_sv2v_reg;
  assign mem[2880] = mem_2880_sv2v_reg;
  assign mem[2879] = mem_2879_sv2v_reg;
  assign mem[2878] = mem_2878_sv2v_reg;
  assign mem[2877] = mem_2877_sv2v_reg;
  assign mem[2876] = mem_2876_sv2v_reg;
  assign mem[2875] = mem_2875_sv2v_reg;
  assign mem[2874] = mem_2874_sv2v_reg;
  assign mem[2873] = mem_2873_sv2v_reg;
  assign mem[2872] = mem_2872_sv2v_reg;
  assign mem[2871] = mem_2871_sv2v_reg;
  assign mem[2870] = mem_2870_sv2v_reg;
  assign mem[2869] = mem_2869_sv2v_reg;
  assign mem[2868] = mem_2868_sv2v_reg;
  assign mem[2867] = mem_2867_sv2v_reg;
  assign mem[2866] = mem_2866_sv2v_reg;
  assign mem[2865] = mem_2865_sv2v_reg;
  assign mem[2864] = mem_2864_sv2v_reg;
  assign mem[2863] = mem_2863_sv2v_reg;
  assign mem[2862] = mem_2862_sv2v_reg;
  assign mem[2861] = mem_2861_sv2v_reg;
  assign mem[2860] = mem_2860_sv2v_reg;
  assign mem[2859] = mem_2859_sv2v_reg;
  assign mem[2858] = mem_2858_sv2v_reg;
  assign mem[2857] = mem_2857_sv2v_reg;
  assign mem[2856] = mem_2856_sv2v_reg;
  assign mem[2855] = mem_2855_sv2v_reg;
  assign mem[2854] = mem_2854_sv2v_reg;
  assign mem[2853] = mem_2853_sv2v_reg;
  assign mem[2852] = mem_2852_sv2v_reg;
  assign mem[2851] = mem_2851_sv2v_reg;
  assign mem[2850] = mem_2850_sv2v_reg;
  assign mem[2849] = mem_2849_sv2v_reg;
  assign mem[2848] = mem_2848_sv2v_reg;
  assign mem[2847] = mem_2847_sv2v_reg;
  assign mem[2846] = mem_2846_sv2v_reg;
  assign mem[2845] = mem_2845_sv2v_reg;
  assign mem[2844] = mem_2844_sv2v_reg;
  assign mem[2843] = mem_2843_sv2v_reg;
  assign mem[2842] = mem_2842_sv2v_reg;
  assign mem[2841] = mem_2841_sv2v_reg;
  assign mem[2840] = mem_2840_sv2v_reg;
  assign mem[2839] = mem_2839_sv2v_reg;
  assign mem[2838] = mem_2838_sv2v_reg;
  assign mem[2837] = mem_2837_sv2v_reg;
  assign mem[2836] = mem_2836_sv2v_reg;
  assign mem[2835] = mem_2835_sv2v_reg;
  assign mem[2834] = mem_2834_sv2v_reg;
  assign mem[2833] = mem_2833_sv2v_reg;
  assign mem[2832] = mem_2832_sv2v_reg;
  assign mem[2831] = mem_2831_sv2v_reg;
  assign mem[2830] = mem_2830_sv2v_reg;
  assign mem[2829] = mem_2829_sv2v_reg;
  assign mem[2828] = mem_2828_sv2v_reg;
  assign mem[2827] = mem_2827_sv2v_reg;
  assign mem[2826] = mem_2826_sv2v_reg;
  assign mem[2825] = mem_2825_sv2v_reg;
  assign mem[2824] = mem_2824_sv2v_reg;
  assign mem[2823] = mem_2823_sv2v_reg;
  assign mem[2822] = mem_2822_sv2v_reg;
  assign mem[2821] = mem_2821_sv2v_reg;
  assign mem[2820] = mem_2820_sv2v_reg;
  assign mem[2819] = mem_2819_sv2v_reg;
  assign mem[2818] = mem_2818_sv2v_reg;
  assign mem[2817] = mem_2817_sv2v_reg;
  assign mem[2816] = mem_2816_sv2v_reg;
  assign mem[2815] = mem_2815_sv2v_reg;
  assign mem[2814] = mem_2814_sv2v_reg;
  assign mem[2813] = mem_2813_sv2v_reg;
  assign mem[2812] = mem_2812_sv2v_reg;
  assign mem[2811] = mem_2811_sv2v_reg;
  assign mem[2810] = mem_2810_sv2v_reg;
  assign mem[2809] = mem_2809_sv2v_reg;
  assign mem[2808] = mem_2808_sv2v_reg;
  assign mem[2807] = mem_2807_sv2v_reg;
  assign mem[2806] = mem_2806_sv2v_reg;
  assign mem[2805] = mem_2805_sv2v_reg;
  assign mem[2804] = mem_2804_sv2v_reg;
  assign mem[2803] = mem_2803_sv2v_reg;
  assign mem[2802] = mem_2802_sv2v_reg;
  assign mem[2801] = mem_2801_sv2v_reg;
  assign mem[2800] = mem_2800_sv2v_reg;
  assign mem[2799] = mem_2799_sv2v_reg;
  assign mem[2798] = mem_2798_sv2v_reg;
  assign mem[2797] = mem_2797_sv2v_reg;
  assign mem[2796] = mem_2796_sv2v_reg;
  assign mem[2795] = mem_2795_sv2v_reg;
  assign mem[2794] = mem_2794_sv2v_reg;
  assign mem[2793] = mem_2793_sv2v_reg;
  assign mem[2792] = mem_2792_sv2v_reg;
  assign mem[2791] = mem_2791_sv2v_reg;
  assign mem[2790] = mem_2790_sv2v_reg;
  assign mem[2789] = mem_2789_sv2v_reg;
  assign mem[2788] = mem_2788_sv2v_reg;
  assign mem[2787] = mem_2787_sv2v_reg;
  assign mem[2786] = mem_2786_sv2v_reg;
  assign mem[2785] = mem_2785_sv2v_reg;
  assign mem[2784] = mem_2784_sv2v_reg;
  assign mem[2783] = mem_2783_sv2v_reg;
  assign mem[2782] = mem_2782_sv2v_reg;
  assign mem[2781] = mem_2781_sv2v_reg;
  assign mem[2780] = mem_2780_sv2v_reg;
  assign mem[2779] = mem_2779_sv2v_reg;
  assign mem[2778] = mem_2778_sv2v_reg;
  assign mem[2777] = mem_2777_sv2v_reg;
  assign mem[2776] = mem_2776_sv2v_reg;
  assign mem[2775] = mem_2775_sv2v_reg;
  assign mem[2774] = mem_2774_sv2v_reg;
  assign mem[2773] = mem_2773_sv2v_reg;
  assign mem[2772] = mem_2772_sv2v_reg;
  assign mem[2771] = mem_2771_sv2v_reg;
  assign mem[2770] = mem_2770_sv2v_reg;
  assign mem[2769] = mem_2769_sv2v_reg;
  assign mem[2768] = mem_2768_sv2v_reg;
  assign mem[2767] = mem_2767_sv2v_reg;
  assign mem[2766] = mem_2766_sv2v_reg;
  assign mem[2765] = mem_2765_sv2v_reg;
  assign mem[2764] = mem_2764_sv2v_reg;
  assign mem[2763] = mem_2763_sv2v_reg;
  assign mem[2762] = mem_2762_sv2v_reg;
  assign mem[2761] = mem_2761_sv2v_reg;
  assign mem[2760] = mem_2760_sv2v_reg;
  assign mem[2759] = mem_2759_sv2v_reg;
  assign mem[2758] = mem_2758_sv2v_reg;
  assign mem[2757] = mem_2757_sv2v_reg;
  assign mem[2756] = mem_2756_sv2v_reg;
  assign mem[2755] = mem_2755_sv2v_reg;
  assign mem[2754] = mem_2754_sv2v_reg;
  assign mem[2753] = mem_2753_sv2v_reg;
  assign mem[2752] = mem_2752_sv2v_reg;
  assign mem[2751] = mem_2751_sv2v_reg;
  assign mem[2750] = mem_2750_sv2v_reg;
  assign mem[2749] = mem_2749_sv2v_reg;
  assign mem[2748] = mem_2748_sv2v_reg;
  assign mem[2747] = mem_2747_sv2v_reg;
  assign mem[2746] = mem_2746_sv2v_reg;
  assign mem[2745] = mem_2745_sv2v_reg;
  assign mem[2744] = mem_2744_sv2v_reg;
  assign mem[2743] = mem_2743_sv2v_reg;
  assign mem[2742] = mem_2742_sv2v_reg;
  assign mem[2741] = mem_2741_sv2v_reg;
  assign mem[2740] = mem_2740_sv2v_reg;
  assign mem[2739] = mem_2739_sv2v_reg;
  assign mem[2738] = mem_2738_sv2v_reg;
  assign mem[2737] = mem_2737_sv2v_reg;
  assign mem[2736] = mem_2736_sv2v_reg;
  assign mem[2735] = mem_2735_sv2v_reg;
  assign mem[2734] = mem_2734_sv2v_reg;
  assign mem[2733] = mem_2733_sv2v_reg;
  assign mem[2732] = mem_2732_sv2v_reg;
  assign mem[2731] = mem_2731_sv2v_reg;
  assign mem[2730] = mem_2730_sv2v_reg;
  assign mem[2729] = mem_2729_sv2v_reg;
  assign mem[2728] = mem_2728_sv2v_reg;
  assign mem[2727] = mem_2727_sv2v_reg;
  assign mem[2726] = mem_2726_sv2v_reg;
  assign mem[2725] = mem_2725_sv2v_reg;
  assign mem[2724] = mem_2724_sv2v_reg;
  assign mem[2723] = mem_2723_sv2v_reg;
  assign mem[2722] = mem_2722_sv2v_reg;
  assign mem[2721] = mem_2721_sv2v_reg;
  assign mem[2720] = mem_2720_sv2v_reg;
  assign mem[2719] = mem_2719_sv2v_reg;
  assign mem[2718] = mem_2718_sv2v_reg;
  assign mem[2717] = mem_2717_sv2v_reg;
  assign mem[2716] = mem_2716_sv2v_reg;
  assign mem[2715] = mem_2715_sv2v_reg;
  assign mem[2714] = mem_2714_sv2v_reg;
  assign mem[2713] = mem_2713_sv2v_reg;
  assign mem[2712] = mem_2712_sv2v_reg;
  assign mem[2711] = mem_2711_sv2v_reg;
  assign mem[2710] = mem_2710_sv2v_reg;
  assign mem[2709] = mem_2709_sv2v_reg;
  assign mem[2708] = mem_2708_sv2v_reg;
  assign mem[2707] = mem_2707_sv2v_reg;
  assign mem[2706] = mem_2706_sv2v_reg;
  assign mem[2705] = mem_2705_sv2v_reg;
  assign mem[2704] = mem_2704_sv2v_reg;
  assign mem[2703] = mem_2703_sv2v_reg;
  assign mem[2702] = mem_2702_sv2v_reg;
  assign mem[2701] = mem_2701_sv2v_reg;
  assign mem[2700] = mem_2700_sv2v_reg;
  assign mem[2699] = mem_2699_sv2v_reg;
  assign mem[2698] = mem_2698_sv2v_reg;
  assign mem[2697] = mem_2697_sv2v_reg;
  assign mem[2696] = mem_2696_sv2v_reg;
  assign mem[2695] = mem_2695_sv2v_reg;
  assign mem[2694] = mem_2694_sv2v_reg;
  assign mem[2693] = mem_2693_sv2v_reg;
  assign mem[2692] = mem_2692_sv2v_reg;
  assign mem[2691] = mem_2691_sv2v_reg;
  assign mem[2690] = mem_2690_sv2v_reg;
  assign mem[2689] = mem_2689_sv2v_reg;
  assign mem[2688] = mem_2688_sv2v_reg;
  assign mem[2687] = mem_2687_sv2v_reg;
  assign mem[2686] = mem_2686_sv2v_reg;
  assign mem[2685] = mem_2685_sv2v_reg;
  assign mem[2684] = mem_2684_sv2v_reg;
  assign mem[2683] = mem_2683_sv2v_reg;
  assign mem[2682] = mem_2682_sv2v_reg;
  assign mem[2681] = mem_2681_sv2v_reg;
  assign mem[2680] = mem_2680_sv2v_reg;
  assign mem[2679] = mem_2679_sv2v_reg;
  assign mem[2678] = mem_2678_sv2v_reg;
  assign mem[2677] = mem_2677_sv2v_reg;
  assign mem[2676] = mem_2676_sv2v_reg;
  assign mem[2675] = mem_2675_sv2v_reg;
  assign mem[2674] = mem_2674_sv2v_reg;
  assign mem[2673] = mem_2673_sv2v_reg;
  assign mem[2672] = mem_2672_sv2v_reg;
  assign mem[2671] = mem_2671_sv2v_reg;
  assign mem[2670] = mem_2670_sv2v_reg;
  assign mem[2669] = mem_2669_sv2v_reg;
  assign mem[2668] = mem_2668_sv2v_reg;
  assign mem[2667] = mem_2667_sv2v_reg;
  assign mem[2666] = mem_2666_sv2v_reg;
  assign mem[2665] = mem_2665_sv2v_reg;
  assign mem[2664] = mem_2664_sv2v_reg;
  assign mem[2663] = mem_2663_sv2v_reg;
  assign mem[2662] = mem_2662_sv2v_reg;
  assign mem[2661] = mem_2661_sv2v_reg;
  assign mem[2660] = mem_2660_sv2v_reg;
  assign mem[2659] = mem_2659_sv2v_reg;
  assign mem[2658] = mem_2658_sv2v_reg;
  assign mem[2657] = mem_2657_sv2v_reg;
  assign mem[2656] = mem_2656_sv2v_reg;
  assign mem[2655] = mem_2655_sv2v_reg;
  assign mem[2654] = mem_2654_sv2v_reg;
  assign mem[2653] = mem_2653_sv2v_reg;
  assign mem[2652] = mem_2652_sv2v_reg;
  assign mem[2651] = mem_2651_sv2v_reg;
  assign mem[2650] = mem_2650_sv2v_reg;
  assign mem[2649] = mem_2649_sv2v_reg;
  assign mem[2648] = mem_2648_sv2v_reg;
  assign mem[2647] = mem_2647_sv2v_reg;
  assign mem[2646] = mem_2646_sv2v_reg;
  assign mem[2645] = mem_2645_sv2v_reg;
  assign mem[2644] = mem_2644_sv2v_reg;
  assign mem[2643] = mem_2643_sv2v_reg;
  assign mem[2642] = mem_2642_sv2v_reg;
  assign mem[2641] = mem_2641_sv2v_reg;
  assign mem[2640] = mem_2640_sv2v_reg;
  assign mem[2639] = mem_2639_sv2v_reg;
  assign mem[2638] = mem_2638_sv2v_reg;
  assign mem[2637] = mem_2637_sv2v_reg;
  assign mem[2636] = mem_2636_sv2v_reg;
  assign mem[2635] = mem_2635_sv2v_reg;
  assign mem[2634] = mem_2634_sv2v_reg;
  assign mem[2633] = mem_2633_sv2v_reg;
  assign mem[2632] = mem_2632_sv2v_reg;
  assign mem[2631] = mem_2631_sv2v_reg;
  assign mem[2630] = mem_2630_sv2v_reg;
  assign mem[2629] = mem_2629_sv2v_reg;
  assign mem[2628] = mem_2628_sv2v_reg;
  assign mem[2627] = mem_2627_sv2v_reg;
  assign mem[2626] = mem_2626_sv2v_reg;
  assign mem[2625] = mem_2625_sv2v_reg;
  assign mem[2624] = mem_2624_sv2v_reg;
  assign mem[2623] = mem_2623_sv2v_reg;
  assign mem[2622] = mem_2622_sv2v_reg;
  assign mem[2621] = mem_2621_sv2v_reg;
  assign mem[2620] = mem_2620_sv2v_reg;
  assign mem[2619] = mem_2619_sv2v_reg;
  assign mem[2618] = mem_2618_sv2v_reg;
  assign mem[2617] = mem_2617_sv2v_reg;
  assign mem[2616] = mem_2616_sv2v_reg;
  assign mem[2615] = mem_2615_sv2v_reg;
  assign mem[2614] = mem_2614_sv2v_reg;
  assign mem[2613] = mem_2613_sv2v_reg;
  assign mem[2612] = mem_2612_sv2v_reg;
  assign mem[2611] = mem_2611_sv2v_reg;
  assign mem[2610] = mem_2610_sv2v_reg;
  assign mem[2609] = mem_2609_sv2v_reg;
  assign mem[2608] = mem_2608_sv2v_reg;
  assign mem[2607] = mem_2607_sv2v_reg;
  assign mem[2606] = mem_2606_sv2v_reg;
  assign mem[2605] = mem_2605_sv2v_reg;
  assign mem[2604] = mem_2604_sv2v_reg;
  assign mem[2603] = mem_2603_sv2v_reg;
  assign mem[2602] = mem_2602_sv2v_reg;
  assign mem[2601] = mem_2601_sv2v_reg;
  assign mem[2600] = mem_2600_sv2v_reg;
  assign mem[2599] = mem_2599_sv2v_reg;
  assign mem[2598] = mem_2598_sv2v_reg;
  assign mem[2597] = mem_2597_sv2v_reg;
  assign mem[2596] = mem_2596_sv2v_reg;
  assign mem[2595] = mem_2595_sv2v_reg;
  assign mem[2594] = mem_2594_sv2v_reg;
  assign mem[2593] = mem_2593_sv2v_reg;
  assign mem[2592] = mem_2592_sv2v_reg;
  assign mem[2591] = mem_2591_sv2v_reg;
  assign mem[2590] = mem_2590_sv2v_reg;
  assign mem[2589] = mem_2589_sv2v_reg;
  assign mem[2588] = mem_2588_sv2v_reg;
  assign mem[2587] = mem_2587_sv2v_reg;
  assign mem[2586] = mem_2586_sv2v_reg;
  assign mem[2585] = mem_2585_sv2v_reg;
  assign mem[2584] = mem_2584_sv2v_reg;
  assign mem[2583] = mem_2583_sv2v_reg;
  assign mem[2582] = mem_2582_sv2v_reg;
  assign mem[2581] = mem_2581_sv2v_reg;
  assign mem[2580] = mem_2580_sv2v_reg;
  assign mem[2579] = mem_2579_sv2v_reg;
  assign mem[2578] = mem_2578_sv2v_reg;
  assign mem[2577] = mem_2577_sv2v_reg;
  assign mem[2576] = mem_2576_sv2v_reg;
  assign mem[2575] = mem_2575_sv2v_reg;
  assign mem[2574] = mem_2574_sv2v_reg;
  assign mem[2573] = mem_2573_sv2v_reg;
  assign mem[2572] = mem_2572_sv2v_reg;
  assign mem[2571] = mem_2571_sv2v_reg;
  assign mem[2570] = mem_2570_sv2v_reg;
  assign mem[2569] = mem_2569_sv2v_reg;
  assign mem[2568] = mem_2568_sv2v_reg;
  assign mem[2567] = mem_2567_sv2v_reg;
  assign mem[2566] = mem_2566_sv2v_reg;
  assign mem[2565] = mem_2565_sv2v_reg;
  assign mem[2564] = mem_2564_sv2v_reg;
  assign mem[2563] = mem_2563_sv2v_reg;
  assign mem[2562] = mem_2562_sv2v_reg;
  assign mem[2561] = mem_2561_sv2v_reg;
  assign mem[2560] = mem_2560_sv2v_reg;
  assign mem[2559] = mem_2559_sv2v_reg;
  assign mem[2558] = mem_2558_sv2v_reg;
  assign mem[2557] = mem_2557_sv2v_reg;
  assign mem[2556] = mem_2556_sv2v_reg;
  assign mem[2555] = mem_2555_sv2v_reg;
  assign mem[2554] = mem_2554_sv2v_reg;
  assign mem[2553] = mem_2553_sv2v_reg;
  assign mem[2552] = mem_2552_sv2v_reg;
  assign mem[2551] = mem_2551_sv2v_reg;
  assign mem[2550] = mem_2550_sv2v_reg;
  assign mem[2549] = mem_2549_sv2v_reg;
  assign mem[2548] = mem_2548_sv2v_reg;
  assign mem[2547] = mem_2547_sv2v_reg;
  assign mem[2546] = mem_2546_sv2v_reg;
  assign mem[2545] = mem_2545_sv2v_reg;
  assign mem[2544] = mem_2544_sv2v_reg;
  assign mem[2543] = mem_2543_sv2v_reg;
  assign mem[2542] = mem_2542_sv2v_reg;
  assign mem[2541] = mem_2541_sv2v_reg;
  assign mem[2540] = mem_2540_sv2v_reg;
  assign mem[2539] = mem_2539_sv2v_reg;
  assign mem[2538] = mem_2538_sv2v_reg;
  assign mem[2537] = mem_2537_sv2v_reg;
  assign mem[2536] = mem_2536_sv2v_reg;
  assign mem[2535] = mem_2535_sv2v_reg;
  assign mem[2534] = mem_2534_sv2v_reg;
  assign mem[2533] = mem_2533_sv2v_reg;
  assign mem[2532] = mem_2532_sv2v_reg;
  assign mem[2531] = mem_2531_sv2v_reg;
  assign mem[2530] = mem_2530_sv2v_reg;
  assign mem[2529] = mem_2529_sv2v_reg;
  assign mem[2528] = mem_2528_sv2v_reg;
  assign mem[2527] = mem_2527_sv2v_reg;
  assign mem[2526] = mem_2526_sv2v_reg;
  assign mem[2525] = mem_2525_sv2v_reg;
  assign mem[2524] = mem_2524_sv2v_reg;
  assign mem[2523] = mem_2523_sv2v_reg;
  assign mem[2522] = mem_2522_sv2v_reg;
  assign mem[2521] = mem_2521_sv2v_reg;
  assign mem[2520] = mem_2520_sv2v_reg;
  assign mem[2519] = mem_2519_sv2v_reg;
  assign mem[2518] = mem_2518_sv2v_reg;
  assign mem[2517] = mem_2517_sv2v_reg;
  assign mem[2516] = mem_2516_sv2v_reg;
  assign mem[2515] = mem_2515_sv2v_reg;
  assign mem[2514] = mem_2514_sv2v_reg;
  assign mem[2513] = mem_2513_sv2v_reg;
  assign mem[2512] = mem_2512_sv2v_reg;
  assign mem[2511] = mem_2511_sv2v_reg;
  assign mem[2510] = mem_2510_sv2v_reg;
  assign mem[2509] = mem_2509_sv2v_reg;
  assign mem[2508] = mem_2508_sv2v_reg;
  assign mem[2507] = mem_2507_sv2v_reg;
  assign mem[2506] = mem_2506_sv2v_reg;
  assign mem[2505] = mem_2505_sv2v_reg;
  assign mem[2504] = mem_2504_sv2v_reg;
  assign mem[2503] = mem_2503_sv2v_reg;
  assign mem[2502] = mem_2502_sv2v_reg;
  assign mem[2501] = mem_2501_sv2v_reg;
  assign mem[2500] = mem_2500_sv2v_reg;
  assign mem[2499] = mem_2499_sv2v_reg;
  assign mem[2498] = mem_2498_sv2v_reg;
  assign mem[2497] = mem_2497_sv2v_reg;
  assign mem[2496] = mem_2496_sv2v_reg;
  assign mem[2495] = mem_2495_sv2v_reg;
  assign mem[2494] = mem_2494_sv2v_reg;
  assign mem[2493] = mem_2493_sv2v_reg;
  assign mem[2492] = mem_2492_sv2v_reg;
  assign mem[2491] = mem_2491_sv2v_reg;
  assign mem[2490] = mem_2490_sv2v_reg;
  assign mem[2489] = mem_2489_sv2v_reg;
  assign mem[2488] = mem_2488_sv2v_reg;
  assign mem[2487] = mem_2487_sv2v_reg;
  assign mem[2486] = mem_2486_sv2v_reg;
  assign mem[2485] = mem_2485_sv2v_reg;
  assign mem[2484] = mem_2484_sv2v_reg;
  assign mem[2483] = mem_2483_sv2v_reg;
  assign mem[2482] = mem_2482_sv2v_reg;
  assign mem[2481] = mem_2481_sv2v_reg;
  assign mem[2480] = mem_2480_sv2v_reg;
  assign mem[2479] = mem_2479_sv2v_reg;
  assign mem[2478] = mem_2478_sv2v_reg;
  assign mem[2477] = mem_2477_sv2v_reg;
  assign mem[2476] = mem_2476_sv2v_reg;
  assign mem[2475] = mem_2475_sv2v_reg;
  assign mem[2474] = mem_2474_sv2v_reg;
  assign mem[2473] = mem_2473_sv2v_reg;
  assign mem[2472] = mem_2472_sv2v_reg;
  assign mem[2471] = mem_2471_sv2v_reg;
  assign mem[2470] = mem_2470_sv2v_reg;
  assign mem[2469] = mem_2469_sv2v_reg;
  assign mem[2468] = mem_2468_sv2v_reg;
  assign mem[2467] = mem_2467_sv2v_reg;
  assign mem[2466] = mem_2466_sv2v_reg;
  assign mem[2465] = mem_2465_sv2v_reg;
  assign mem[2464] = mem_2464_sv2v_reg;
  assign mem[2463] = mem_2463_sv2v_reg;
  assign mem[2462] = mem_2462_sv2v_reg;
  assign mem[2461] = mem_2461_sv2v_reg;
  assign mem[2460] = mem_2460_sv2v_reg;
  assign mem[2459] = mem_2459_sv2v_reg;
  assign mem[2458] = mem_2458_sv2v_reg;
  assign mem[2457] = mem_2457_sv2v_reg;
  assign mem[2456] = mem_2456_sv2v_reg;
  assign mem[2455] = mem_2455_sv2v_reg;
  assign mem[2454] = mem_2454_sv2v_reg;
  assign mem[2453] = mem_2453_sv2v_reg;
  assign mem[2452] = mem_2452_sv2v_reg;
  assign mem[2451] = mem_2451_sv2v_reg;
  assign mem[2450] = mem_2450_sv2v_reg;
  assign mem[2449] = mem_2449_sv2v_reg;
  assign mem[2448] = mem_2448_sv2v_reg;
  assign mem[2447] = mem_2447_sv2v_reg;
  assign mem[2446] = mem_2446_sv2v_reg;
  assign mem[2445] = mem_2445_sv2v_reg;
  assign mem[2444] = mem_2444_sv2v_reg;
  assign mem[2443] = mem_2443_sv2v_reg;
  assign mem[2442] = mem_2442_sv2v_reg;
  assign mem[2441] = mem_2441_sv2v_reg;
  assign mem[2440] = mem_2440_sv2v_reg;
  assign mem[2439] = mem_2439_sv2v_reg;
  assign mem[2438] = mem_2438_sv2v_reg;
  assign mem[2437] = mem_2437_sv2v_reg;
  assign mem[2436] = mem_2436_sv2v_reg;
  assign mem[2435] = mem_2435_sv2v_reg;
  assign mem[2434] = mem_2434_sv2v_reg;
  assign mem[2433] = mem_2433_sv2v_reg;
  assign mem[2432] = mem_2432_sv2v_reg;
  assign mem[2431] = mem_2431_sv2v_reg;
  assign mem[2430] = mem_2430_sv2v_reg;
  assign mem[2429] = mem_2429_sv2v_reg;
  assign mem[2428] = mem_2428_sv2v_reg;
  assign mem[2427] = mem_2427_sv2v_reg;
  assign mem[2426] = mem_2426_sv2v_reg;
  assign mem[2425] = mem_2425_sv2v_reg;
  assign mem[2424] = mem_2424_sv2v_reg;
  assign mem[2423] = mem_2423_sv2v_reg;
  assign mem[2422] = mem_2422_sv2v_reg;
  assign mem[2421] = mem_2421_sv2v_reg;
  assign mem[2420] = mem_2420_sv2v_reg;
  assign mem[2419] = mem_2419_sv2v_reg;
  assign mem[2418] = mem_2418_sv2v_reg;
  assign mem[2417] = mem_2417_sv2v_reg;
  assign mem[2416] = mem_2416_sv2v_reg;
  assign mem[2415] = mem_2415_sv2v_reg;
  assign mem[2414] = mem_2414_sv2v_reg;
  assign mem[2413] = mem_2413_sv2v_reg;
  assign mem[2412] = mem_2412_sv2v_reg;
  assign mem[2411] = mem_2411_sv2v_reg;
  assign mem[2410] = mem_2410_sv2v_reg;
  assign mem[2409] = mem_2409_sv2v_reg;
  assign mem[2408] = mem_2408_sv2v_reg;
  assign mem[2407] = mem_2407_sv2v_reg;
  assign mem[2406] = mem_2406_sv2v_reg;
  assign mem[2405] = mem_2405_sv2v_reg;
  assign mem[2404] = mem_2404_sv2v_reg;
  assign mem[2403] = mem_2403_sv2v_reg;
  assign mem[2402] = mem_2402_sv2v_reg;
  assign mem[2401] = mem_2401_sv2v_reg;
  assign mem[2400] = mem_2400_sv2v_reg;
  assign mem[2399] = mem_2399_sv2v_reg;
  assign mem[2398] = mem_2398_sv2v_reg;
  assign mem[2397] = mem_2397_sv2v_reg;
  assign mem[2396] = mem_2396_sv2v_reg;
  assign mem[2395] = mem_2395_sv2v_reg;
  assign mem[2394] = mem_2394_sv2v_reg;
  assign mem[2393] = mem_2393_sv2v_reg;
  assign mem[2392] = mem_2392_sv2v_reg;
  assign mem[2391] = mem_2391_sv2v_reg;
  assign mem[2390] = mem_2390_sv2v_reg;
  assign mem[2389] = mem_2389_sv2v_reg;
  assign mem[2388] = mem_2388_sv2v_reg;
  assign mem[2387] = mem_2387_sv2v_reg;
  assign mem[2386] = mem_2386_sv2v_reg;
  assign mem[2385] = mem_2385_sv2v_reg;
  assign mem[2384] = mem_2384_sv2v_reg;
  assign mem[2383] = mem_2383_sv2v_reg;
  assign mem[2382] = mem_2382_sv2v_reg;
  assign mem[2381] = mem_2381_sv2v_reg;
  assign mem[2380] = mem_2380_sv2v_reg;
  assign mem[2379] = mem_2379_sv2v_reg;
  assign mem[2378] = mem_2378_sv2v_reg;
  assign mem[2377] = mem_2377_sv2v_reg;
  assign mem[2376] = mem_2376_sv2v_reg;
  assign mem[2375] = mem_2375_sv2v_reg;
  assign mem[2374] = mem_2374_sv2v_reg;
  assign mem[2373] = mem_2373_sv2v_reg;
  assign mem[2372] = mem_2372_sv2v_reg;
  assign mem[2371] = mem_2371_sv2v_reg;
  assign mem[2370] = mem_2370_sv2v_reg;
  assign mem[2369] = mem_2369_sv2v_reg;
  assign mem[2368] = mem_2368_sv2v_reg;
  assign mem[2367] = mem_2367_sv2v_reg;
  assign mem[2366] = mem_2366_sv2v_reg;
  assign mem[2365] = mem_2365_sv2v_reg;
  assign mem[2364] = mem_2364_sv2v_reg;
  assign mem[2363] = mem_2363_sv2v_reg;
  assign mem[2362] = mem_2362_sv2v_reg;
  assign mem[2361] = mem_2361_sv2v_reg;
  assign mem[2360] = mem_2360_sv2v_reg;
  assign mem[2359] = mem_2359_sv2v_reg;
  assign mem[2358] = mem_2358_sv2v_reg;
  assign mem[2357] = mem_2357_sv2v_reg;
  assign mem[2356] = mem_2356_sv2v_reg;
  assign mem[2355] = mem_2355_sv2v_reg;
  assign mem[2354] = mem_2354_sv2v_reg;
  assign mem[2353] = mem_2353_sv2v_reg;
  assign mem[2352] = mem_2352_sv2v_reg;
  assign mem[2351] = mem_2351_sv2v_reg;
  assign mem[2350] = mem_2350_sv2v_reg;
  assign mem[2349] = mem_2349_sv2v_reg;
  assign mem[2348] = mem_2348_sv2v_reg;
  assign mem[2347] = mem_2347_sv2v_reg;
  assign mem[2346] = mem_2346_sv2v_reg;
  assign mem[2345] = mem_2345_sv2v_reg;
  assign mem[2344] = mem_2344_sv2v_reg;
  assign mem[2343] = mem_2343_sv2v_reg;
  assign mem[2342] = mem_2342_sv2v_reg;
  assign mem[2341] = mem_2341_sv2v_reg;
  assign mem[2340] = mem_2340_sv2v_reg;
  assign mem[2339] = mem_2339_sv2v_reg;
  assign mem[2338] = mem_2338_sv2v_reg;
  assign mem[2337] = mem_2337_sv2v_reg;
  assign mem[2336] = mem_2336_sv2v_reg;
  assign mem[2335] = mem_2335_sv2v_reg;
  assign mem[2334] = mem_2334_sv2v_reg;
  assign mem[2333] = mem_2333_sv2v_reg;
  assign mem[2332] = mem_2332_sv2v_reg;
  assign mem[2331] = mem_2331_sv2v_reg;
  assign mem[2330] = mem_2330_sv2v_reg;
  assign mem[2329] = mem_2329_sv2v_reg;
  assign mem[2328] = mem_2328_sv2v_reg;
  assign mem[2327] = mem_2327_sv2v_reg;
  assign mem[2326] = mem_2326_sv2v_reg;
  assign mem[2325] = mem_2325_sv2v_reg;
  assign mem[2324] = mem_2324_sv2v_reg;
  assign mem[2323] = mem_2323_sv2v_reg;
  assign mem[2322] = mem_2322_sv2v_reg;
  assign mem[2321] = mem_2321_sv2v_reg;
  assign mem[2320] = mem_2320_sv2v_reg;
  assign mem[2319] = mem_2319_sv2v_reg;
  assign mem[2318] = mem_2318_sv2v_reg;
  assign mem[2317] = mem_2317_sv2v_reg;
  assign mem[2316] = mem_2316_sv2v_reg;
  assign mem[2315] = mem_2315_sv2v_reg;
  assign mem[2314] = mem_2314_sv2v_reg;
  assign mem[2313] = mem_2313_sv2v_reg;
  assign mem[2312] = mem_2312_sv2v_reg;
  assign mem[2311] = mem_2311_sv2v_reg;
  assign mem[2310] = mem_2310_sv2v_reg;
  assign mem[2309] = mem_2309_sv2v_reg;
  assign mem[2308] = mem_2308_sv2v_reg;
  assign mem[2307] = mem_2307_sv2v_reg;
  assign mem[2306] = mem_2306_sv2v_reg;
  assign mem[2305] = mem_2305_sv2v_reg;
  assign mem[2304] = mem_2304_sv2v_reg;
  assign mem[2303] = mem_2303_sv2v_reg;
  assign mem[2302] = mem_2302_sv2v_reg;
  assign mem[2301] = mem_2301_sv2v_reg;
  assign mem[2300] = mem_2300_sv2v_reg;
  assign mem[2299] = mem_2299_sv2v_reg;
  assign mem[2298] = mem_2298_sv2v_reg;
  assign mem[2297] = mem_2297_sv2v_reg;
  assign mem[2296] = mem_2296_sv2v_reg;
  assign mem[2295] = mem_2295_sv2v_reg;
  assign mem[2294] = mem_2294_sv2v_reg;
  assign mem[2293] = mem_2293_sv2v_reg;
  assign mem[2292] = mem_2292_sv2v_reg;
  assign mem[2291] = mem_2291_sv2v_reg;
  assign mem[2290] = mem_2290_sv2v_reg;
  assign mem[2289] = mem_2289_sv2v_reg;
  assign mem[2288] = mem_2288_sv2v_reg;
  assign mem[2287] = mem_2287_sv2v_reg;
  assign mem[2286] = mem_2286_sv2v_reg;
  assign mem[2285] = mem_2285_sv2v_reg;
  assign mem[2284] = mem_2284_sv2v_reg;
  assign mem[2283] = mem_2283_sv2v_reg;
  assign mem[2282] = mem_2282_sv2v_reg;
  assign mem[2281] = mem_2281_sv2v_reg;
  assign mem[2280] = mem_2280_sv2v_reg;
  assign mem[2279] = mem_2279_sv2v_reg;
  assign mem[2278] = mem_2278_sv2v_reg;
  assign mem[2277] = mem_2277_sv2v_reg;
  assign mem[2276] = mem_2276_sv2v_reg;
  assign mem[2275] = mem_2275_sv2v_reg;
  assign mem[2274] = mem_2274_sv2v_reg;
  assign mem[2273] = mem_2273_sv2v_reg;
  assign mem[2272] = mem_2272_sv2v_reg;
  assign mem[2271] = mem_2271_sv2v_reg;
  assign mem[2270] = mem_2270_sv2v_reg;
  assign mem[2269] = mem_2269_sv2v_reg;
  assign mem[2268] = mem_2268_sv2v_reg;
  assign mem[2267] = mem_2267_sv2v_reg;
  assign mem[2266] = mem_2266_sv2v_reg;
  assign mem[2265] = mem_2265_sv2v_reg;
  assign mem[2264] = mem_2264_sv2v_reg;
  assign mem[2263] = mem_2263_sv2v_reg;
  assign mem[2262] = mem_2262_sv2v_reg;
  assign mem[2261] = mem_2261_sv2v_reg;
  assign mem[2260] = mem_2260_sv2v_reg;
  assign mem[2259] = mem_2259_sv2v_reg;
  assign mem[2258] = mem_2258_sv2v_reg;
  assign mem[2257] = mem_2257_sv2v_reg;
  assign mem[2256] = mem_2256_sv2v_reg;
  assign mem[2255] = mem_2255_sv2v_reg;
  assign mem[2254] = mem_2254_sv2v_reg;
  assign mem[2253] = mem_2253_sv2v_reg;
  assign mem[2252] = mem_2252_sv2v_reg;
  assign mem[2251] = mem_2251_sv2v_reg;
  assign mem[2250] = mem_2250_sv2v_reg;
  assign mem[2249] = mem_2249_sv2v_reg;
  assign mem[2248] = mem_2248_sv2v_reg;
  assign mem[2247] = mem_2247_sv2v_reg;
  assign mem[2246] = mem_2246_sv2v_reg;
  assign mem[2245] = mem_2245_sv2v_reg;
  assign mem[2244] = mem_2244_sv2v_reg;
  assign mem[2243] = mem_2243_sv2v_reg;
  assign mem[2242] = mem_2242_sv2v_reg;
  assign mem[2241] = mem_2241_sv2v_reg;
  assign mem[2240] = mem_2240_sv2v_reg;
  assign mem[2239] = mem_2239_sv2v_reg;
  assign mem[2238] = mem_2238_sv2v_reg;
  assign mem[2237] = mem_2237_sv2v_reg;
  assign mem[2236] = mem_2236_sv2v_reg;
  assign mem[2235] = mem_2235_sv2v_reg;
  assign mem[2234] = mem_2234_sv2v_reg;
  assign mem[2233] = mem_2233_sv2v_reg;
  assign mem[2232] = mem_2232_sv2v_reg;
  assign mem[2231] = mem_2231_sv2v_reg;
  assign mem[2230] = mem_2230_sv2v_reg;
  assign mem[2229] = mem_2229_sv2v_reg;
  assign mem[2228] = mem_2228_sv2v_reg;
  assign mem[2227] = mem_2227_sv2v_reg;
  assign mem[2226] = mem_2226_sv2v_reg;
  assign mem[2225] = mem_2225_sv2v_reg;
  assign mem[2224] = mem_2224_sv2v_reg;
  assign mem[2223] = mem_2223_sv2v_reg;
  assign mem[2222] = mem_2222_sv2v_reg;
  assign mem[2221] = mem_2221_sv2v_reg;
  assign mem[2220] = mem_2220_sv2v_reg;
  assign mem[2219] = mem_2219_sv2v_reg;
  assign mem[2218] = mem_2218_sv2v_reg;
  assign mem[2217] = mem_2217_sv2v_reg;
  assign mem[2216] = mem_2216_sv2v_reg;
  assign mem[2215] = mem_2215_sv2v_reg;
  assign mem[2214] = mem_2214_sv2v_reg;
  assign mem[2213] = mem_2213_sv2v_reg;
  assign mem[2212] = mem_2212_sv2v_reg;
  assign mem[2211] = mem_2211_sv2v_reg;
  assign mem[2210] = mem_2210_sv2v_reg;
  assign mem[2209] = mem_2209_sv2v_reg;
  assign mem[2208] = mem_2208_sv2v_reg;
  assign mem[2207] = mem_2207_sv2v_reg;
  assign mem[2206] = mem_2206_sv2v_reg;
  assign mem[2205] = mem_2205_sv2v_reg;
  assign mem[2204] = mem_2204_sv2v_reg;
  assign mem[2203] = mem_2203_sv2v_reg;
  assign mem[2202] = mem_2202_sv2v_reg;
  assign mem[2201] = mem_2201_sv2v_reg;
  assign mem[2200] = mem_2200_sv2v_reg;
  assign mem[2199] = mem_2199_sv2v_reg;
  assign mem[2198] = mem_2198_sv2v_reg;
  assign mem[2197] = mem_2197_sv2v_reg;
  assign mem[2196] = mem_2196_sv2v_reg;
  assign mem[2195] = mem_2195_sv2v_reg;
  assign mem[2194] = mem_2194_sv2v_reg;
  assign mem[2193] = mem_2193_sv2v_reg;
  assign mem[2192] = mem_2192_sv2v_reg;
  assign mem[2191] = mem_2191_sv2v_reg;
  assign mem[2190] = mem_2190_sv2v_reg;
  assign mem[2189] = mem_2189_sv2v_reg;
  assign mem[2188] = mem_2188_sv2v_reg;
  assign mem[2187] = mem_2187_sv2v_reg;
  assign mem[2186] = mem_2186_sv2v_reg;
  assign mem[2185] = mem_2185_sv2v_reg;
  assign mem[2184] = mem_2184_sv2v_reg;
  assign mem[2183] = mem_2183_sv2v_reg;
  assign mem[2182] = mem_2182_sv2v_reg;
  assign mem[2181] = mem_2181_sv2v_reg;
  assign mem[2180] = mem_2180_sv2v_reg;
  assign mem[2179] = mem_2179_sv2v_reg;
  assign mem[2178] = mem_2178_sv2v_reg;
  assign mem[2177] = mem_2177_sv2v_reg;
  assign mem[2176] = mem_2176_sv2v_reg;
  assign mem[2175] = mem_2175_sv2v_reg;
  assign mem[2174] = mem_2174_sv2v_reg;
  assign mem[2173] = mem_2173_sv2v_reg;
  assign mem[2172] = mem_2172_sv2v_reg;
  assign mem[2171] = mem_2171_sv2v_reg;
  assign mem[2170] = mem_2170_sv2v_reg;
  assign mem[2169] = mem_2169_sv2v_reg;
  assign mem[2168] = mem_2168_sv2v_reg;
  assign mem[2167] = mem_2167_sv2v_reg;
  assign mem[2166] = mem_2166_sv2v_reg;
  assign mem[2165] = mem_2165_sv2v_reg;
  assign mem[2164] = mem_2164_sv2v_reg;
  assign mem[2163] = mem_2163_sv2v_reg;
  assign mem[2162] = mem_2162_sv2v_reg;
  assign mem[2161] = mem_2161_sv2v_reg;
  assign mem[2160] = mem_2160_sv2v_reg;
  assign mem[2159] = mem_2159_sv2v_reg;
  assign mem[2158] = mem_2158_sv2v_reg;
  assign mem[2157] = mem_2157_sv2v_reg;
  assign mem[2156] = mem_2156_sv2v_reg;
  assign mem[2155] = mem_2155_sv2v_reg;
  assign mem[2154] = mem_2154_sv2v_reg;
  assign mem[2153] = mem_2153_sv2v_reg;
  assign mem[2152] = mem_2152_sv2v_reg;
  assign mem[2151] = mem_2151_sv2v_reg;
  assign mem[2150] = mem_2150_sv2v_reg;
  assign mem[2149] = mem_2149_sv2v_reg;
  assign mem[2148] = mem_2148_sv2v_reg;
  assign mem[2147] = mem_2147_sv2v_reg;
  assign mem[2146] = mem_2146_sv2v_reg;
  assign mem[2145] = mem_2145_sv2v_reg;
  assign mem[2144] = mem_2144_sv2v_reg;
  assign mem[2143] = mem_2143_sv2v_reg;
  assign mem[2142] = mem_2142_sv2v_reg;
  assign mem[2141] = mem_2141_sv2v_reg;
  assign mem[2140] = mem_2140_sv2v_reg;
  assign mem[2139] = mem_2139_sv2v_reg;
  assign mem[2138] = mem_2138_sv2v_reg;
  assign mem[2137] = mem_2137_sv2v_reg;
  assign mem[2136] = mem_2136_sv2v_reg;
  assign mem[2135] = mem_2135_sv2v_reg;
  assign mem[2134] = mem_2134_sv2v_reg;
  assign mem[2133] = mem_2133_sv2v_reg;
  assign mem[2132] = mem_2132_sv2v_reg;
  assign mem[2131] = mem_2131_sv2v_reg;
  assign mem[2130] = mem_2130_sv2v_reg;
  assign mem[2129] = mem_2129_sv2v_reg;
  assign mem[2128] = mem_2128_sv2v_reg;
  assign mem[2127] = mem_2127_sv2v_reg;
  assign mem[2126] = mem_2126_sv2v_reg;
  assign mem[2125] = mem_2125_sv2v_reg;
  assign mem[2124] = mem_2124_sv2v_reg;
  assign mem[2123] = mem_2123_sv2v_reg;
  assign mem[2122] = mem_2122_sv2v_reg;
  assign mem[2121] = mem_2121_sv2v_reg;
  assign mem[2120] = mem_2120_sv2v_reg;
  assign mem[2119] = mem_2119_sv2v_reg;
  assign mem[2118] = mem_2118_sv2v_reg;
  assign mem[2117] = mem_2117_sv2v_reg;
  assign mem[2116] = mem_2116_sv2v_reg;
  assign mem[2115] = mem_2115_sv2v_reg;
  assign mem[2114] = mem_2114_sv2v_reg;
  assign mem[2113] = mem_2113_sv2v_reg;
  assign mem[2112] = mem_2112_sv2v_reg;
  assign mem[2111] = mem_2111_sv2v_reg;
  assign mem[2110] = mem_2110_sv2v_reg;
  assign mem[2109] = mem_2109_sv2v_reg;
  assign mem[2108] = mem_2108_sv2v_reg;
  assign mem[2107] = mem_2107_sv2v_reg;
  assign mem[2106] = mem_2106_sv2v_reg;
  assign mem[2105] = mem_2105_sv2v_reg;
  assign mem[2104] = mem_2104_sv2v_reg;
  assign mem[2103] = mem_2103_sv2v_reg;
  assign mem[2102] = mem_2102_sv2v_reg;
  assign mem[2101] = mem_2101_sv2v_reg;
  assign mem[2100] = mem_2100_sv2v_reg;
  assign mem[2099] = mem_2099_sv2v_reg;
  assign mem[2098] = mem_2098_sv2v_reg;
  assign mem[2097] = mem_2097_sv2v_reg;
  assign mem[2096] = mem_2096_sv2v_reg;
  assign mem[2095] = mem_2095_sv2v_reg;
  assign mem[2094] = mem_2094_sv2v_reg;
  assign mem[2093] = mem_2093_sv2v_reg;
  assign mem[2092] = mem_2092_sv2v_reg;
  assign mem[2091] = mem_2091_sv2v_reg;
  assign mem[2090] = mem_2090_sv2v_reg;
  assign mem[2089] = mem_2089_sv2v_reg;
  assign mem[2088] = mem_2088_sv2v_reg;
  assign mem[2087] = mem_2087_sv2v_reg;
  assign mem[2086] = mem_2086_sv2v_reg;
  assign mem[2085] = mem_2085_sv2v_reg;
  assign mem[2084] = mem_2084_sv2v_reg;
  assign mem[2083] = mem_2083_sv2v_reg;
  assign mem[2082] = mem_2082_sv2v_reg;
  assign mem[2081] = mem_2081_sv2v_reg;
  assign mem[2080] = mem_2080_sv2v_reg;
  assign mem[2079] = mem_2079_sv2v_reg;
  assign mem[2078] = mem_2078_sv2v_reg;
  assign mem[2077] = mem_2077_sv2v_reg;
  assign mem[2076] = mem_2076_sv2v_reg;
  assign mem[2075] = mem_2075_sv2v_reg;
  assign mem[2074] = mem_2074_sv2v_reg;
  assign mem[2073] = mem_2073_sv2v_reg;
  assign mem[2072] = mem_2072_sv2v_reg;
  assign mem[2071] = mem_2071_sv2v_reg;
  assign mem[2070] = mem_2070_sv2v_reg;
  assign mem[2069] = mem_2069_sv2v_reg;
  assign mem[2068] = mem_2068_sv2v_reg;
  assign mem[2067] = mem_2067_sv2v_reg;
  assign mem[2066] = mem_2066_sv2v_reg;
  assign mem[2065] = mem_2065_sv2v_reg;
  assign mem[2064] = mem_2064_sv2v_reg;
  assign mem[2063] = mem_2063_sv2v_reg;
  assign mem[2062] = mem_2062_sv2v_reg;
  assign mem[2061] = mem_2061_sv2v_reg;
  assign mem[2060] = mem_2060_sv2v_reg;
  assign mem[2059] = mem_2059_sv2v_reg;
  assign mem[2058] = mem_2058_sv2v_reg;
  assign mem[2057] = mem_2057_sv2v_reg;
  assign mem[2056] = mem_2056_sv2v_reg;
  assign mem[2055] = mem_2055_sv2v_reg;
  assign mem[2054] = mem_2054_sv2v_reg;
  assign mem[2053] = mem_2053_sv2v_reg;
  assign mem[2052] = mem_2052_sv2v_reg;
  assign mem[2051] = mem_2051_sv2v_reg;
  assign mem[2050] = mem_2050_sv2v_reg;
  assign mem[2049] = mem_2049_sv2v_reg;
  assign mem[2048] = mem_2048_sv2v_reg;
  assign mem[2047] = mem_2047_sv2v_reg;
  assign mem[2046] = mem_2046_sv2v_reg;
  assign mem[2045] = mem_2045_sv2v_reg;
  assign mem[2044] = mem_2044_sv2v_reg;
  assign mem[2043] = mem_2043_sv2v_reg;
  assign mem[2042] = mem_2042_sv2v_reg;
  assign mem[2041] = mem_2041_sv2v_reg;
  assign mem[2040] = mem_2040_sv2v_reg;
  assign mem[2039] = mem_2039_sv2v_reg;
  assign mem[2038] = mem_2038_sv2v_reg;
  assign mem[2037] = mem_2037_sv2v_reg;
  assign mem[2036] = mem_2036_sv2v_reg;
  assign mem[2035] = mem_2035_sv2v_reg;
  assign mem[2034] = mem_2034_sv2v_reg;
  assign mem[2033] = mem_2033_sv2v_reg;
  assign mem[2032] = mem_2032_sv2v_reg;
  assign mem[2031] = mem_2031_sv2v_reg;
  assign mem[2030] = mem_2030_sv2v_reg;
  assign mem[2029] = mem_2029_sv2v_reg;
  assign mem[2028] = mem_2028_sv2v_reg;
  assign mem[2027] = mem_2027_sv2v_reg;
  assign mem[2026] = mem_2026_sv2v_reg;
  assign mem[2025] = mem_2025_sv2v_reg;
  assign mem[2024] = mem_2024_sv2v_reg;
  assign mem[2023] = mem_2023_sv2v_reg;
  assign mem[2022] = mem_2022_sv2v_reg;
  assign mem[2021] = mem_2021_sv2v_reg;
  assign mem[2020] = mem_2020_sv2v_reg;
  assign mem[2019] = mem_2019_sv2v_reg;
  assign mem[2018] = mem_2018_sv2v_reg;
  assign mem[2017] = mem_2017_sv2v_reg;
  assign mem[2016] = mem_2016_sv2v_reg;
  assign mem[2015] = mem_2015_sv2v_reg;
  assign mem[2014] = mem_2014_sv2v_reg;
  assign mem[2013] = mem_2013_sv2v_reg;
  assign mem[2012] = mem_2012_sv2v_reg;
  assign mem[2011] = mem_2011_sv2v_reg;
  assign mem[2010] = mem_2010_sv2v_reg;
  assign mem[2009] = mem_2009_sv2v_reg;
  assign mem[2008] = mem_2008_sv2v_reg;
  assign mem[2007] = mem_2007_sv2v_reg;
  assign mem[2006] = mem_2006_sv2v_reg;
  assign mem[2005] = mem_2005_sv2v_reg;
  assign mem[2004] = mem_2004_sv2v_reg;
  assign mem[2003] = mem_2003_sv2v_reg;
  assign mem[2002] = mem_2002_sv2v_reg;
  assign mem[2001] = mem_2001_sv2v_reg;
  assign mem[2000] = mem_2000_sv2v_reg;
  assign mem[1999] = mem_1999_sv2v_reg;
  assign mem[1998] = mem_1998_sv2v_reg;
  assign mem[1997] = mem_1997_sv2v_reg;
  assign mem[1996] = mem_1996_sv2v_reg;
  assign mem[1995] = mem_1995_sv2v_reg;
  assign mem[1994] = mem_1994_sv2v_reg;
  assign mem[1993] = mem_1993_sv2v_reg;
  assign mem[1992] = mem_1992_sv2v_reg;
  assign mem[1991] = mem_1991_sv2v_reg;
  assign mem[1990] = mem_1990_sv2v_reg;
  assign mem[1989] = mem_1989_sv2v_reg;
  assign mem[1988] = mem_1988_sv2v_reg;
  assign mem[1987] = mem_1987_sv2v_reg;
  assign mem[1986] = mem_1986_sv2v_reg;
  assign mem[1985] = mem_1985_sv2v_reg;
  assign mem[1984] = mem_1984_sv2v_reg;
  assign mem[1983] = mem_1983_sv2v_reg;
  assign mem[1982] = mem_1982_sv2v_reg;
  assign mem[1981] = mem_1981_sv2v_reg;
  assign mem[1980] = mem_1980_sv2v_reg;
  assign mem[1979] = mem_1979_sv2v_reg;
  assign mem[1978] = mem_1978_sv2v_reg;
  assign mem[1977] = mem_1977_sv2v_reg;
  assign mem[1976] = mem_1976_sv2v_reg;
  assign mem[1975] = mem_1975_sv2v_reg;
  assign mem[1974] = mem_1974_sv2v_reg;
  assign mem[1973] = mem_1973_sv2v_reg;
  assign mem[1972] = mem_1972_sv2v_reg;
  assign mem[1971] = mem_1971_sv2v_reg;
  assign mem[1970] = mem_1970_sv2v_reg;
  assign mem[1969] = mem_1969_sv2v_reg;
  assign mem[1968] = mem_1968_sv2v_reg;
  assign mem[1967] = mem_1967_sv2v_reg;
  assign mem[1966] = mem_1966_sv2v_reg;
  assign mem[1965] = mem_1965_sv2v_reg;
  assign mem[1964] = mem_1964_sv2v_reg;
  assign mem[1963] = mem_1963_sv2v_reg;
  assign mem[1962] = mem_1962_sv2v_reg;
  assign mem[1961] = mem_1961_sv2v_reg;
  assign mem[1960] = mem_1960_sv2v_reg;
  assign mem[1959] = mem_1959_sv2v_reg;
  assign mem[1958] = mem_1958_sv2v_reg;
  assign mem[1957] = mem_1957_sv2v_reg;
  assign mem[1956] = mem_1956_sv2v_reg;
  assign mem[1955] = mem_1955_sv2v_reg;
  assign mem[1954] = mem_1954_sv2v_reg;
  assign mem[1953] = mem_1953_sv2v_reg;
  assign mem[1952] = mem_1952_sv2v_reg;
  assign mem[1951] = mem_1951_sv2v_reg;
  assign mem[1950] = mem_1950_sv2v_reg;
  assign mem[1949] = mem_1949_sv2v_reg;
  assign mem[1948] = mem_1948_sv2v_reg;
  assign mem[1947] = mem_1947_sv2v_reg;
  assign mem[1946] = mem_1946_sv2v_reg;
  assign mem[1945] = mem_1945_sv2v_reg;
  assign mem[1944] = mem_1944_sv2v_reg;
  assign mem[1943] = mem_1943_sv2v_reg;
  assign mem[1942] = mem_1942_sv2v_reg;
  assign mem[1941] = mem_1941_sv2v_reg;
  assign mem[1940] = mem_1940_sv2v_reg;
  assign mem[1939] = mem_1939_sv2v_reg;
  assign mem[1938] = mem_1938_sv2v_reg;
  assign mem[1937] = mem_1937_sv2v_reg;
  assign mem[1936] = mem_1936_sv2v_reg;
  assign mem[1935] = mem_1935_sv2v_reg;
  assign mem[1934] = mem_1934_sv2v_reg;
  assign mem[1933] = mem_1933_sv2v_reg;
  assign mem[1932] = mem_1932_sv2v_reg;
  assign mem[1931] = mem_1931_sv2v_reg;
  assign mem[1930] = mem_1930_sv2v_reg;
  assign mem[1929] = mem_1929_sv2v_reg;
  assign mem[1928] = mem_1928_sv2v_reg;
  assign mem[1927] = mem_1927_sv2v_reg;
  assign mem[1926] = mem_1926_sv2v_reg;
  assign mem[1925] = mem_1925_sv2v_reg;
  assign mem[1924] = mem_1924_sv2v_reg;
  assign mem[1923] = mem_1923_sv2v_reg;
  assign mem[1922] = mem_1922_sv2v_reg;
  assign mem[1921] = mem_1921_sv2v_reg;
  assign mem[1920] = mem_1920_sv2v_reg;
  assign mem[1919] = mem_1919_sv2v_reg;
  assign mem[1918] = mem_1918_sv2v_reg;
  assign mem[1917] = mem_1917_sv2v_reg;
  assign mem[1916] = mem_1916_sv2v_reg;
  assign mem[1915] = mem_1915_sv2v_reg;
  assign mem[1914] = mem_1914_sv2v_reg;
  assign mem[1913] = mem_1913_sv2v_reg;
  assign mem[1912] = mem_1912_sv2v_reg;
  assign mem[1911] = mem_1911_sv2v_reg;
  assign mem[1910] = mem_1910_sv2v_reg;
  assign mem[1909] = mem_1909_sv2v_reg;
  assign mem[1908] = mem_1908_sv2v_reg;
  assign mem[1907] = mem_1907_sv2v_reg;
  assign mem[1906] = mem_1906_sv2v_reg;
  assign mem[1905] = mem_1905_sv2v_reg;
  assign mem[1904] = mem_1904_sv2v_reg;
  assign mem[1903] = mem_1903_sv2v_reg;
  assign mem[1902] = mem_1902_sv2v_reg;
  assign mem[1901] = mem_1901_sv2v_reg;
  assign mem[1900] = mem_1900_sv2v_reg;
  assign mem[1899] = mem_1899_sv2v_reg;
  assign mem[1898] = mem_1898_sv2v_reg;
  assign mem[1897] = mem_1897_sv2v_reg;
  assign mem[1896] = mem_1896_sv2v_reg;
  assign mem[1895] = mem_1895_sv2v_reg;
  assign mem[1894] = mem_1894_sv2v_reg;
  assign mem[1893] = mem_1893_sv2v_reg;
  assign mem[1892] = mem_1892_sv2v_reg;
  assign mem[1891] = mem_1891_sv2v_reg;
  assign mem[1890] = mem_1890_sv2v_reg;
  assign mem[1889] = mem_1889_sv2v_reg;
  assign mem[1888] = mem_1888_sv2v_reg;
  assign mem[1887] = mem_1887_sv2v_reg;
  assign mem[1886] = mem_1886_sv2v_reg;
  assign mem[1885] = mem_1885_sv2v_reg;
  assign mem[1884] = mem_1884_sv2v_reg;
  assign mem[1883] = mem_1883_sv2v_reg;
  assign mem[1882] = mem_1882_sv2v_reg;
  assign mem[1881] = mem_1881_sv2v_reg;
  assign mem[1880] = mem_1880_sv2v_reg;
  assign mem[1879] = mem_1879_sv2v_reg;
  assign mem[1878] = mem_1878_sv2v_reg;
  assign mem[1877] = mem_1877_sv2v_reg;
  assign mem[1876] = mem_1876_sv2v_reg;
  assign mem[1875] = mem_1875_sv2v_reg;
  assign mem[1874] = mem_1874_sv2v_reg;
  assign mem[1873] = mem_1873_sv2v_reg;
  assign mem[1872] = mem_1872_sv2v_reg;
  assign mem[1871] = mem_1871_sv2v_reg;
  assign mem[1870] = mem_1870_sv2v_reg;
  assign mem[1869] = mem_1869_sv2v_reg;
  assign mem[1868] = mem_1868_sv2v_reg;
  assign mem[1867] = mem_1867_sv2v_reg;
  assign mem[1866] = mem_1866_sv2v_reg;
  assign mem[1865] = mem_1865_sv2v_reg;
  assign mem[1864] = mem_1864_sv2v_reg;
  assign mem[1863] = mem_1863_sv2v_reg;
  assign mem[1862] = mem_1862_sv2v_reg;
  assign mem[1861] = mem_1861_sv2v_reg;
  assign mem[1860] = mem_1860_sv2v_reg;
  assign mem[1859] = mem_1859_sv2v_reg;
  assign mem[1858] = mem_1858_sv2v_reg;
  assign mem[1857] = mem_1857_sv2v_reg;
  assign mem[1856] = mem_1856_sv2v_reg;
  assign mem[1855] = mem_1855_sv2v_reg;
  assign mem[1854] = mem_1854_sv2v_reg;
  assign mem[1853] = mem_1853_sv2v_reg;
  assign mem[1852] = mem_1852_sv2v_reg;
  assign mem[1851] = mem_1851_sv2v_reg;
  assign mem[1850] = mem_1850_sv2v_reg;
  assign mem[1849] = mem_1849_sv2v_reg;
  assign mem[1848] = mem_1848_sv2v_reg;
  assign mem[1847] = mem_1847_sv2v_reg;
  assign mem[1846] = mem_1846_sv2v_reg;
  assign mem[1845] = mem_1845_sv2v_reg;
  assign mem[1844] = mem_1844_sv2v_reg;
  assign mem[1843] = mem_1843_sv2v_reg;
  assign mem[1842] = mem_1842_sv2v_reg;
  assign mem[1841] = mem_1841_sv2v_reg;
  assign mem[1840] = mem_1840_sv2v_reg;
  assign mem[1839] = mem_1839_sv2v_reg;
  assign mem[1838] = mem_1838_sv2v_reg;
  assign mem[1837] = mem_1837_sv2v_reg;
  assign mem[1836] = mem_1836_sv2v_reg;
  assign mem[1835] = mem_1835_sv2v_reg;
  assign mem[1834] = mem_1834_sv2v_reg;
  assign mem[1833] = mem_1833_sv2v_reg;
  assign mem[1832] = mem_1832_sv2v_reg;
  assign mem[1831] = mem_1831_sv2v_reg;
  assign mem[1830] = mem_1830_sv2v_reg;
  assign mem[1829] = mem_1829_sv2v_reg;
  assign mem[1828] = mem_1828_sv2v_reg;
  assign mem[1827] = mem_1827_sv2v_reg;
  assign mem[1826] = mem_1826_sv2v_reg;
  assign mem[1825] = mem_1825_sv2v_reg;
  assign mem[1824] = mem_1824_sv2v_reg;
  assign mem[1823] = mem_1823_sv2v_reg;
  assign mem[1822] = mem_1822_sv2v_reg;
  assign mem[1821] = mem_1821_sv2v_reg;
  assign mem[1820] = mem_1820_sv2v_reg;
  assign mem[1819] = mem_1819_sv2v_reg;
  assign mem[1818] = mem_1818_sv2v_reg;
  assign mem[1817] = mem_1817_sv2v_reg;
  assign mem[1816] = mem_1816_sv2v_reg;
  assign mem[1815] = mem_1815_sv2v_reg;
  assign mem[1814] = mem_1814_sv2v_reg;
  assign mem[1813] = mem_1813_sv2v_reg;
  assign mem[1812] = mem_1812_sv2v_reg;
  assign mem[1811] = mem_1811_sv2v_reg;
  assign mem[1810] = mem_1810_sv2v_reg;
  assign mem[1809] = mem_1809_sv2v_reg;
  assign mem[1808] = mem_1808_sv2v_reg;
  assign mem[1807] = mem_1807_sv2v_reg;
  assign mem[1806] = mem_1806_sv2v_reg;
  assign mem[1805] = mem_1805_sv2v_reg;
  assign mem[1804] = mem_1804_sv2v_reg;
  assign mem[1803] = mem_1803_sv2v_reg;
  assign mem[1802] = mem_1802_sv2v_reg;
  assign mem[1801] = mem_1801_sv2v_reg;
  assign mem[1800] = mem_1800_sv2v_reg;
  assign mem[1799] = mem_1799_sv2v_reg;
  assign mem[1798] = mem_1798_sv2v_reg;
  assign mem[1797] = mem_1797_sv2v_reg;
  assign mem[1796] = mem_1796_sv2v_reg;
  assign mem[1795] = mem_1795_sv2v_reg;
  assign mem[1794] = mem_1794_sv2v_reg;
  assign mem[1793] = mem_1793_sv2v_reg;
  assign mem[1792] = mem_1792_sv2v_reg;
  assign mem[1791] = mem_1791_sv2v_reg;
  assign mem[1790] = mem_1790_sv2v_reg;
  assign mem[1789] = mem_1789_sv2v_reg;
  assign mem[1788] = mem_1788_sv2v_reg;
  assign mem[1787] = mem_1787_sv2v_reg;
  assign mem[1786] = mem_1786_sv2v_reg;
  assign mem[1785] = mem_1785_sv2v_reg;
  assign mem[1784] = mem_1784_sv2v_reg;
  assign mem[1783] = mem_1783_sv2v_reg;
  assign mem[1782] = mem_1782_sv2v_reg;
  assign mem[1781] = mem_1781_sv2v_reg;
  assign mem[1780] = mem_1780_sv2v_reg;
  assign mem[1779] = mem_1779_sv2v_reg;
  assign mem[1778] = mem_1778_sv2v_reg;
  assign mem[1777] = mem_1777_sv2v_reg;
  assign mem[1776] = mem_1776_sv2v_reg;
  assign mem[1775] = mem_1775_sv2v_reg;
  assign mem[1774] = mem_1774_sv2v_reg;
  assign mem[1773] = mem_1773_sv2v_reg;
  assign mem[1772] = mem_1772_sv2v_reg;
  assign mem[1771] = mem_1771_sv2v_reg;
  assign mem[1770] = mem_1770_sv2v_reg;
  assign mem[1769] = mem_1769_sv2v_reg;
  assign mem[1768] = mem_1768_sv2v_reg;
  assign mem[1767] = mem_1767_sv2v_reg;
  assign mem[1766] = mem_1766_sv2v_reg;
  assign mem[1765] = mem_1765_sv2v_reg;
  assign mem[1764] = mem_1764_sv2v_reg;
  assign mem[1763] = mem_1763_sv2v_reg;
  assign mem[1762] = mem_1762_sv2v_reg;
  assign mem[1761] = mem_1761_sv2v_reg;
  assign mem[1760] = mem_1760_sv2v_reg;
  assign mem[1759] = mem_1759_sv2v_reg;
  assign mem[1758] = mem_1758_sv2v_reg;
  assign mem[1757] = mem_1757_sv2v_reg;
  assign mem[1756] = mem_1756_sv2v_reg;
  assign mem[1755] = mem_1755_sv2v_reg;
  assign mem[1754] = mem_1754_sv2v_reg;
  assign mem[1753] = mem_1753_sv2v_reg;
  assign mem[1752] = mem_1752_sv2v_reg;
  assign mem[1751] = mem_1751_sv2v_reg;
  assign mem[1750] = mem_1750_sv2v_reg;
  assign mem[1749] = mem_1749_sv2v_reg;
  assign mem[1748] = mem_1748_sv2v_reg;
  assign mem[1747] = mem_1747_sv2v_reg;
  assign mem[1746] = mem_1746_sv2v_reg;
  assign mem[1745] = mem_1745_sv2v_reg;
  assign mem[1744] = mem_1744_sv2v_reg;
  assign mem[1743] = mem_1743_sv2v_reg;
  assign mem[1742] = mem_1742_sv2v_reg;
  assign mem[1741] = mem_1741_sv2v_reg;
  assign mem[1740] = mem_1740_sv2v_reg;
  assign mem[1739] = mem_1739_sv2v_reg;
  assign mem[1738] = mem_1738_sv2v_reg;
  assign mem[1737] = mem_1737_sv2v_reg;
  assign mem[1736] = mem_1736_sv2v_reg;
  assign mem[1735] = mem_1735_sv2v_reg;
  assign mem[1734] = mem_1734_sv2v_reg;
  assign mem[1733] = mem_1733_sv2v_reg;
  assign mem[1732] = mem_1732_sv2v_reg;
  assign mem[1731] = mem_1731_sv2v_reg;
  assign mem[1730] = mem_1730_sv2v_reg;
  assign mem[1729] = mem_1729_sv2v_reg;
  assign mem[1728] = mem_1728_sv2v_reg;
  assign mem[1727] = mem_1727_sv2v_reg;
  assign mem[1726] = mem_1726_sv2v_reg;
  assign mem[1725] = mem_1725_sv2v_reg;
  assign mem[1724] = mem_1724_sv2v_reg;
  assign mem[1723] = mem_1723_sv2v_reg;
  assign mem[1722] = mem_1722_sv2v_reg;
  assign mem[1721] = mem_1721_sv2v_reg;
  assign mem[1720] = mem_1720_sv2v_reg;
  assign mem[1719] = mem_1719_sv2v_reg;
  assign mem[1718] = mem_1718_sv2v_reg;
  assign mem[1717] = mem_1717_sv2v_reg;
  assign mem[1716] = mem_1716_sv2v_reg;
  assign mem[1715] = mem_1715_sv2v_reg;
  assign mem[1714] = mem_1714_sv2v_reg;
  assign mem[1713] = mem_1713_sv2v_reg;
  assign mem[1712] = mem_1712_sv2v_reg;
  assign mem[1711] = mem_1711_sv2v_reg;
  assign mem[1710] = mem_1710_sv2v_reg;
  assign mem[1709] = mem_1709_sv2v_reg;
  assign mem[1708] = mem_1708_sv2v_reg;
  assign mem[1707] = mem_1707_sv2v_reg;
  assign mem[1706] = mem_1706_sv2v_reg;
  assign mem[1705] = mem_1705_sv2v_reg;
  assign mem[1704] = mem_1704_sv2v_reg;
  assign mem[1703] = mem_1703_sv2v_reg;
  assign mem[1702] = mem_1702_sv2v_reg;
  assign mem[1701] = mem_1701_sv2v_reg;
  assign mem[1700] = mem_1700_sv2v_reg;
  assign mem[1699] = mem_1699_sv2v_reg;
  assign mem[1698] = mem_1698_sv2v_reg;
  assign mem[1697] = mem_1697_sv2v_reg;
  assign mem[1696] = mem_1696_sv2v_reg;
  assign mem[1695] = mem_1695_sv2v_reg;
  assign mem[1694] = mem_1694_sv2v_reg;
  assign mem[1693] = mem_1693_sv2v_reg;
  assign mem[1692] = mem_1692_sv2v_reg;
  assign mem[1691] = mem_1691_sv2v_reg;
  assign mem[1690] = mem_1690_sv2v_reg;
  assign mem[1689] = mem_1689_sv2v_reg;
  assign mem[1688] = mem_1688_sv2v_reg;
  assign mem[1687] = mem_1687_sv2v_reg;
  assign mem[1686] = mem_1686_sv2v_reg;
  assign mem[1685] = mem_1685_sv2v_reg;
  assign mem[1684] = mem_1684_sv2v_reg;
  assign mem[1683] = mem_1683_sv2v_reg;
  assign mem[1682] = mem_1682_sv2v_reg;
  assign mem[1681] = mem_1681_sv2v_reg;
  assign mem[1680] = mem_1680_sv2v_reg;
  assign mem[1679] = mem_1679_sv2v_reg;
  assign mem[1678] = mem_1678_sv2v_reg;
  assign mem[1677] = mem_1677_sv2v_reg;
  assign mem[1676] = mem_1676_sv2v_reg;
  assign mem[1675] = mem_1675_sv2v_reg;
  assign mem[1674] = mem_1674_sv2v_reg;
  assign mem[1673] = mem_1673_sv2v_reg;
  assign mem[1672] = mem_1672_sv2v_reg;
  assign mem[1671] = mem_1671_sv2v_reg;
  assign mem[1670] = mem_1670_sv2v_reg;
  assign mem[1669] = mem_1669_sv2v_reg;
  assign mem[1668] = mem_1668_sv2v_reg;
  assign mem[1667] = mem_1667_sv2v_reg;
  assign mem[1666] = mem_1666_sv2v_reg;
  assign mem[1665] = mem_1665_sv2v_reg;
  assign mem[1664] = mem_1664_sv2v_reg;
  assign mem[1663] = mem_1663_sv2v_reg;
  assign mem[1662] = mem_1662_sv2v_reg;
  assign mem[1661] = mem_1661_sv2v_reg;
  assign mem[1660] = mem_1660_sv2v_reg;
  assign mem[1659] = mem_1659_sv2v_reg;
  assign mem[1658] = mem_1658_sv2v_reg;
  assign mem[1657] = mem_1657_sv2v_reg;
  assign mem[1656] = mem_1656_sv2v_reg;
  assign mem[1655] = mem_1655_sv2v_reg;
  assign mem[1654] = mem_1654_sv2v_reg;
  assign mem[1653] = mem_1653_sv2v_reg;
  assign mem[1652] = mem_1652_sv2v_reg;
  assign mem[1651] = mem_1651_sv2v_reg;
  assign mem[1650] = mem_1650_sv2v_reg;
  assign mem[1649] = mem_1649_sv2v_reg;
  assign mem[1648] = mem_1648_sv2v_reg;
  assign mem[1647] = mem_1647_sv2v_reg;
  assign mem[1646] = mem_1646_sv2v_reg;
  assign mem[1645] = mem_1645_sv2v_reg;
  assign mem[1644] = mem_1644_sv2v_reg;
  assign mem[1643] = mem_1643_sv2v_reg;
  assign mem[1642] = mem_1642_sv2v_reg;
  assign mem[1641] = mem_1641_sv2v_reg;
  assign mem[1640] = mem_1640_sv2v_reg;
  assign mem[1639] = mem_1639_sv2v_reg;
  assign mem[1638] = mem_1638_sv2v_reg;
  assign mem[1637] = mem_1637_sv2v_reg;
  assign mem[1636] = mem_1636_sv2v_reg;
  assign mem[1635] = mem_1635_sv2v_reg;
  assign mem[1634] = mem_1634_sv2v_reg;
  assign mem[1633] = mem_1633_sv2v_reg;
  assign mem[1632] = mem_1632_sv2v_reg;
  assign mem[1631] = mem_1631_sv2v_reg;
  assign mem[1630] = mem_1630_sv2v_reg;
  assign mem[1629] = mem_1629_sv2v_reg;
  assign mem[1628] = mem_1628_sv2v_reg;
  assign mem[1627] = mem_1627_sv2v_reg;
  assign mem[1626] = mem_1626_sv2v_reg;
  assign mem[1625] = mem_1625_sv2v_reg;
  assign mem[1624] = mem_1624_sv2v_reg;
  assign mem[1623] = mem_1623_sv2v_reg;
  assign mem[1622] = mem_1622_sv2v_reg;
  assign mem[1621] = mem_1621_sv2v_reg;
  assign mem[1620] = mem_1620_sv2v_reg;
  assign mem[1619] = mem_1619_sv2v_reg;
  assign mem[1618] = mem_1618_sv2v_reg;
  assign mem[1617] = mem_1617_sv2v_reg;
  assign mem[1616] = mem_1616_sv2v_reg;
  assign mem[1615] = mem_1615_sv2v_reg;
  assign mem[1614] = mem_1614_sv2v_reg;
  assign mem[1613] = mem_1613_sv2v_reg;
  assign mem[1612] = mem_1612_sv2v_reg;
  assign mem[1611] = mem_1611_sv2v_reg;
  assign mem[1610] = mem_1610_sv2v_reg;
  assign mem[1609] = mem_1609_sv2v_reg;
  assign mem[1608] = mem_1608_sv2v_reg;
  assign mem[1607] = mem_1607_sv2v_reg;
  assign mem[1606] = mem_1606_sv2v_reg;
  assign mem[1605] = mem_1605_sv2v_reg;
  assign mem[1604] = mem_1604_sv2v_reg;
  assign mem[1603] = mem_1603_sv2v_reg;
  assign mem[1602] = mem_1602_sv2v_reg;
  assign mem[1601] = mem_1601_sv2v_reg;
  assign mem[1600] = mem_1600_sv2v_reg;
  assign mem[1599] = mem_1599_sv2v_reg;
  assign mem[1598] = mem_1598_sv2v_reg;
  assign mem[1597] = mem_1597_sv2v_reg;
  assign mem[1596] = mem_1596_sv2v_reg;
  assign mem[1595] = mem_1595_sv2v_reg;
  assign mem[1594] = mem_1594_sv2v_reg;
  assign mem[1593] = mem_1593_sv2v_reg;
  assign mem[1592] = mem_1592_sv2v_reg;
  assign mem[1591] = mem_1591_sv2v_reg;
  assign mem[1590] = mem_1590_sv2v_reg;
  assign mem[1589] = mem_1589_sv2v_reg;
  assign mem[1588] = mem_1588_sv2v_reg;
  assign mem[1587] = mem_1587_sv2v_reg;
  assign mem[1586] = mem_1586_sv2v_reg;
  assign mem[1585] = mem_1585_sv2v_reg;
  assign mem[1584] = mem_1584_sv2v_reg;
  assign mem[1583] = mem_1583_sv2v_reg;
  assign mem[1582] = mem_1582_sv2v_reg;
  assign mem[1581] = mem_1581_sv2v_reg;
  assign mem[1580] = mem_1580_sv2v_reg;
  assign mem[1579] = mem_1579_sv2v_reg;
  assign mem[1578] = mem_1578_sv2v_reg;
  assign mem[1577] = mem_1577_sv2v_reg;
  assign mem[1576] = mem_1576_sv2v_reg;
  assign mem[1575] = mem_1575_sv2v_reg;
  assign mem[1574] = mem_1574_sv2v_reg;
  assign mem[1573] = mem_1573_sv2v_reg;
  assign mem[1572] = mem_1572_sv2v_reg;
  assign mem[1571] = mem_1571_sv2v_reg;
  assign mem[1570] = mem_1570_sv2v_reg;
  assign mem[1569] = mem_1569_sv2v_reg;
  assign mem[1568] = mem_1568_sv2v_reg;
  assign mem[1567] = mem_1567_sv2v_reg;
  assign mem[1566] = mem_1566_sv2v_reg;
  assign mem[1565] = mem_1565_sv2v_reg;
  assign mem[1564] = mem_1564_sv2v_reg;
  assign mem[1563] = mem_1563_sv2v_reg;
  assign mem[1562] = mem_1562_sv2v_reg;
  assign mem[1561] = mem_1561_sv2v_reg;
  assign mem[1560] = mem_1560_sv2v_reg;
  assign mem[1559] = mem_1559_sv2v_reg;
  assign mem[1558] = mem_1558_sv2v_reg;
  assign mem[1557] = mem_1557_sv2v_reg;
  assign mem[1556] = mem_1556_sv2v_reg;
  assign mem[1555] = mem_1555_sv2v_reg;
  assign mem[1554] = mem_1554_sv2v_reg;
  assign mem[1553] = mem_1553_sv2v_reg;
  assign mem[1552] = mem_1552_sv2v_reg;
  assign mem[1551] = mem_1551_sv2v_reg;
  assign mem[1550] = mem_1550_sv2v_reg;
  assign mem[1549] = mem_1549_sv2v_reg;
  assign mem[1548] = mem_1548_sv2v_reg;
  assign mem[1547] = mem_1547_sv2v_reg;
  assign mem[1546] = mem_1546_sv2v_reg;
  assign mem[1545] = mem_1545_sv2v_reg;
  assign mem[1544] = mem_1544_sv2v_reg;
  assign mem[1543] = mem_1543_sv2v_reg;
  assign mem[1542] = mem_1542_sv2v_reg;
  assign mem[1541] = mem_1541_sv2v_reg;
  assign mem[1540] = mem_1540_sv2v_reg;
  assign mem[1539] = mem_1539_sv2v_reg;
  assign mem[1538] = mem_1538_sv2v_reg;
  assign mem[1537] = mem_1537_sv2v_reg;
  assign mem[1536] = mem_1536_sv2v_reg;
  assign mem[1535] = mem_1535_sv2v_reg;
  assign mem[1534] = mem_1534_sv2v_reg;
  assign mem[1533] = mem_1533_sv2v_reg;
  assign mem[1532] = mem_1532_sv2v_reg;
  assign mem[1531] = mem_1531_sv2v_reg;
  assign mem[1530] = mem_1530_sv2v_reg;
  assign mem[1529] = mem_1529_sv2v_reg;
  assign mem[1528] = mem_1528_sv2v_reg;
  assign mem[1527] = mem_1527_sv2v_reg;
  assign mem[1526] = mem_1526_sv2v_reg;
  assign mem[1525] = mem_1525_sv2v_reg;
  assign mem[1524] = mem_1524_sv2v_reg;
  assign mem[1523] = mem_1523_sv2v_reg;
  assign mem[1522] = mem_1522_sv2v_reg;
  assign mem[1521] = mem_1521_sv2v_reg;
  assign mem[1520] = mem_1520_sv2v_reg;
  assign mem[1519] = mem_1519_sv2v_reg;
  assign mem[1518] = mem_1518_sv2v_reg;
  assign mem[1517] = mem_1517_sv2v_reg;
  assign mem[1516] = mem_1516_sv2v_reg;
  assign mem[1515] = mem_1515_sv2v_reg;
  assign mem[1514] = mem_1514_sv2v_reg;
  assign mem[1513] = mem_1513_sv2v_reg;
  assign mem[1512] = mem_1512_sv2v_reg;
  assign mem[1511] = mem_1511_sv2v_reg;
  assign mem[1510] = mem_1510_sv2v_reg;
  assign mem[1509] = mem_1509_sv2v_reg;
  assign mem[1508] = mem_1508_sv2v_reg;
  assign mem[1507] = mem_1507_sv2v_reg;
  assign mem[1506] = mem_1506_sv2v_reg;
  assign mem[1505] = mem_1505_sv2v_reg;
  assign mem[1504] = mem_1504_sv2v_reg;
  assign mem[1503] = mem_1503_sv2v_reg;
  assign mem[1502] = mem_1502_sv2v_reg;
  assign mem[1501] = mem_1501_sv2v_reg;
  assign mem[1500] = mem_1500_sv2v_reg;
  assign mem[1499] = mem_1499_sv2v_reg;
  assign mem[1498] = mem_1498_sv2v_reg;
  assign mem[1497] = mem_1497_sv2v_reg;
  assign mem[1496] = mem_1496_sv2v_reg;
  assign mem[1495] = mem_1495_sv2v_reg;
  assign mem[1494] = mem_1494_sv2v_reg;
  assign mem[1493] = mem_1493_sv2v_reg;
  assign mem[1492] = mem_1492_sv2v_reg;
  assign mem[1491] = mem_1491_sv2v_reg;
  assign mem[1490] = mem_1490_sv2v_reg;
  assign mem[1489] = mem_1489_sv2v_reg;
  assign mem[1488] = mem_1488_sv2v_reg;
  assign mem[1487] = mem_1487_sv2v_reg;
  assign mem[1486] = mem_1486_sv2v_reg;
  assign mem[1485] = mem_1485_sv2v_reg;
  assign mem[1484] = mem_1484_sv2v_reg;
  assign mem[1483] = mem_1483_sv2v_reg;
  assign mem[1482] = mem_1482_sv2v_reg;
  assign mem[1481] = mem_1481_sv2v_reg;
  assign mem[1480] = mem_1480_sv2v_reg;
  assign mem[1479] = mem_1479_sv2v_reg;
  assign mem[1478] = mem_1478_sv2v_reg;
  assign mem[1477] = mem_1477_sv2v_reg;
  assign mem[1476] = mem_1476_sv2v_reg;
  assign mem[1475] = mem_1475_sv2v_reg;
  assign mem[1474] = mem_1474_sv2v_reg;
  assign mem[1473] = mem_1473_sv2v_reg;
  assign mem[1472] = mem_1472_sv2v_reg;
  assign mem[1471] = mem_1471_sv2v_reg;
  assign mem[1470] = mem_1470_sv2v_reg;
  assign mem[1469] = mem_1469_sv2v_reg;
  assign mem[1468] = mem_1468_sv2v_reg;
  assign mem[1467] = mem_1467_sv2v_reg;
  assign mem[1466] = mem_1466_sv2v_reg;
  assign mem[1465] = mem_1465_sv2v_reg;
  assign mem[1464] = mem_1464_sv2v_reg;
  assign mem[1463] = mem_1463_sv2v_reg;
  assign mem[1462] = mem_1462_sv2v_reg;
  assign mem[1461] = mem_1461_sv2v_reg;
  assign mem[1460] = mem_1460_sv2v_reg;
  assign mem[1459] = mem_1459_sv2v_reg;
  assign mem[1458] = mem_1458_sv2v_reg;
  assign mem[1457] = mem_1457_sv2v_reg;
  assign mem[1456] = mem_1456_sv2v_reg;
  assign mem[1455] = mem_1455_sv2v_reg;
  assign mem[1454] = mem_1454_sv2v_reg;
  assign mem[1453] = mem_1453_sv2v_reg;
  assign mem[1452] = mem_1452_sv2v_reg;
  assign mem[1451] = mem_1451_sv2v_reg;
  assign mem[1450] = mem_1450_sv2v_reg;
  assign mem[1449] = mem_1449_sv2v_reg;
  assign mem[1448] = mem_1448_sv2v_reg;
  assign mem[1447] = mem_1447_sv2v_reg;
  assign mem[1446] = mem_1446_sv2v_reg;
  assign mem[1445] = mem_1445_sv2v_reg;
  assign mem[1444] = mem_1444_sv2v_reg;
  assign mem[1443] = mem_1443_sv2v_reg;
  assign mem[1442] = mem_1442_sv2v_reg;
  assign mem[1441] = mem_1441_sv2v_reg;
  assign mem[1440] = mem_1440_sv2v_reg;
  assign mem[1439] = mem_1439_sv2v_reg;
  assign mem[1438] = mem_1438_sv2v_reg;
  assign mem[1437] = mem_1437_sv2v_reg;
  assign mem[1436] = mem_1436_sv2v_reg;
  assign mem[1435] = mem_1435_sv2v_reg;
  assign mem[1434] = mem_1434_sv2v_reg;
  assign mem[1433] = mem_1433_sv2v_reg;
  assign mem[1432] = mem_1432_sv2v_reg;
  assign mem[1431] = mem_1431_sv2v_reg;
  assign mem[1430] = mem_1430_sv2v_reg;
  assign mem[1429] = mem_1429_sv2v_reg;
  assign mem[1428] = mem_1428_sv2v_reg;
  assign mem[1427] = mem_1427_sv2v_reg;
  assign mem[1426] = mem_1426_sv2v_reg;
  assign mem[1425] = mem_1425_sv2v_reg;
  assign mem[1424] = mem_1424_sv2v_reg;
  assign mem[1423] = mem_1423_sv2v_reg;
  assign mem[1422] = mem_1422_sv2v_reg;
  assign mem[1421] = mem_1421_sv2v_reg;
  assign mem[1420] = mem_1420_sv2v_reg;
  assign mem[1419] = mem_1419_sv2v_reg;
  assign mem[1418] = mem_1418_sv2v_reg;
  assign mem[1417] = mem_1417_sv2v_reg;
  assign mem[1416] = mem_1416_sv2v_reg;
  assign mem[1415] = mem_1415_sv2v_reg;
  assign mem[1414] = mem_1414_sv2v_reg;
  assign mem[1413] = mem_1413_sv2v_reg;
  assign mem[1412] = mem_1412_sv2v_reg;
  assign mem[1411] = mem_1411_sv2v_reg;
  assign mem[1410] = mem_1410_sv2v_reg;
  assign mem[1409] = mem_1409_sv2v_reg;
  assign mem[1408] = mem_1408_sv2v_reg;
  assign mem[1407] = mem_1407_sv2v_reg;
  assign mem[1406] = mem_1406_sv2v_reg;
  assign mem[1405] = mem_1405_sv2v_reg;
  assign mem[1404] = mem_1404_sv2v_reg;
  assign mem[1403] = mem_1403_sv2v_reg;
  assign mem[1402] = mem_1402_sv2v_reg;
  assign mem[1401] = mem_1401_sv2v_reg;
  assign mem[1400] = mem_1400_sv2v_reg;
  assign mem[1399] = mem_1399_sv2v_reg;
  assign mem[1398] = mem_1398_sv2v_reg;
  assign mem[1397] = mem_1397_sv2v_reg;
  assign mem[1396] = mem_1396_sv2v_reg;
  assign mem[1395] = mem_1395_sv2v_reg;
  assign mem[1394] = mem_1394_sv2v_reg;
  assign mem[1393] = mem_1393_sv2v_reg;
  assign mem[1392] = mem_1392_sv2v_reg;
  assign mem[1391] = mem_1391_sv2v_reg;
  assign mem[1390] = mem_1390_sv2v_reg;
  assign mem[1389] = mem_1389_sv2v_reg;
  assign mem[1388] = mem_1388_sv2v_reg;
  assign mem[1387] = mem_1387_sv2v_reg;
  assign mem[1386] = mem_1386_sv2v_reg;
  assign mem[1385] = mem_1385_sv2v_reg;
  assign mem[1384] = mem_1384_sv2v_reg;
  assign mem[1383] = mem_1383_sv2v_reg;
  assign mem[1382] = mem_1382_sv2v_reg;
  assign mem[1381] = mem_1381_sv2v_reg;
  assign mem[1380] = mem_1380_sv2v_reg;
  assign mem[1379] = mem_1379_sv2v_reg;
  assign mem[1378] = mem_1378_sv2v_reg;
  assign mem[1377] = mem_1377_sv2v_reg;
  assign mem[1376] = mem_1376_sv2v_reg;
  assign mem[1375] = mem_1375_sv2v_reg;
  assign mem[1374] = mem_1374_sv2v_reg;
  assign mem[1373] = mem_1373_sv2v_reg;
  assign mem[1372] = mem_1372_sv2v_reg;
  assign mem[1371] = mem_1371_sv2v_reg;
  assign mem[1370] = mem_1370_sv2v_reg;
  assign mem[1369] = mem_1369_sv2v_reg;
  assign mem[1368] = mem_1368_sv2v_reg;
  assign mem[1367] = mem_1367_sv2v_reg;
  assign mem[1366] = mem_1366_sv2v_reg;
  assign mem[1365] = mem_1365_sv2v_reg;
  assign mem[1364] = mem_1364_sv2v_reg;
  assign mem[1363] = mem_1363_sv2v_reg;
  assign mem[1362] = mem_1362_sv2v_reg;
  assign mem[1361] = mem_1361_sv2v_reg;
  assign mem[1360] = mem_1360_sv2v_reg;
  assign mem[1359] = mem_1359_sv2v_reg;
  assign mem[1358] = mem_1358_sv2v_reg;
  assign mem[1357] = mem_1357_sv2v_reg;
  assign mem[1356] = mem_1356_sv2v_reg;
  assign mem[1355] = mem_1355_sv2v_reg;
  assign mem[1354] = mem_1354_sv2v_reg;
  assign mem[1353] = mem_1353_sv2v_reg;
  assign mem[1352] = mem_1352_sv2v_reg;
  assign mem[1351] = mem_1351_sv2v_reg;
  assign mem[1350] = mem_1350_sv2v_reg;
  assign mem[1349] = mem_1349_sv2v_reg;
  assign mem[1348] = mem_1348_sv2v_reg;
  assign mem[1347] = mem_1347_sv2v_reg;
  assign mem[1346] = mem_1346_sv2v_reg;
  assign mem[1345] = mem_1345_sv2v_reg;
  assign mem[1344] = mem_1344_sv2v_reg;
  assign mem[1343] = mem_1343_sv2v_reg;
  assign mem[1342] = mem_1342_sv2v_reg;
  assign mem[1341] = mem_1341_sv2v_reg;
  assign mem[1340] = mem_1340_sv2v_reg;
  assign mem[1339] = mem_1339_sv2v_reg;
  assign mem[1338] = mem_1338_sv2v_reg;
  assign mem[1337] = mem_1337_sv2v_reg;
  assign mem[1336] = mem_1336_sv2v_reg;
  assign mem[1335] = mem_1335_sv2v_reg;
  assign mem[1334] = mem_1334_sv2v_reg;
  assign mem[1333] = mem_1333_sv2v_reg;
  assign mem[1332] = mem_1332_sv2v_reg;
  assign mem[1331] = mem_1331_sv2v_reg;
  assign mem[1330] = mem_1330_sv2v_reg;
  assign mem[1329] = mem_1329_sv2v_reg;
  assign mem[1328] = mem_1328_sv2v_reg;
  assign mem[1327] = mem_1327_sv2v_reg;
  assign mem[1326] = mem_1326_sv2v_reg;
  assign mem[1325] = mem_1325_sv2v_reg;
  assign mem[1324] = mem_1324_sv2v_reg;
  assign mem[1323] = mem_1323_sv2v_reg;
  assign mem[1322] = mem_1322_sv2v_reg;
  assign mem[1321] = mem_1321_sv2v_reg;
  assign mem[1320] = mem_1320_sv2v_reg;
  assign mem[1319] = mem_1319_sv2v_reg;
  assign mem[1318] = mem_1318_sv2v_reg;
  assign mem[1317] = mem_1317_sv2v_reg;
  assign mem[1316] = mem_1316_sv2v_reg;
  assign mem[1315] = mem_1315_sv2v_reg;
  assign mem[1314] = mem_1314_sv2v_reg;
  assign mem[1313] = mem_1313_sv2v_reg;
  assign mem[1312] = mem_1312_sv2v_reg;
  assign mem[1311] = mem_1311_sv2v_reg;
  assign mem[1310] = mem_1310_sv2v_reg;
  assign mem[1309] = mem_1309_sv2v_reg;
  assign mem[1308] = mem_1308_sv2v_reg;
  assign mem[1307] = mem_1307_sv2v_reg;
  assign mem[1306] = mem_1306_sv2v_reg;
  assign mem[1305] = mem_1305_sv2v_reg;
  assign mem[1304] = mem_1304_sv2v_reg;
  assign mem[1303] = mem_1303_sv2v_reg;
  assign mem[1302] = mem_1302_sv2v_reg;
  assign mem[1301] = mem_1301_sv2v_reg;
  assign mem[1300] = mem_1300_sv2v_reg;
  assign mem[1299] = mem_1299_sv2v_reg;
  assign mem[1298] = mem_1298_sv2v_reg;
  assign mem[1297] = mem_1297_sv2v_reg;
  assign mem[1296] = mem_1296_sv2v_reg;
  assign mem[1295] = mem_1295_sv2v_reg;
  assign mem[1294] = mem_1294_sv2v_reg;
  assign mem[1293] = mem_1293_sv2v_reg;
  assign mem[1292] = mem_1292_sv2v_reg;
  assign mem[1291] = mem_1291_sv2v_reg;
  assign mem[1290] = mem_1290_sv2v_reg;
  assign mem[1289] = mem_1289_sv2v_reg;
  assign mem[1288] = mem_1288_sv2v_reg;
  assign mem[1287] = mem_1287_sv2v_reg;
  assign mem[1286] = mem_1286_sv2v_reg;
  assign mem[1285] = mem_1285_sv2v_reg;
  assign mem[1284] = mem_1284_sv2v_reg;
  assign mem[1283] = mem_1283_sv2v_reg;
  assign mem[1282] = mem_1282_sv2v_reg;
  assign mem[1281] = mem_1281_sv2v_reg;
  assign mem[1280] = mem_1280_sv2v_reg;
  assign mem[1279] = mem_1279_sv2v_reg;
  assign mem[1278] = mem_1278_sv2v_reg;
  assign mem[1277] = mem_1277_sv2v_reg;
  assign mem[1276] = mem_1276_sv2v_reg;
  assign mem[1275] = mem_1275_sv2v_reg;
  assign mem[1274] = mem_1274_sv2v_reg;
  assign mem[1273] = mem_1273_sv2v_reg;
  assign mem[1272] = mem_1272_sv2v_reg;
  assign mem[1271] = mem_1271_sv2v_reg;
  assign mem[1270] = mem_1270_sv2v_reg;
  assign mem[1269] = mem_1269_sv2v_reg;
  assign mem[1268] = mem_1268_sv2v_reg;
  assign mem[1267] = mem_1267_sv2v_reg;
  assign mem[1266] = mem_1266_sv2v_reg;
  assign mem[1265] = mem_1265_sv2v_reg;
  assign mem[1264] = mem_1264_sv2v_reg;
  assign mem[1263] = mem_1263_sv2v_reg;
  assign mem[1262] = mem_1262_sv2v_reg;
  assign mem[1261] = mem_1261_sv2v_reg;
  assign mem[1260] = mem_1260_sv2v_reg;
  assign mem[1259] = mem_1259_sv2v_reg;
  assign mem[1258] = mem_1258_sv2v_reg;
  assign mem[1257] = mem_1257_sv2v_reg;
  assign mem[1256] = mem_1256_sv2v_reg;
  assign mem[1255] = mem_1255_sv2v_reg;
  assign mem[1254] = mem_1254_sv2v_reg;
  assign mem[1253] = mem_1253_sv2v_reg;
  assign mem[1252] = mem_1252_sv2v_reg;
  assign mem[1251] = mem_1251_sv2v_reg;
  assign mem[1250] = mem_1250_sv2v_reg;
  assign mem[1249] = mem_1249_sv2v_reg;
  assign mem[1248] = mem_1248_sv2v_reg;
  assign mem[1247] = mem_1247_sv2v_reg;
  assign mem[1246] = mem_1246_sv2v_reg;
  assign mem[1245] = mem_1245_sv2v_reg;
  assign mem[1244] = mem_1244_sv2v_reg;
  assign mem[1243] = mem_1243_sv2v_reg;
  assign mem[1242] = mem_1242_sv2v_reg;
  assign mem[1241] = mem_1241_sv2v_reg;
  assign mem[1240] = mem_1240_sv2v_reg;
  assign mem[1239] = mem_1239_sv2v_reg;
  assign mem[1238] = mem_1238_sv2v_reg;
  assign mem[1237] = mem_1237_sv2v_reg;
  assign mem[1236] = mem_1236_sv2v_reg;
  assign mem[1235] = mem_1235_sv2v_reg;
  assign mem[1234] = mem_1234_sv2v_reg;
  assign mem[1233] = mem_1233_sv2v_reg;
  assign mem[1232] = mem_1232_sv2v_reg;
  assign mem[1231] = mem_1231_sv2v_reg;
  assign mem[1230] = mem_1230_sv2v_reg;
  assign mem[1229] = mem_1229_sv2v_reg;
  assign mem[1228] = mem_1228_sv2v_reg;
  assign mem[1227] = mem_1227_sv2v_reg;
  assign mem[1226] = mem_1226_sv2v_reg;
  assign mem[1225] = mem_1225_sv2v_reg;
  assign mem[1224] = mem_1224_sv2v_reg;
  assign mem[1223] = mem_1223_sv2v_reg;
  assign mem[1222] = mem_1222_sv2v_reg;
  assign mem[1221] = mem_1221_sv2v_reg;
  assign mem[1220] = mem_1220_sv2v_reg;
  assign mem[1219] = mem_1219_sv2v_reg;
  assign mem[1218] = mem_1218_sv2v_reg;
  assign mem[1217] = mem_1217_sv2v_reg;
  assign mem[1216] = mem_1216_sv2v_reg;
  assign mem[1215] = mem_1215_sv2v_reg;
  assign mem[1214] = mem_1214_sv2v_reg;
  assign mem[1213] = mem_1213_sv2v_reg;
  assign mem[1212] = mem_1212_sv2v_reg;
  assign mem[1211] = mem_1211_sv2v_reg;
  assign mem[1210] = mem_1210_sv2v_reg;
  assign mem[1209] = mem_1209_sv2v_reg;
  assign mem[1208] = mem_1208_sv2v_reg;
  assign mem[1207] = mem_1207_sv2v_reg;
  assign mem[1206] = mem_1206_sv2v_reg;
  assign mem[1205] = mem_1205_sv2v_reg;
  assign mem[1204] = mem_1204_sv2v_reg;
  assign mem[1203] = mem_1203_sv2v_reg;
  assign mem[1202] = mem_1202_sv2v_reg;
  assign mem[1201] = mem_1201_sv2v_reg;
  assign mem[1200] = mem_1200_sv2v_reg;
  assign mem[1199] = mem_1199_sv2v_reg;
  assign mem[1198] = mem_1198_sv2v_reg;
  assign mem[1197] = mem_1197_sv2v_reg;
  assign mem[1196] = mem_1196_sv2v_reg;
  assign mem[1195] = mem_1195_sv2v_reg;
  assign mem[1194] = mem_1194_sv2v_reg;
  assign mem[1193] = mem_1193_sv2v_reg;
  assign mem[1192] = mem_1192_sv2v_reg;
  assign mem[1191] = mem_1191_sv2v_reg;
  assign mem[1190] = mem_1190_sv2v_reg;
  assign mem[1189] = mem_1189_sv2v_reg;
  assign mem[1188] = mem_1188_sv2v_reg;
  assign mem[1187] = mem_1187_sv2v_reg;
  assign mem[1186] = mem_1186_sv2v_reg;
  assign mem[1185] = mem_1185_sv2v_reg;
  assign mem[1184] = mem_1184_sv2v_reg;
  assign mem[1183] = mem_1183_sv2v_reg;
  assign mem[1182] = mem_1182_sv2v_reg;
  assign mem[1181] = mem_1181_sv2v_reg;
  assign mem[1180] = mem_1180_sv2v_reg;
  assign mem[1179] = mem_1179_sv2v_reg;
  assign mem[1178] = mem_1178_sv2v_reg;
  assign mem[1177] = mem_1177_sv2v_reg;
  assign mem[1176] = mem_1176_sv2v_reg;
  assign mem[1175] = mem_1175_sv2v_reg;
  assign mem[1174] = mem_1174_sv2v_reg;
  assign mem[1173] = mem_1173_sv2v_reg;
  assign mem[1172] = mem_1172_sv2v_reg;
  assign mem[1171] = mem_1171_sv2v_reg;
  assign mem[1170] = mem_1170_sv2v_reg;
  assign mem[1169] = mem_1169_sv2v_reg;
  assign mem[1168] = mem_1168_sv2v_reg;
  assign mem[1167] = mem_1167_sv2v_reg;
  assign mem[1166] = mem_1166_sv2v_reg;
  assign mem[1165] = mem_1165_sv2v_reg;
  assign mem[1164] = mem_1164_sv2v_reg;
  assign mem[1163] = mem_1163_sv2v_reg;
  assign mem[1162] = mem_1162_sv2v_reg;
  assign mem[1161] = mem_1161_sv2v_reg;
  assign mem[1160] = mem_1160_sv2v_reg;
  assign mem[1159] = mem_1159_sv2v_reg;
  assign mem[1158] = mem_1158_sv2v_reg;
  assign mem[1157] = mem_1157_sv2v_reg;
  assign mem[1156] = mem_1156_sv2v_reg;
  assign mem[1155] = mem_1155_sv2v_reg;
  assign mem[1154] = mem_1154_sv2v_reg;
  assign mem[1153] = mem_1153_sv2v_reg;
  assign mem[1152] = mem_1152_sv2v_reg;
  assign mem[1151] = mem_1151_sv2v_reg;
  assign mem[1150] = mem_1150_sv2v_reg;
  assign mem[1149] = mem_1149_sv2v_reg;
  assign mem[1148] = mem_1148_sv2v_reg;
  assign mem[1147] = mem_1147_sv2v_reg;
  assign mem[1146] = mem_1146_sv2v_reg;
  assign mem[1145] = mem_1145_sv2v_reg;
  assign mem[1144] = mem_1144_sv2v_reg;
  assign mem[1143] = mem_1143_sv2v_reg;
  assign mem[1142] = mem_1142_sv2v_reg;
  assign mem[1141] = mem_1141_sv2v_reg;
  assign mem[1140] = mem_1140_sv2v_reg;
  assign mem[1139] = mem_1139_sv2v_reg;
  assign mem[1138] = mem_1138_sv2v_reg;
  assign mem[1137] = mem_1137_sv2v_reg;
  assign mem[1136] = mem_1136_sv2v_reg;
  assign mem[1135] = mem_1135_sv2v_reg;
  assign mem[1134] = mem_1134_sv2v_reg;
  assign mem[1133] = mem_1133_sv2v_reg;
  assign mem[1132] = mem_1132_sv2v_reg;
  assign mem[1131] = mem_1131_sv2v_reg;
  assign mem[1130] = mem_1130_sv2v_reg;
  assign mem[1129] = mem_1129_sv2v_reg;
  assign mem[1128] = mem_1128_sv2v_reg;
  assign mem[1127] = mem_1127_sv2v_reg;
  assign mem[1126] = mem_1126_sv2v_reg;
  assign mem[1125] = mem_1125_sv2v_reg;
  assign mem[1124] = mem_1124_sv2v_reg;
  assign mem[1123] = mem_1123_sv2v_reg;
  assign mem[1122] = mem_1122_sv2v_reg;
  assign mem[1121] = mem_1121_sv2v_reg;
  assign mem[1120] = mem_1120_sv2v_reg;
  assign mem[1119] = mem_1119_sv2v_reg;
  assign mem[1118] = mem_1118_sv2v_reg;
  assign mem[1117] = mem_1117_sv2v_reg;
  assign mem[1116] = mem_1116_sv2v_reg;
  assign mem[1115] = mem_1115_sv2v_reg;
  assign mem[1114] = mem_1114_sv2v_reg;
  assign mem[1113] = mem_1113_sv2v_reg;
  assign mem[1112] = mem_1112_sv2v_reg;
  assign mem[1111] = mem_1111_sv2v_reg;
  assign mem[1110] = mem_1110_sv2v_reg;
  assign mem[1109] = mem_1109_sv2v_reg;
  assign mem[1108] = mem_1108_sv2v_reg;
  assign mem[1107] = mem_1107_sv2v_reg;
  assign mem[1106] = mem_1106_sv2v_reg;
  assign mem[1105] = mem_1105_sv2v_reg;
  assign mem[1104] = mem_1104_sv2v_reg;
  assign mem[1103] = mem_1103_sv2v_reg;
  assign mem[1102] = mem_1102_sv2v_reg;
  assign mem[1101] = mem_1101_sv2v_reg;
  assign mem[1100] = mem_1100_sv2v_reg;
  assign mem[1099] = mem_1099_sv2v_reg;
  assign mem[1098] = mem_1098_sv2v_reg;
  assign mem[1097] = mem_1097_sv2v_reg;
  assign mem[1096] = mem_1096_sv2v_reg;
  assign mem[1095] = mem_1095_sv2v_reg;
  assign mem[1094] = mem_1094_sv2v_reg;
  assign mem[1093] = mem_1093_sv2v_reg;
  assign mem[1092] = mem_1092_sv2v_reg;
  assign mem[1091] = mem_1091_sv2v_reg;
  assign mem[1090] = mem_1090_sv2v_reg;
  assign mem[1089] = mem_1089_sv2v_reg;
  assign mem[1088] = mem_1088_sv2v_reg;
  assign mem[1087] = mem_1087_sv2v_reg;
  assign mem[1086] = mem_1086_sv2v_reg;
  assign mem[1085] = mem_1085_sv2v_reg;
  assign mem[1084] = mem_1084_sv2v_reg;
  assign mem[1083] = mem_1083_sv2v_reg;
  assign mem[1082] = mem_1082_sv2v_reg;
  assign mem[1081] = mem_1081_sv2v_reg;
  assign mem[1080] = mem_1080_sv2v_reg;
  assign mem[1079] = mem_1079_sv2v_reg;
  assign mem[1078] = mem_1078_sv2v_reg;
  assign mem[1077] = mem_1077_sv2v_reg;
  assign mem[1076] = mem_1076_sv2v_reg;
  assign mem[1075] = mem_1075_sv2v_reg;
  assign mem[1074] = mem_1074_sv2v_reg;
  assign mem[1073] = mem_1073_sv2v_reg;
  assign mem[1072] = mem_1072_sv2v_reg;
  assign mem[1071] = mem_1071_sv2v_reg;
  assign mem[1070] = mem_1070_sv2v_reg;
  assign mem[1069] = mem_1069_sv2v_reg;
  assign mem[1068] = mem_1068_sv2v_reg;
  assign mem[1067] = mem_1067_sv2v_reg;
  assign mem[1066] = mem_1066_sv2v_reg;
  assign mem[1065] = mem_1065_sv2v_reg;
  assign mem[1064] = mem_1064_sv2v_reg;
  assign mem[1063] = mem_1063_sv2v_reg;
  assign mem[1062] = mem_1062_sv2v_reg;
  assign mem[1061] = mem_1061_sv2v_reg;
  assign mem[1060] = mem_1060_sv2v_reg;
  assign mem[1059] = mem_1059_sv2v_reg;
  assign mem[1058] = mem_1058_sv2v_reg;
  assign mem[1057] = mem_1057_sv2v_reg;
  assign mem[1056] = mem_1056_sv2v_reg;
  assign mem[1055] = mem_1055_sv2v_reg;
  assign mem[1054] = mem_1054_sv2v_reg;
  assign mem[1053] = mem_1053_sv2v_reg;
  assign mem[1052] = mem_1052_sv2v_reg;
  assign mem[1051] = mem_1051_sv2v_reg;
  assign mem[1050] = mem_1050_sv2v_reg;
  assign mem[1049] = mem_1049_sv2v_reg;
  assign mem[1048] = mem_1048_sv2v_reg;
  assign mem[1047] = mem_1047_sv2v_reg;
  assign mem[1046] = mem_1046_sv2v_reg;
  assign mem[1045] = mem_1045_sv2v_reg;
  assign mem[1044] = mem_1044_sv2v_reg;
  assign mem[1043] = mem_1043_sv2v_reg;
  assign mem[1042] = mem_1042_sv2v_reg;
  assign mem[1041] = mem_1041_sv2v_reg;
  assign mem[1040] = mem_1040_sv2v_reg;
  assign mem[1039] = mem_1039_sv2v_reg;
  assign mem[1038] = mem_1038_sv2v_reg;
  assign mem[1037] = mem_1037_sv2v_reg;
  assign mem[1036] = mem_1036_sv2v_reg;
  assign mem[1035] = mem_1035_sv2v_reg;
  assign mem[1034] = mem_1034_sv2v_reg;
  assign mem[1033] = mem_1033_sv2v_reg;
  assign mem[1032] = mem_1032_sv2v_reg;
  assign mem[1031] = mem_1031_sv2v_reg;
  assign mem[1030] = mem_1030_sv2v_reg;
  assign mem[1029] = mem_1029_sv2v_reg;
  assign mem[1028] = mem_1028_sv2v_reg;
  assign mem[1027] = mem_1027_sv2v_reg;
  assign mem[1026] = mem_1026_sv2v_reg;
  assign mem[1025] = mem_1025_sv2v_reg;
  assign mem[1024] = mem_1024_sv2v_reg;
  assign mem[1023] = mem_1023_sv2v_reg;
  assign mem[1022] = mem_1022_sv2v_reg;
  assign mem[1021] = mem_1021_sv2v_reg;
  assign mem[1020] = mem_1020_sv2v_reg;
  assign mem[1019] = mem_1019_sv2v_reg;
  assign mem[1018] = mem_1018_sv2v_reg;
  assign mem[1017] = mem_1017_sv2v_reg;
  assign mem[1016] = mem_1016_sv2v_reg;
  assign mem[1015] = mem_1015_sv2v_reg;
  assign mem[1014] = mem_1014_sv2v_reg;
  assign mem[1013] = mem_1013_sv2v_reg;
  assign mem[1012] = mem_1012_sv2v_reg;
  assign mem[1011] = mem_1011_sv2v_reg;
  assign mem[1010] = mem_1010_sv2v_reg;
  assign mem[1009] = mem_1009_sv2v_reg;
  assign mem[1008] = mem_1008_sv2v_reg;
  assign mem[1007] = mem_1007_sv2v_reg;
  assign mem[1006] = mem_1006_sv2v_reg;
  assign mem[1005] = mem_1005_sv2v_reg;
  assign mem[1004] = mem_1004_sv2v_reg;
  assign mem[1003] = mem_1003_sv2v_reg;
  assign mem[1002] = mem_1002_sv2v_reg;
  assign mem[1001] = mem_1001_sv2v_reg;
  assign mem[1000] = mem_1000_sv2v_reg;
  assign mem[999] = mem_999_sv2v_reg;
  assign mem[998] = mem_998_sv2v_reg;
  assign mem[997] = mem_997_sv2v_reg;
  assign mem[996] = mem_996_sv2v_reg;
  assign mem[995] = mem_995_sv2v_reg;
  assign mem[994] = mem_994_sv2v_reg;
  assign mem[993] = mem_993_sv2v_reg;
  assign mem[992] = mem_992_sv2v_reg;
  assign mem[991] = mem_991_sv2v_reg;
  assign mem[990] = mem_990_sv2v_reg;
  assign mem[989] = mem_989_sv2v_reg;
  assign mem[988] = mem_988_sv2v_reg;
  assign mem[987] = mem_987_sv2v_reg;
  assign mem[986] = mem_986_sv2v_reg;
  assign mem[985] = mem_985_sv2v_reg;
  assign mem[984] = mem_984_sv2v_reg;
  assign mem[983] = mem_983_sv2v_reg;
  assign mem[982] = mem_982_sv2v_reg;
  assign mem[981] = mem_981_sv2v_reg;
  assign mem[980] = mem_980_sv2v_reg;
  assign mem[979] = mem_979_sv2v_reg;
  assign mem[978] = mem_978_sv2v_reg;
  assign mem[977] = mem_977_sv2v_reg;
  assign mem[976] = mem_976_sv2v_reg;
  assign mem[975] = mem_975_sv2v_reg;
  assign mem[974] = mem_974_sv2v_reg;
  assign mem[973] = mem_973_sv2v_reg;
  assign mem[972] = mem_972_sv2v_reg;
  assign mem[971] = mem_971_sv2v_reg;
  assign mem[970] = mem_970_sv2v_reg;
  assign mem[969] = mem_969_sv2v_reg;
  assign mem[968] = mem_968_sv2v_reg;
  assign mem[967] = mem_967_sv2v_reg;
  assign mem[966] = mem_966_sv2v_reg;
  assign mem[965] = mem_965_sv2v_reg;
  assign mem[964] = mem_964_sv2v_reg;
  assign mem[963] = mem_963_sv2v_reg;
  assign mem[962] = mem_962_sv2v_reg;
  assign mem[961] = mem_961_sv2v_reg;
  assign mem[960] = mem_960_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[61] = (N76)? mem[61] : 
                        (N78)? mem[123] : 
                        (N80)? mem[185] : 
                        (N82)? mem[247] : 
                        (N84)? mem[309] : 
                        (N86)? mem[371] : 
                        (N88)? mem[433] : 
                        (N90)? mem[495] : 
                        (N92)? mem[557] : 
                        (N94)? mem[619] : 
                        (N96)? mem[681] : 
                        (N98)? mem[743] : 
                        (N100)? mem[805] : 
                        (N102)? mem[867] : 
                        (N104)? mem[929] : 
                        (N106)? mem[991] : 
                        (N108)? mem[1053] : 
                        (N110)? mem[1115] : 
                        (N112)? mem[1177] : 
                        (N114)? mem[1239] : 
                        (N116)? mem[1301] : 
                        (N118)? mem[1363] : 
                        (N120)? mem[1425] : 
                        (N122)? mem[1487] : 
                        (N124)? mem[1549] : 
                        (N126)? mem[1611] : 
                        (N128)? mem[1673] : 
                        (N130)? mem[1735] : 
                        (N132)? mem[1797] : 
                        (N134)? mem[1859] : 
                        (N136)? mem[1921] : 
                        (N138)? mem[1983] : 
                        (N77)? mem[2045] : 
                        (N79)? mem[2107] : 
                        (N81)? mem[2169] : 
                        (N83)? mem[2231] : 
                        (N85)? mem[2293] : 
                        (N87)? mem[2355] : 
                        (N89)? mem[2417] : 
                        (N91)? mem[2479] : 
                        (N93)? mem[2541] : 
                        (N95)? mem[2603] : 
                        (N97)? mem[2665] : 
                        (N99)? mem[2727] : 
                        (N101)? mem[2789] : 
                        (N103)? mem[2851] : 
                        (N105)? mem[2913] : 
                        (N107)? mem[2975] : 
                        (N109)? mem[3037] : 
                        (N111)? mem[3099] : 
                        (N113)? mem[3161] : 
                        (N115)? mem[3223] : 
                        (N117)? mem[3285] : 
                        (N119)? mem[3347] : 
                        (N121)? mem[3409] : 
                        (N123)? mem[3471] : 
                        (N125)? mem[3533] : 
                        (N127)? mem[3595] : 
                        (N129)? mem[3657] : 
                        (N131)? mem[3719] : 
                        (N133)? mem[3781] : 
                        (N135)? mem[3843] : 
                        (N137)? mem[3905] : 
                        (N139)? mem[3967] : 1'b0;
  assign r_data_o[60] = (N76)? mem[60] : 
                        (N78)? mem[122] : 
                        (N80)? mem[184] : 
                        (N82)? mem[246] : 
                        (N84)? mem[308] : 
                        (N86)? mem[370] : 
                        (N88)? mem[432] : 
                        (N90)? mem[494] : 
                        (N92)? mem[556] : 
                        (N94)? mem[618] : 
                        (N96)? mem[680] : 
                        (N98)? mem[742] : 
                        (N100)? mem[804] : 
                        (N102)? mem[866] : 
                        (N104)? mem[928] : 
                        (N106)? mem[990] : 
                        (N108)? mem[1052] : 
                        (N110)? mem[1114] : 
                        (N112)? mem[1176] : 
                        (N114)? mem[1238] : 
                        (N116)? mem[1300] : 
                        (N118)? mem[1362] : 
                        (N120)? mem[1424] : 
                        (N122)? mem[1486] : 
                        (N124)? mem[1548] : 
                        (N126)? mem[1610] : 
                        (N128)? mem[1672] : 
                        (N130)? mem[1734] : 
                        (N132)? mem[1796] : 
                        (N134)? mem[1858] : 
                        (N136)? mem[1920] : 
                        (N138)? mem[1982] : 
                        (N77)? mem[2044] : 
                        (N79)? mem[2106] : 
                        (N81)? mem[2168] : 
                        (N83)? mem[2230] : 
                        (N85)? mem[2292] : 
                        (N87)? mem[2354] : 
                        (N89)? mem[2416] : 
                        (N91)? mem[2478] : 
                        (N93)? mem[2540] : 
                        (N95)? mem[2602] : 
                        (N97)? mem[2664] : 
                        (N99)? mem[2726] : 
                        (N101)? mem[2788] : 
                        (N103)? mem[2850] : 
                        (N105)? mem[2912] : 
                        (N107)? mem[2974] : 
                        (N109)? mem[3036] : 
                        (N111)? mem[3098] : 
                        (N113)? mem[3160] : 
                        (N115)? mem[3222] : 
                        (N117)? mem[3284] : 
                        (N119)? mem[3346] : 
                        (N121)? mem[3408] : 
                        (N123)? mem[3470] : 
                        (N125)? mem[3532] : 
                        (N127)? mem[3594] : 
                        (N129)? mem[3656] : 
                        (N131)? mem[3718] : 
                        (N133)? mem[3780] : 
                        (N135)? mem[3842] : 
                        (N137)? mem[3904] : 
                        (N139)? mem[3966] : 1'b0;
  assign r_data_o[59] = (N76)? mem[59] : 
                        (N78)? mem[121] : 
                        (N80)? mem[183] : 
                        (N82)? mem[245] : 
                        (N84)? mem[307] : 
                        (N86)? mem[369] : 
                        (N88)? mem[431] : 
                        (N90)? mem[493] : 
                        (N92)? mem[555] : 
                        (N94)? mem[617] : 
                        (N96)? mem[679] : 
                        (N98)? mem[741] : 
                        (N100)? mem[803] : 
                        (N102)? mem[865] : 
                        (N104)? mem[927] : 
                        (N106)? mem[989] : 
                        (N108)? mem[1051] : 
                        (N110)? mem[1113] : 
                        (N112)? mem[1175] : 
                        (N114)? mem[1237] : 
                        (N116)? mem[1299] : 
                        (N118)? mem[1361] : 
                        (N120)? mem[1423] : 
                        (N122)? mem[1485] : 
                        (N124)? mem[1547] : 
                        (N126)? mem[1609] : 
                        (N128)? mem[1671] : 
                        (N130)? mem[1733] : 
                        (N132)? mem[1795] : 
                        (N134)? mem[1857] : 
                        (N136)? mem[1919] : 
                        (N138)? mem[1981] : 
                        (N77)? mem[2043] : 
                        (N79)? mem[2105] : 
                        (N81)? mem[2167] : 
                        (N83)? mem[2229] : 
                        (N85)? mem[2291] : 
                        (N87)? mem[2353] : 
                        (N89)? mem[2415] : 
                        (N91)? mem[2477] : 
                        (N93)? mem[2539] : 
                        (N95)? mem[2601] : 
                        (N97)? mem[2663] : 
                        (N99)? mem[2725] : 
                        (N101)? mem[2787] : 
                        (N103)? mem[2849] : 
                        (N105)? mem[2911] : 
                        (N107)? mem[2973] : 
                        (N109)? mem[3035] : 
                        (N111)? mem[3097] : 
                        (N113)? mem[3159] : 
                        (N115)? mem[3221] : 
                        (N117)? mem[3283] : 
                        (N119)? mem[3345] : 
                        (N121)? mem[3407] : 
                        (N123)? mem[3469] : 
                        (N125)? mem[3531] : 
                        (N127)? mem[3593] : 
                        (N129)? mem[3655] : 
                        (N131)? mem[3717] : 
                        (N133)? mem[3779] : 
                        (N135)? mem[3841] : 
                        (N137)? mem[3903] : 
                        (N139)? mem[3965] : 1'b0;
  assign r_data_o[58] = (N76)? mem[58] : 
                        (N78)? mem[120] : 
                        (N80)? mem[182] : 
                        (N82)? mem[244] : 
                        (N84)? mem[306] : 
                        (N86)? mem[368] : 
                        (N88)? mem[430] : 
                        (N90)? mem[492] : 
                        (N92)? mem[554] : 
                        (N94)? mem[616] : 
                        (N96)? mem[678] : 
                        (N98)? mem[740] : 
                        (N100)? mem[802] : 
                        (N102)? mem[864] : 
                        (N104)? mem[926] : 
                        (N106)? mem[988] : 
                        (N108)? mem[1050] : 
                        (N110)? mem[1112] : 
                        (N112)? mem[1174] : 
                        (N114)? mem[1236] : 
                        (N116)? mem[1298] : 
                        (N118)? mem[1360] : 
                        (N120)? mem[1422] : 
                        (N122)? mem[1484] : 
                        (N124)? mem[1546] : 
                        (N126)? mem[1608] : 
                        (N128)? mem[1670] : 
                        (N130)? mem[1732] : 
                        (N132)? mem[1794] : 
                        (N134)? mem[1856] : 
                        (N136)? mem[1918] : 
                        (N138)? mem[1980] : 
                        (N77)? mem[2042] : 
                        (N79)? mem[2104] : 
                        (N81)? mem[2166] : 
                        (N83)? mem[2228] : 
                        (N85)? mem[2290] : 
                        (N87)? mem[2352] : 
                        (N89)? mem[2414] : 
                        (N91)? mem[2476] : 
                        (N93)? mem[2538] : 
                        (N95)? mem[2600] : 
                        (N97)? mem[2662] : 
                        (N99)? mem[2724] : 
                        (N101)? mem[2786] : 
                        (N103)? mem[2848] : 
                        (N105)? mem[2910] : 
                        (N107)? mem[2972] : 
                        (N109)? mem[3034] : 
                        (N111)? mem[3096] : 
                        (N113)? mem[3158] : 
                        (N115)? mem[3220] : 
                        (N117)? mem[3282] : 
                        (N119)? mem[3344] : 
                        (N121)? mem[3406] : 
                        (N123)? mem[3468] : 
                        (N125)? mem[3530] : 
                        (N127)? mem[3592] : 
                        (N129)? mem[3654] : 
                        (N131)? mem[3716] : 
                        (N133)? mem[3778] : 
                        (N135)? mem[3840] : 
                        (N137)? mem[3902] : 
                        (N139)? mem[3964] : 1'b0;
  assign r_data_o[57] = (N76)? mem[57] : 
                        (N78)? mem[119] : 
                        (N80)? mem[181] : 
                        (N82)? mem[243] : 
                        (N84)? mem[305] : 
                        (N86)? mem[367] : 
                        (N88)? mem[429] : 
                        (N90)? mem[491] : 
                        (N92)? mem[553] : 
                        (N94)? mem[615] : 
                        (N96)? mem[677] : 
                        (N98)? mem[739] : 
                        (N100)? mem[801] : 
                        (N102)? mem[863] : 
                        (N104)? mem[925] : 
                        (N106)? mem[987] : 
                        (N108)? mem[1049] : 
                        (N110)? mem[1111] : 
                        (N112)? mem[1173] : 
                        (N114)? mem[1235] : 
                        (N116)? mem[1297] : 
                        (N118)? mem[1359] : 
                        (N120)? mem[1421] : 
                        (N122)? mem[1483] : 
                        (N124)? mem[1545] : 
                        (N126)? mem[1607] : 
                        (N128)? mem[1669] : 
                        (N130)? mem[1731] : 
                        (N132)? mem[1793] : 
                        (N134)? mem[1855] : 
                        (N136)? mem[1917] : 
                        (N138)? mem[1979] : 
                        (N77)? mem[2041] : 
                        (N79)? mem[2103] : 
                        (N81)? mem[2165] : 
                        (N83)? mem[2227] : 
                        (N85)? mem[2289] : 
                        (N87)? mem[2351] : 
                        (N89)? mem[2413] : 
                        (N91)? mem[2475] : 
                        (N93)? mem[2537] : 
                        (N95)? mem[2599] : 
                        (N97)? mem[2661] : 
                        (N99)? mem[2723] : 
                        (N101)? mem[2785] : 
                        (N103)? mem[2847] : 
                        (N105)? mem[2909] : 
                        (N107)? mem[2971] : 
                        (N109)? mem[3033] : 
                        (N111)? mem[3095] : 
                        (N113)? mem[3157] : 
                        (N115)? mem[3219] : 
                        (N117)? mem[3281] : 
                        (N119)? mem[3343] : 
                        (N121)? mem[3405] : 
                        (N123)? mem[3467] : 
                        (N125)? mem[3529] : 
                        (N127)? mem[3591] : 
                        (N129)? mem[3653] : 
                        (N131)? mem[3715] : 
                        (N133)? mem[3777] : 
                        (N135)? mem[3839] : 
                        (N137)? mem[3901] : 
                        (N139)? mem[3963] : 1'b0;
  assign r_data_o[56] = (N76)? mem[56] : 
                        (N78)? mem[118] : 
                        (N80)? mem[180] : 
                        (N82)? mem[242] : 
                        (N84)? mem[304] : 
                        (N86)? mem[366] : 
                        (N88)? mem[428] : 
                        (N90)? mem[490] : 
                        (N92)? mem[552] : 
                        (N94)? mem[614] : 
                        (N96)? mem[676] : 
                        (N98)? mem[738] : 
                        (N100)? mem[800] : 
                        (N102)? mem[862] : 
                        (N104)? mem[924] : 
                        (N106)? mem[986] : 
                        (N108)? mem[1048] : 
                        (N110)? mem[1110] : 
                        (N112)? mem[1172] : 
                        (N114)? mem[1234] : 
                        (N116)? mem[1296] : 
                        (N118)? mem[1358] : 
                        (N120)? mem[1420] : 
                        (N122)? mem[1482] : 
                        (N124)? mem[1544] : 
                        (N126)? mem[1606] : 
                        (N128)? mem[1668] : 
                        (N130)? mem[1730] : 
                        (N132)? mem[1792] : 
                        (N134)? mem[1854] : 
                        (N136)? mem[1916] : 
                        (N138)? mem[1978] : 
                        (N77)? mem[2040] : 
                        (N79)? mem[2102] : 
                        (N81)? mem[2164] : 
                        (N83)? mem[2226] : 
                        (N85)? mem[2288] : 
                        (N87)? mem[2350] : 
                        (N89)? mem[2412] : 
                        (N91)? mem[2474] : 
                        (N93)? mem[2536] : 
                        (N95)? mem[2598] : 
                        (N97)? mem[2660] : 
                        (N99)? mem[2722] : 
                        (N101)? mem[2784] : 
                        (N103)? mem[2846] : 
                        (N105)? mem[2908] : 
                        (N107)? mem[2970] : 
                        (N109)? mem[3032] : 
                        (N111)? mem[3094] : 
                        (N113)? mem[3156] : 
                        (N115)? mem[3218] : 
                        (N117)? mem[3280] : 
                        (N119)? mem[3342] : 
                        (N121)? mem[3404] : 
                        (N123)? mem[3466] : 
                        (N125)? mem[3528] : 
                        (N127)? mem[3590] : 
                        (N129)? mem[3652] : 
                        (N131)? mem[3714] : 
                        (N133)? mem[3776] : 
                        (N135)? mem[3838] : 
                        (N137)? mem[3900] : 
                        (N139)? mem[3962] : 1'b0;
  assign r_data_o[55] = (N76)? mem[55] : 
                        (N78)? mem[117] : 
                        (N80)? mem[179] : 
                        (N82)? mem[241] : 
                        (N84)? mem[303] : 
                        (N86)? mem[365] : 
                        (N88)? mem[427] : 
                        (N90)? mem[489] : 
                        (N92)? mem[551] : 
                        (N94)? mem[613] : 
                        (N96)? mem[675] : 
                        (N98)? mem[737] : 
                        (N100)? mem[799] : 
                        (N102)? mem[861] : 
                        (N104)? mem[923] : 
                        (N106)? mem[985] : 
                        (N108)? mem[1047] : 
                        (N110)? mem[1109] : 
                        (N112)? mem[1171] : 
                        (N114)? mem[1233] : 
                        (N116)? mem[1295] : 
                        (N118)? mem[1357] : 
                        (N120)? mem[1419] : 
                        (N122)? mem[1481] : 
                        (N124)? mem[1543] : 
                        (N126)? mem[1605] : 
                        (N128)? mem[1667] : 
                        (N130)? mem[1729] : 
                        (N132)? mem[1791] : 
                        (N134)? mem[1853] : 
                        (N136)? mem[1915] : 
                        (N138)? mem[1977] : 
                        (N77)? mem[2039] : 
                        (N79)? mem[2101] : 
                        (N81)? mem[2163] : 
                        (N83)? mem[2225] : 
                        (N85)? mem[2287] : 
                        (N87)? mem[2349] : 
                        (N89)? mem[2411] : 
                        (N91)? mem[2473] : 
                        (N93)? mem[2535] : 
                        (N95)? mem[2597] : 
                        (N97)? mem[2659] : 
                        (N99)? mem[2721] : 
                        (N101)? mem[2783] : 
                        (N103)? mem[2845] : 
                        (N105)? mem[2907] : 
                        (N107)? mem[2969] : 
                        (N109)? mem[3031] : 
                        (N111)? mem[3093] : 
                        (N113)? mem[3155] : 
                        (N115)? mem[3217] : 
                        (N117)? mem[3279] : 
                        (N119)? mem[3341] : 
                        (N121)? mem[3403] : 
                        (N123)? mem[3465] : 
                        (N125)? mem[3527] : 
                        (N127)? mem[3589] : 
                        (N129)? mem[3651] : 
                        (N131)? mem[3713] : 
                        (N133)? mem[3775] : 
                        (N135)? mem[3837] : 
                        (N137)? mem[3899] : 
                        (N139)? mem[3961] : 1'b0;
  assign r_data_o[54] = (N76)? mem[54] : 
                        (N78)? mem[116] : 
                        (N80)? mem[178] : 
                        (N82)? mem[240] : 
                        (N84)? mem[302] : 
                        (N86)? mem[364] : 
                        (N88)? mem[426] : 
                        (N90)? mem[488] : 
                        (N92)? mem[550] : 
                        (N94)? mem[612] : 
                        (N96)? mem[674] : 
                        (N98)? mem[736] : 
                        (N100)? mem[798] : 
                        (N102)? mem[860] : 
                        (N104)? mem[922] : 
                        (N106)? mem[984] : 
                        (N108)? mem[1046] : 
                        (N110)? mem[1108] : 
                        (N112)? mem[1170] : 
                        (N114)? mem[1232] : 
                        (N116)? mem[1294] : 
                        (N118)? mem[1356] : 
                        (N120)? mem[1418] : 
                        (N122)? mem[1480] : 
                        (N124)? mem[1542] : 
                        (N126)? mem[1604] : 
                        (N128)? mem[1666] : 
                        (N130)? mem[1728] : 
                        (N132)? mem[1790] : 
                        (N134)? mem[1852] : 
                        (N136)? mem[1914] : 
                        (N138)? mem[1976] : 
                        (N77)? mem[2038] : 
                        (N79)? mem[2100] : 
                        (N81)? mem[2162] : 
                        (N83)? mem[2224] : 
                        (N85)? mem[2286] : 
                        (N87)? mem[2348] : 
                        (N89)? mem[2410] : 
                        (N91)? mem[2472] : 
                        (N93)? mem[2534] : 
                        (N95)? mem[2596] : 
                        (N97)? mem[2658] : 
                        (N99)? mem[2720] : 
                        (N101)? mem[2782] : 
                        (N103)? mem[2844] : 
                        (N105)? mem[2906] : 
                        (N107)? mem[2968] : 
                        (N109)? mem[3030] : 
                        (N111)? mem[3092] : 
                        (N113)? mem[3154] : 
                        (N115)? mem[3216] : 
                        (N117)? mem[3278] : 
                        (N119)? mem[3340] : 
                        (N121)? mem[3402] : 
                        (N123)? mem[3464] : 
                        (N125)? mem[3526] : 
                        (N127)? mem[3588] : 
                        (N129)? mem[3650] : 
                        (N131)? mem[3712] : 
                        (N133)? mem[3774] : 
                        (N135)? mem[3836] : 
                        (N137)? mem[3898] : 
                        (N139)? mem[3960] : 1'b0;
  assign r_data_o[53] = (N76)? mem[53] : 
                        (N78)? mem[115] : 
                        (N80)? mem[177] : 
                        (N82)? mem[239] : 
                        (N84)? mem[301] : 
                        (N86)? mem[363] : 
                        (N88)? mem[425] : 
                        (N90)? mem[487] : 
                        (N92)? mem[549] : 
                        (N94)? mem[611] : 
                        (N96)? mem[673] : 
                        (N98)? mem[735] : 
                        (N100)? mem[797] : 
                        (N102)? mem[859] : 
                        (N104)? mem[921] : 
                        (N106)? mem[983] : 
                        (N108)? mem[1045] : 
                        (N110)? mem[1107] : 
                        (N112)? mem[1169] : 
                        (N114)? mem[1231] : 
                        (N116)? mem[1293] : 
                        (N118)? mem[1355] : 
                        (N120)? mem[1417] : 
                        (N122)? mem[1479] : 
                        (N124)? mem[1541] : 
                        (N126)? mem[1603] : 
                        (N128)? mem[1665] : 
                        (N130)? mem[1727] : 
                        (N132)? mem[1789] : 
                        (N134)? mem[1851] : 
                        (N136)? mem[1913] : 
                        (N138)? mem[1975] : 
                        (N77)? mem[2037] : 
                        (N79)? mem[2099] : 
                        (N81)? mem[2161] : 
                        (N83)? mem[2223] : 
                        (N85)? mem[2285] : 
                        (N87)? mem[2347] : 
                        (N89)? mem[2409] : 
                        (N91)? mem[2471] : 
                        (N93)? mem[2533] : 
                        (N95)? mem[2595] : 
                        (N97)? mem[2657] : 
                        (N99)? mem[2719] : 
                        (N101)? mem[2781] : 
                        (N103)? mem[2843] : 
                        (N105)? mem[2905] : 
                        (N107)? mem[2967] : 
                        (N109)? mem[3029] : 
                        (N111)? mem[3091] : 
                        (N113)? mem[3153] : 
                        (N115)? mem[3215] : 
                        (N117)? mem[3277] : 
                        (N119)? mem[3339] : 
                        (N121)? mem[3401] : 
                        (N123)? mem[3463] : 
                        (N125)? mem[3525] : 
                        (N127)? mem[3587] : 
                        (N129)? mem[3649] : 
                        (N131)? mem[3711] : 
                        (N133)? mem[3773] : 
                        (N135)? mem[3835] : 
                        (N137)? mem[3897] : 
                        (N139)? mem[3959] : 1'b0;
  assign r_data_o[52] = (N76)? mem[52] : 
                        (N78)? mem[114] : 
                        (N80)? mem[176] : 
                        (N82)? mem[238] : 
                        (N84)? mem[300] : 
                        (N86)? mem[362] : 
                        (N88)? mem[424] : 
                        (N90)? mem[486] : 
                        (N92)? mem[548] : 
                        (N94)? mem[610] : 
                        (N96)? mem[672] : 
                        (N98)? mem[734] : 
                        (N100)? mem[796] : 
                        (N102)? mem[858] : 
                        (N104)? mem[920] : 
                        (N106)? mem[982] : 
                        (N108)? mem[1044] : 
                        (N110)? mem[1106] : 
                        (N112)? mem[1168] : 
                        (N114)? mem[1230] : 
                        (N116)? mem[1292] : 
                        (N118)? mem[1354] : 
                        (N120)? mem[1416] : 
                        (N122)? mem[1478] : 
                        (N124)? mem[1540] : 
                        (N126)? mem[1602] : 
                        (N128)? mem[1664] : 
                        (N130)? mem[1726] : 
                        (N132)? mem[1788] : 
                        (N134)? mem[1850] : 
                        (N136)? mem[1912] : 
                        (N138)? mem[1974] : 
                        (N77)? mem[2036] : 
                        (N79)? mem[2098] : 
                        (N81)? mem[2160] : 
                        (N83)? mem[2222] : 
                        (N85)? mem[2284] : 
                        (N87)? mem[2346] : 
                        (N89)? mem[2408] : 
                        (N91)? mem[2470] : 
                        (N93)? mem[2532] : 
                        (N95)? mem[2594] : 
                        (N97)? mem[2656] : 
                        (N99)? mem[2718] : 
                        (N101)? mem[2780] : 
                        (N103)? mem[2842] : 
                        (N105)? mem[2904] : 
                        (N107)? mem[2966] : 
                        (N109)? mem[3028] : 
                        (N111)? mem[3090] : 
                        (N113)? mem[3152] : 
                        (N115)? mem[3214] : 
                        (N117)? mem[3276] : 
                        (N119)? mem[3338] : 
                        (N121)? mem[3400] : 
                        (N123)? mem[3462] : 
                        (N125)? mem[3524] : 
                        (N127)? mem[3586] : 
                        (N129)? mem[3648] : 
                        (N131)? mem[3710] : 
                        (N133)? mem[3772] : 
                        (N135)? mem[3834] : 
                        (N137)? mem[3896] : 
                        (N139)? mem[3958] : 1'b0;
  assign r_data_o[51] = (N76)? mem[51] : 
                        (N78)? mem[113] : 
                        (N80)? mem[175] : 
                        (N82)? mem[237] : 
                        (N84)? mem[299] : 
                        (N86)? mem[361] : 
                        (N88)? mem[423] : 
                        (N90)? mem[485] : 
                        (N92)? mem[547] : 
                        (N94)? mem[609] : 
                        (N96)? mem[671] : 
                        (N98)? mem[733] : 
                        (N100)? mem[795] : 
                        (N102)? mem[857] : 
                        (N104)? mem[919] : 
                        (N106)? mem[981] : 
                        (N108)? mem[1043] : 
                        (N110)? mem[1105] : 
                        (N112)? mem[1167] : 
                        (N114)? mem[1229] : 
                        (N116)? mem[1291] : 
                        (N118)? mem[1353] : 
                        (N120)? mem[1415] : 
                        (N122)? mem[1477] : 
                        (N124)? mem[1539] : 
                        (N126)? mem[1601] : 
                        (N128)? mem[1663] : 
                        (N130)? mem[1725] : 
                        (N132)? mem[1787] : 
                        (N134)? mem[1849] : 
                        (N136)? mem[1911] : 
                        (N138)? mem[1973] : 
                        (N77)? mem[2035] : 
                        (N79)? mem[2097] : 
                        (N81)? mem[2159] : 
                        (N83)? mem[2221] : 
                        (N85)? mem[2283] : 
                        (N87)? mem[2345] : 
                        (N89)? mem[2407] : 
                        (N91)? mem[2469] : 
                        (N93)? mem[2531] : 
                        (N95)? mem[2593] : 
                        (N97)? mem[2655] : 
                        (N99)? mem[2717] : 
                        (N101)? mem[2779] : 
                        (N103)? mem[2841] : 
                        (N105)? mem[2903] : 
                        (N107)? mem[2965] : 
                        (N109)? mem[3027] : 
                        (N111)? mem[3089] : 
                        (N113)? mem[3151] : 
                        (N115)? mem[3213] : 
                        (N117)? mem[3275] : 
                        (N119)? mem[3337] : 
                        (N121)? mem[3399] : 
                        (N123)? mem[3461] : 
                        (N125)? mem[3523] : 
                        (N127)? mem[3585] : 
                        (N129)? mem[3647] : 
                        (N131)? mem[3709] : 
                        (N133)? mem[3771] : 
                        (N135)? mem[3833] : 
                        (N137)? mem[3895] : 
                        (N139)? mem[3957] : 1'b0;
  assign r_data_o[50] = (N76)? mem[50] : 
                        (N78)? mem[112] : 
                        (N80)? mem[174] : 
                        (N82)? mem[236] : 
                        (N84)? mem[298] : 
                        (N86)? mem[360] : 
                        (N88)? mem[422] : 
                        (N90)? mem[484] : 
                        (N92)? mem[546] : 
                        (N94)? mem[608] : 
                        (N96)? mem[670] : 
                        (N98)? mem[732] : 
                        (N100)? mem[794] : 
                        (N102)? mem[856] : 
                        (N104)? mem[918] : 
                        (N106)? mem[980] : 
                        (N108)? mem[1042] : 
                        (N110)? mem[1104] : 
                        (N112)? mem[1166] : 
                        (N114)? mem[1228] : 
                        (N116)? mem[1290] : 
                        (N118)? mem[1352] : 
                        (N120)? mem[1414] : 
                        (N122)? mem[1476] : 
                        (N124)? mem[1538] : 
                        (N126)? mem[1600] : 
                        (N128)? mem[1662] : 
                        (N130)? mem[1724] : 
                        (N132)? mem[1786] : 
                        (N134)? mem[1848] : 
                        (N136)? mem[1910] : 
                        (N138)? mem[1972] : 
                        (N77)? mem[2034] : 
                        (N79)? mem[2096] : 
                        (N81)? mem[2158] : 
                        (N83)? mem[2220] : 
                        (N85)? mem[2282] : 
                        (N87)? mem[2344] : 
                        (N89)? mem[2406] : 
                        (N91)? mem[2468] : 
                        (N93)? mem[2530] : 
                        (N95)? mem[2592] : 
                        (N97)? mem[2654] : 
                        (N99)? mem[2716] : 
                        (N101)? mem[2778] : 
                        (N103)? mem[2840] : 
                        (N105)? mem[2902] : 
                        (N107)? mem[2964] : 
                        (N109)? mem[3026] : 
                        (N111)? mem[3088] : 
                        (N113)? mem[3150] : 
                        (N115)? mem[3212] : 
                        (N117)? mem[3274] : 
                        (N119)? mem[3336] : 
                        (N121)? mem[3398] : 
                        (N123)? mem[3460] : 
                        (N125)? mem[3522] : 
                        (N127)? mem[3584] : 
                        (N129)? mem[3646] : 
                        (N131)? mem[3708] : 
                        (N133)? mem[3770] : 
                        (N135)? mem[3832] : 
                        (N137)? mem[3894] : 
                        (N139)? mem[3956] : 1'b0;
  assign r_data_o[49] = (N76)? mem[49] : 
                        (N78)? mem[111] : 
                        (N80)? mem[173] : 
                        (N82)? mem[235] : 
                        (N84)? mem[297] : 
                        (N86)? mem[359] : 
                        (N88)? mem[421] : 
                        (N90)? mem[483] : 
                        (N92)? mem[545] : 
                        (N94)? mem[607] : 
                        (N96)? mem[669] : 
                        (N98)? mem[731] : 
                        (N100)? mem[793] : 
                        (N102)? mem[855] : 
                        (N104)? mem[917] : 
                        (N106)? mem[979] : 
                        (N108)? mem[1041] : 
                        (N110)? mem[1103] : 
                        (N112)? mem[1165] : 
                        (N114)? mem[1227] : 
                        (N116)? mem[1289] : 
                        (N118)? mem[1351] : 
                        (N120)? mem[1413] : 
                        (N122)? mem[1475] : 
                        (N124)? mem[1537] : 
                        (N126)? mem[1599] : 
                        (N128)? mem[1661] : 
                        (N130)? mem[1723] : 
                        (N132)? mem[1785] : 
                        (N134)? mem[1847] : 
                        (N136)? mem[1909] : 
                        (N138)? mem[1971] : 
                        (N77)? mem[2033] : 
                        (N79)? mem[2095] : 
                        (N81)? mem[2157] : 
                        (N83)? mem[2219] : 
                        (N85)? mem[2281] : 
                        (N87)? mem[2343] : 
                        (N89)? mem[2405] : 
                        (N91)? mem[2467] : 
                        (N93)? mem[2529] : 
                        (N95)? mem[2591] : 
                        (N97)? mem[2653] : 
                        (N99)? mem[2715] : 
                        (N101)? mem[2777] : 
                        (N103)? mem[2839] : 
                        (N105)? mem[2901] : 
                        (N107)? mem[2963] : 
                        (N109)? mem[3025] : 
                        (N111)? mem[3087] : 
                        (N113)? mem[3149] : 
                        (N115)? mem[3211] : 
                        (N117)? mem[3273] : 
                        (N119)? mem[3335] : 
                        (N121)? mem[3397] : 
                        (N123)? mem[3459] : 
                        (N125)? mem[3521] : 
                        (N127)? mem[3583] : 
                        (N129)? mem[3645] : 
                        (N131)? mem[3707] : 
                        (N133)? mem[3769] : 
                        (N135)? mem[3831] : 
                        (N137)? mem[3893] : 
                        (N139)? mem[3955] : 1'b0;
  assign r_data_o[48] = (N76)? mem[48] : 
                        (N78)? mem[110] : 
                        (N80)? mem[172] : 
                        (N82)? mem[234] : 
                        (N84)? mem[296] : 
                        (N86)? mem[358] : 
                        (N88)? mem[420] : 
                        (N90)? mem[482] : 
                        (N92)? mem[544] : 
                        (N94)? mem[606] : 
                        (N96)? mem[668] : 
                        (N98)? mem[730] : 
                        (N100)? mem[792] : 
                        (N102)? mem[854] : 
                        (N104)? mem[916] : 
                        (N106)? mem[978] : 
                        (N108)? mem[1040] : 
                        (N110)? mem[1102] : 
                        (N112)? mem[1164] : 
                        (N114)? mem[1226] : 
                        (N116)? mem[1288] : 
                        (N118)? mem[1350] : 
                        (N120)? mem[1412] : 
                        (N122)? mem[1474] : 
                        (N124)? mem[1536] : 
                        (N126)? mem[1598] : 
                        (N128)? mem[1660] : 
                        (N130)? mem[1722] : 
                        (N132)? mem[1784] : 
                        (N134)? mem[1846] : 
                        (N136)? mem[1908] : 
                        (N138)? mem[1970] : 
                        (N77)? mem[2032] : 
                        (N79)? mem[2094] : 
                        (N81)? mem[2156] : 
                        (N83)? mem[2218] : 
                        (N85)? mem[2280] : 
                        (N87)? mem[2342] : 
                        (N89)? mem[2404] : 
                        (N91)? mem[2466] : 
                        (N93)? mem[2528] : 
                        (N95)? mem[2590] : 
                        (N97)? mem[2652] : 
                        (N99)? mem[2714] : 
                        (N101)? mem[2776] : 
                        (N103)? mem[2838] : 
                        (N105)? mem[2900] : 
                        (N107)? mem[2962] : 
                        (N109)? mem[3024] : 
                        (N111)? mem[3086] : 
                        (N113)? mem[3148] : 
                        (N115)? mem[3210] : 
                        (N117)? mem[3272] : 
                        (N119)? mem[3334] : 
                        (N121)? mem[3396] : 
                        (N123)? mem[3458] : 
                        (N125)? mem[3520] : 
                        (N127)? mem[3582] : 
                        (N129)? mem[3644] : 
                        (N131)? mem[3706] : 
                        (N133)? mem[3768] : 
                        (N135)? mem[3830] : 
                        (N137)? mem[3892] : 
                        (N139)? mem[3954] : 1'b0;
  assign r_data_o[47] = (N76)? mem[47] : 
                        (N78)? mem[109] : 
                        (N80)? mem[171] : 
                        (N82)? mem[233] : 
                        (N84)? mem[295] : 
                        (N86)? mem[357] : 
                        (N88)? mem[419] : 
                        (N90)? mem[481] : 
                        (N92)? mem[543] : 
                        (N94)? mem[605] : 
                        (N96)? mem[667] : 
                        (N98)? mem[729] : 
                        (N100)? mem[791] : 
                        (N102)? mem[853] : 
                        (N104)? mem[915] : 
                        (N106)? mem[977] : 
                        (N108)? mem[1039] : 
                        (N110)? mem[1101] : 
                        (N112)? mem[1163] : 
                        (N114)? mem[1225] : 
                        (N116)? mem[1287] : 
                        (N118)? mem[1349] : 
                        (N120)? mem[1411] : 
                        (N122)? mem[1473] : 
                        (N124)? mem[1535] : 
                        (N126)? mem[1597] : 
                        (N128)? mem[1659] : 
                        (N130)? mem[1721] : 
                        (N132)? mem[1783] : 
                        (N134)? mem[1845] : 
                        (N136)? mem[1907] : 
                        (N138)? mem[1969] : 
                        (N77)? mem[2031] : 
                        (N79)? mem[2093] : 
                        (N81)? mem[2155] : 
                        (N83)? mem[2217] : 
                        (N85)? mem[2279] : 
                        (N87)? mem[2341] : 
                        (N89)? mem[2403] : 
                        (N91)? mem[2465] : 
                        (N93)? mem[2527] : 
                        (N95)? mem[2589] : 
                        (N97)? mem[2651] : 
                        (N99)? mem[2713] : 
                        (N101)? mem[2775] : 
                        (N103)? mem[2837] : 
                        (N105)? mem[2899] : 
                        (N107)? mem[2961] : 
                        (N109)? mem[3023] : 
                        (N111)? mem[3085] : 
                        (N113)? mem[3147] : 
                        (N115)? mem[3209] : 
                        (N117)? mem[3271] : 
                        (N119)? mem[3333] : 
                        (N121)? mem[3395] : 
                        (N123)? mem[3457] : 
                        (N125)? mem[3519] : 
                        (N127)? mem[3581] : 
                        (N129)? mem[3643] : 
                        (N131)? mem[3705] : 
                        (N133)? mem[3767] : 
                        (N135)? mem[3829] : 
                        (N137)? mem[3891] : 
                        (N139)? mem[3953] : 1'b0;
  assign r_data_o[46] = (N76)? mem[46] : 
                        (N78)? mem[108] : 
                        (N80)? mem[170] : 
                        (N82)? mem[232] : 
                        (N84)? mem[294] : 
                        (N86)? mem[356] : 
                        (N88)? mem[418] : 
                        (N90)? mem[480] : 
                        (N92)? mem[542] : 
                        (N94)? mem[604] : 
                        (N96)? mem[666] : 
                        (N98)? mem[728] : 
                        (N100)? mem[790] : 
                        (N102)? mem[852] : 
                        (N104)? mem[914] : 
                        (N106)? mem[976] : 
                        (N108)? mem[1038] : 
                        (N110)? mem[1100] : 
                        (N112)? mem[1162] : 
                        (N114)? mem[1224] : 
                        (N116)? mem[1286] : 
                        (N118)? mem[1348] : 
                        (N120)? mem[1410] : 
                        (N122)? mem[1472] : 
                        (N124)? mem[1534] : 
                        (N126)? mem[1596] : 
                        (N128)? mem[1658] : 
                        (N130)? mem[1720] : 
                        (N132)? mem[1782] : 
                        (N134)? mem[1844] : 
                        (N136)? mem[1906] : 
                        (N138)? mem[1968] : 
                        (N77)? mem[2030] : 
                        (N79)? mem[2092] : 
                        (N81)? mem[2154] : 
                        (N83)? mem[2216] : 
                        (N85)? mem[2278] : 
                        (N87)? mem[2340] : 
                        (N89)? mem[2402] : 
                        (N91)? mem[2464] : 
                        (N93)? mem[2526] : 
                        (N95)? mem[2588] : 
                        (N97)? mem[2650] : 
                        (N99)? mem[2712] : 
                        (N101)? mem[2774] : 
                        (N103)? mem[2836] : 
                        (N105)? mem[2898] : 
                        (N107)? mem[2960] : 
                        (N109)? mem[3022] : 
                        (N111)? mem[3084] : 
                        (N113)? mem[3146] : 
                        (N115)? mem[3208] : 
                        (N117)? mem[3270] : 
                        (N119)? mem[3332] : 
                        (N121)? mem[3394] : 
                        (N123)? mem[3456] : 
                        (N125)? mem[3518] : 
                        (N127)? mem[3580] : 
                        (N129)? mem[3642] : 
                        (N131)? mem[3704] : 
                        (N133)? mem[3766] : 
                        (N135)? mem[3828] : 
                        (N137)? mem[3890] : 
                        (N139)? mem[3952] : 1'b0;
  assign r_data_o[45] = (N76)? mem[45] : 
                        (N78)? mem[107] : 
                        (N80)? mem[169] : 
                        (N82)? mem[231] : 
                        (N84)? mem[293] : 
                        (N86)? mem[355] : 
                        (N88)? mem[417] : 
                        (N90)? mem[479] : 
                        (N92)? mem[541] : 
                        (N94)? mem[603] : 
                        (N96)? mem[665] : 
                        (N98)? mem[727] : 
                        (N100)? mem[789] : 
                        (N102)? mem[851] : 
                        (N104)? mem[913] : 
                        (N106)? mem[975] : 
                        (N108)? mem[1037] : 
                        (N110)? mem[1099] : 
                        (N112)? mem[1161] : 
                        (N114)? mem[1223] : 
                        (N116)? mem[1285] : 
                        (N118)? mem[1347] : 
                        (N120)? mem[1409] : 
                        (N122)? mem[1471] : 
                        (N124)? mem[1533] : 
                        (N126)? mem[1595] : 
                        (N128)? mem[1657] : 
                        (N130)? mem[1719] : 
                        (N132)? mem[1781] : 
                        (N134)? mem[1843] : 
                        (N136)? mem[1905] : 
                        (N138)? mem[1967] : 
                        (N77)? mem[2029] : 
                        (N79)? mem[2091] : 
                        (N81)? mem[2153] : 
                        (N83)? mem[2215] : 
                        (N85)? mem[2277] : 
                        (N87)? mem[2339] : 
                        (N89)? mem[2401] : 
                        (N91)? mem[2463] : 
                        (N93)? mem[2525] : 
                        (N95)? mem[2587] : 
                        (N97)? mem[2649] : 
                        (N99)? mem[2711] : 
                        (N101)? mem[2773] : 
                        (N103)? mem[2835] : 
                        (N105)? mem[2897] : 
                        (N107)? mem[2959] : 
                        (N109)? mem[3021] : 
                        (N111)? mem[3083] : 
                        (N113)? mem[3145] : 
                        (N115)? mem[3207] : 
                        (N117)? mem[3269] : 
                        (N119)? mem[3331] : 
                        (N121)? mem[3393] : 
                        (N123)? mem[3455] : 
                        (N125)? mem[3517] : 
                        (N127)? mem[3579] : 
                        (N129)? mem[3641] : 
                        (N131)? mem[3703] : 
                        (N133)? mem[3765] : 
                        (N135)? mem[3827] : 
                        (N137)? mem[3889] : 
                        (N139)? mem[3951] : 1'b0;
  assign r_data_o[44] = (N76)? mem[44] : 
                        (N78)? mem[106] : 
                        (N80)? mem[168] : 
                        (N82)? mem[230] : 
                        (N84)? mem[292] : 
                        (N86)? mem[354] : 
                        (N88)? mem[416] : 
                        (N90)? mem[478] : 
                        (N92)? mem[540] : 
                        (N94)? mem[602] : 
                        (N96)? mem[664] : 
                        (N98)? mem[726] : 
                        (N100)? mem[788] : 
                        (N102)? mem[850] : 
                        (N104)? mem[912] : 
                        (N106)? mem[974] : 
                        (N108)? mem[1036] : 
                        (N110)? mem[1098] : 
                        (N112)? mem[1160] : 
                        (N114)? mem[1222] : 
                        (N116)? mem[1284] : 
                        (N118)? mem[1346] : 
                        (N120)? mem[1408] : 
                        (N122)? mem[1470] : 
                        (N124)? mem[1532] : 
                        (N126)? mem[1594] : 
                        (N128)? mem[1656] : 
                        (N130)? mem[1718] : 
                        (N132)? mem[1780] : 
                        (N134)? mem[1842] : 
                        (N136)? mem[1904] : 
                        (N138)? mem[1966] : 
                        (N77)? mem[2028] : 
                        (N79)? mem[2090] : 
                        (N81)? mem[2152] : 
                        (N83)? mem[2214] : 
                        (N85)? mem[2276] : 
                        (N87)? mem[2338] : 
                        (N89)? mem[2400] : 
                        (N91)? mem[2462] : 
                        (N93)? mem[2524] : 
                        (N95)? mem[2586] : 
                        (N97)? mem[2648] : 
                        (N99)? mem[2710] : 
                        (N101)? mem[2772] : 
                        (N103)? mem[2834] : 
                        (N105)? mem[2896] : 
                        (N107)? mem[2958] : 
                        (N109)? mem[3020] : 
                        (N111)? mem[3082] : 
                        (N113)? mem[3144] : 
                        (N115)? mem[3206] : 
                        (N117)? mem[3268] : 
                        (N119)? mem[3330] : 
                        (N121)? mem[3392] : 
                        (N123)? mem[3454] : 
                        (N125)? mem[3516] : 
                        (N127)? mem[3578] : 
                        (N129)? mem[3640] : 
                        (N131)? mem[3702] : 
                        (N133)? mem[3764] : 
                        (N135)? mem[3826] : 
                        (N137)? mem[3888] : 
                        (N139)? mem[3950] : 1'b0;
  assign r_data_o[43] = (N76)? mem[43] : 
                        (N78)? mem[105] : 
                        (N80)? mem[167] : 
                        (N82)? mem[229] : 
                        (N84)? mem[291] : 
                        (N86)? mem[353] : 
                        (N88)? mem[415] : 
                        (N90)? mem[477] : 
                        (N92)? mem[539] : 
                        (N94)? mem[601] : 
                        (N96)? mem[663] : 
                        (N98)? mem[725] : 
                        (N100)? mem[787] : 
                        (N102)? mem[849] : 
                        (N104)? mem[911] : 
                        (N106)? mem[973] : 
                        (N108)? mem[1035] : 
                        (N110)? mem[1097] : 
                        (N112)? mem[1159] : 
                        (N114)? mem[1221] : 
                        (N116)? mem[1283] : 
                        (N118)? mem[1345] : 
                        (N120)? mem[1407] : 
                        (N122)? mem[1469] : 
                        (N124)? mem[1531] : 
                        (N126)? mem[1593] : 
                        (N128)? mem[1655] : 
                        (N130)? mem[1717] : 
                        (N132)? mem[1779] : 
                        (N134)? mem[1841] : 
                        (N136)? mem[1903] : 
                        (N138)? mem[1965] : 
                        (N77)? mem[2027] : 
                        (N79)? mem[2089] : 
                        (N81)? mem[2151] : 
                        (N83)? mem[2213] : 
                        (N85)? mem[2275] : 
                        (N87)? mem[2337] : 
                        (N89)? mem[2399] : 
                        (N91)? mem[2461] : 
                        (N93)? mem[2523] : 
                        (N95)? mem[2585] : 
                        (N97)? mem[2647] : 
                        (N99)? mem[2709] : 
                        (N101)? mem[2771] : 
                        (N103)? mem[2833] : 
                        (N105)? mem[2895] : 
                        (N107)? mem[2957] : 
                        (N109)? mem[3019] : 
                        (N111)? mem[3081] : 
                        (N113)? mem[3143] : 
                        (N115)? mem[3205] : 
                        (N117)? mem[3267] : 
                        (N119)? mem[3329] : 
                        (N121)? mem[3391] : 
                        (N123)? mem[3453] : 
                        (N125)? mem[3515] : 
                        (N127)? mem[3577] : 
                        (N129)? mem[3639] : 
                        (N131)? mem[3701] : 
                        (N133)? mem[3763] : 
                        (N135)? mem[3825] : 
                        (N137)? mem[3887] : 
                        (N139)? mem[3949] : 1'b0;
  assign r_data_o[42] = (N76)? mem[42] : 
                        (N78)? mem[104] : 
                        (N80)? mem[166] : 
                        (N82)? mem[228] : 
                        (N84)? mem[290] : 
                        (N86)? mem[352] : 
                        (N88)? mem[414] : 
                        (N90)? mem[476] : 
                        (N92)? mem[538] : 
                        (N94)? mem[600] : 
                        (N96)? mem[662] : 
                        (N98)? mem[724] : 
                        (N100)? mem[786] : 
                        (N102)? mem[848] : 
                        (N104)? mem[910] : 
                        (N106)? mem[972] : 
                        (N108)? mem[1034] : 
                        (N110)? mem[1096] : 
                        (N112)? mem[1158] : 
                        (N114)? mem[1220] : 
                        (N116)? mem[1282] : 
                        (N118)? mem[1344] : 
                        (N120)? mem[1406] : 
                        (N122)? mem[1468] : 
                        (N124)? mem[1530] : 
                        (N126)? mem[1592] : 
                        (N128)? mem[1654] : 
                        (N130)? mem[1716] : 
                        (N132)? mem[1778] : 
                        (N134)? mem[1840] : 
                        (N136)? mem[1902] : 
                        (N138)? mem[1964] : 
                        (N77)? mem[2026] : 
                        (N79)? mem[2088] : 
                        (N81)? mem[2150] : 
                        (N83)? mem[2212] : 
                        (N85)? mem[2274] : 
                        (N87)? mem[2336] : 
                        (N89)? mem[2398] : 
                        (N91)? mem[2460] : 
                        (N93)? mem[2522] : 
                        (N95)? mem[2584] : 
                        (N97)? mem[2646] : 
                        (N99)? mem[2708] : 
                        (N101)? mem[2770] : 
                        (N103)? mem[2832] : 
                        (N105)? mem[2894] : 
                        (N107)? mem[2956] : 
                        (N109)? mem[3018] : 
                        (N111)? mem[3080] : 
                        (N113)? mem[3142] : 
                        (N115)? mem[3204] : 
                        (N117)? mem[3266] : 
                        (N119)? mem[3328] : 
                        (N121)? mem[3390] : 
                        (N123)? mem[3452] : 
                        (N125)? mem[3514] : 
                        (N127)? mem[3576] : 
                        (N129)? mem[3638] : 
                        (N131)? mem[3700] : 
                        (N133)? mem[3762] : 
                        (N135)? mem[3824] : 
                        (N137)? mem[3886] : 
                        (N139)? mem[3948] : 1'b0;
  assign r_data_o[41] = (N76)? mem[41] : 
                        (N78)? mem[103] : 
                        (N80)? mem[165] : 
                        (N82)? mem[227] : 
                        (N84)? mem[289] : 
                        (N86)? mem[351] : 
                        (N88)? mem[413] : 
                        (N90)? mem[475] : 
                        (N92)? mem[537] : 
                        (N94)? mem[599] : 
                        (N96)? mem[661] : 
                        (N98)? mem[723] : 
                        (N100)? mem[785] : 
                        (N102)? mem[847] : 
                        (N104)? mem[909] : 
                        (N106)? mem[971] : 
                        (N108)? mem[1033] : 
                        (N110)? mem[1095] : 
                        (N112)? mem[1157] : 
                        (N114)? mem[1219] : 
                        (N116)? mem[1281] : 
                        (N118)? mem[1343] : 
                        (N120)? mem[1405] : 
                        (N122)? mem[1467] : 
                        (N124)? mem[1529] : 
                        (N126)? mem[1591] : 
                        (N128)? mem[1653] : 
                        (N130)? mem[1715] : 
                        (N132)? mem[1777] : 
                        (N134)? mem[1839] : 
                        (N136)? mem[1901] : 
                        (N138)? mem[1963] : 
                        (N77)? mem[2025] : 
                        (N79)? mem[2087] : 
                        (N81)? mem[2149] : 
                        (N83)? mem[2211] : 
                        (N85)? mem[2273] : 
                        (N87)? mem[2335] : 
                        (N89)? mem[2397] : 
                        (N91)? mem[2459] : 
                        (N93)? mem[2521] : 
                        (N95)? mem[2583] : 
                        (N97)? mem[2645] : 
                        (N99)? mem[2707] : 
                        (N101)? mem[2769] : 
                        (N103)? mem[2831] : 
                        (N105)? mem[2893] : 
                        (N107)? mem[2955] : 
                        (N109)? mem[3017] : 
                        (N111)? mem[3079] : 
                        (N113)? mem[3141] : 
                        (N115)? mem[3203] : 
                        (N117)? mem[3265] : 
                        (N119)? mem[3327] : 
                        (N121)? mem[3389] : 
                        (N123)? mem[3451] : 
                        (N125)? mem[3513] : 
                        (N127)? mem[3575] : 
                        (N129)? mem[3637] : 
                        (N131)? mem[3699] : 
                        (N133)? mem[3761] : 
                        (N135)? mem[3823] : 
                        (N137)? mem[3885] : 
                        (N139)? mem[3947] : 1'b0;
  assign r_data_o[40] = (N76)? mem[40] : 
                        (N78)? mem[102] : 
                        (N80)? mem[164] : 
                        (N82)? mem[226] : 
                        (N84)? mem[288] : 
                        (N86)? mem[350] : 
                        (N88)? mem[412] : 
                        (N90)? mem[474] : 
                        (N92)? mem[536] : 
                        (N94)? mem[598] : 
                        (N96)? mem[660] : 
                        (N98)? mem[722] : 
                        (N100)? mem[784] : 
                        (N102)? mem[846] : 
                        (N104)? mem[908] : 
                        (N106)? mem[970] : 
                        (N108)? mem[1032] : 
                        (N110)? mem[1094] : 
                        (N112)? mem[1156] : 
                        (N114)? mem[1218] : 
                        (N116)? mem[1280] : 
                        (N118)? mem[1342] : 
                        (N120)? mem[1404] : 
                        (N122)? mem[1466] : 
                        (N124)? mem[1528] : 
                        (N126)? mem[1590] : 
                        (N128)? mem[1652] : 
                        (N130)? mem[1714] : 
                        (N132)? mem[1776] : 
                        (N134)? mem[1838] : 
                        (N136)? mem[1900] : 
                        (N138)? mem[1962] : 
                        (N77)? mem[2024] : 
                        (N79)? mem[2086] : 
                        (N81)? mem[2148] : 
                        (N83)? mem[2210] : 
                        (N85)? mem[2272] : 
                        (N87)? mem[2334] : 
                        (N89)? mem[2396] : 
                        (N91)? mem[2458] : 
                        (N93)? mem[2520] : 
                        (N95)? mem[2582] : 
                        (N97)? mem[2644] : 
                        (N99)? mem[2706] : 
                        (N101)? mem[2768] : 
                        (N103)? mem[2830] : 
                        (N105)? mem[2892] : 
                        (N107)? mem[2954] : 
                        (N109)? mem[3016] : 
                        (N111)? mem[3078] : 
                        (N113)? mem[3140] : 
                        (N115)? mem[3202] : 
                        (N117)? mem[3264] : 
                        (N119)? mem[3326] : 
                        (N121)? mem[3388] : 
                        (N123)? mem[3450] : 
                        (N125)? mem[3512] : 
                        (N127)? mem[3574] : 
                        (N129)? mem[3636] : 
                        (N131)? mem[3698] : 
                        (N133)? mem[3760] : 
                        (N135)? mem[3822] : 
                        (N137)? mem[3884] : 
                        (N139)? mem[3946] : 1'b0;
  assign r_data_o[39] = (N76)? mem[39] : 
                        (N78)? mem[101] : 
                        (N80)? mem[163] : 
                        (N82)? mem[225] : 
                        (N84)? mem[287] : 
                        (N86)? mem[349] : 
                        (N88)? mem[411] : 
                        (N90)? mem[473] : 
                        (N92)? mem[535] : 
                        (N94)? mem[597] : 
                        (N96)? mem[659] : 
                        (N98)? mem[721] : 
                        (N100)? mem[783] : 
                        (N102)? mem[845] : 
                        (N104)? mem[907] : 
                        (N106)? mem[969] : 
                        (N108)? mem[1031] : 
                        (N110)? mem[1093] : 
                        (N112)? mem[1155] : 
                        (N114)? mem[1217] : 
                        (N116)? mem[1279] : 
                        (N118)? mem[1341] : 
                        (N120)? mem[1403] : 
                        (N122)? mem[1465] : 
                        (N124)? mem[1527] : 
                        (N126)? mem[1589] : 
                        (N128)? mem[1651] : 
                        (N130)? mem[1713] : 
                        (N132)? mem[1775] : 
                        (N134)? mem[1837] : 
                        (N136)? mem[1899] : 
                        (N138)? mem[1961] : 
                        (N77)? mem[2023] : 
                        (N79)? mem[2085] : 
                        (N81)? mem[2147] : 
                        (N83)? mem[2209] : 
                        (N85)? mem[2271] : 
                        (N87)? mem[2333] : 
                        (N89)? mem[2395] : 
                        (N91)? mem[2457] : 
                        (N93)? mem[2519] : 
                        (N95)? mem[2581] : 
                        (N97)? mem[2643] : 
                        (N99)? mem[2705] : 
                        (N101)? mem[2767] : 
                        (N103)? mem[2829] : 
                        (N105)? mem[2891] : 
                        (N107)? mem[2953] : 
                        (N109)? mem[3015] : 
                        (N111)? mem[3077] : 
                        (N113)? mem[3139] : 
                        (N115)? mem[3201] : 
                        (N117)? mem[3263] : 
                        (N119)? mem[3325] : 
                        (N121)? mem[3387] : 
                        (N123)? mem[3449] : 
                        (N125)? mem[3511] : 
                        (N127)? mem[3573] : 
                        (N129)? mem[3635] : 
                        (N131)? mem[3697] : 
                        (N133)? mem[3759] : 
                        (N135)? mem[3821] : 
                        (N137)? mem[3883] : 
                        (N139)? mem[3945] : 1'b0;
  assign r_data_o[38] = (N76)? mem[38] : 
                        (N78)? mem[100] : 
                        (N80)? mem[162] : 
                        (N82)? mem[224] : 
                        (N84)? mem[286] : 
                        (N86)? mem[348] : 
                        (N88)? mem[410] : 
                        (N90)? mem[472] : 
                        (N92)? mem[534] : 
                        (N94)? mem[596] : 
                        (N96)? mem[658] : 
                        (N98)? mem[720] : 
                        (N100)? mem[782] : 
                        (N102)? mem[844] : 
                        (N104)? mem[906] : 
                        (N106)? mem[968] : 
                        (N108)? mem[1030] : 
                        (N110)? mem[1092] : 
                        (N112)? mem[1154] : 
                        (N114)? mem[1216] : 
                        (N116)? mem[1278] : 
                        (N118)? mem[1340] : 
                        (N120)? mem[1402] : 
                        (N122)? mem[1464] : 
                        (N124)? mem[1526] : 
                        (N126)? mem[1588] : 
                        (N128)? mem[1650] : 
                        (N130)? mem[1712] : 
                        (N132)? mem[1774] : 
                        (N134)? mem[1836] : 
                        (N136)? mem[1898] : 
                        (N138)? mem[1960] : 
                        (N77)? mem[2022] : 
                        (N79)? mem[2084] : 
                        (N81)? mem[2146] : 
                        (N83)? mem[2208] : 
                        (N85)? mem[2270] : 
                        (N87)? mem[2332] : 
                        (N89)? mem[2394] : 
                        (N91)? mem[2456] : 
                        (N93)? mem[2518] : 
                        (N95)? mem[2580] : 
                        (N97)? mem[2642] : 
                        (N99)? mem[2704] : 
                        (N101)? mem[2766] : 
                        (N103)? mem[2828] : 
                        (N105)? mem[2890] : 
                        (N107)? mem[2952] : 
                        (N109)? mem[3014] : 
                        (N111)? mem[3076] : 
                        (N113)? mem[3138] : 
                        (N115)? mem[3200] : 
                        (N117)? mem[3262] : 
                        (N119)? mem[3324] : 
                        (N121)? mem[3386] : 
                        (N123)? mem[3448] : 
                        (N125)? mem[3510] : 
                        (N127)? mem[3572] : 
                        (N129)? mem[3634] : 
                        (N131)? mem[3696] : 
                        (N133)? mem[3758] : 
                        (N135)? mem[3820] : 
                        (N137)? mem[3882] : 
                        (N139)? mem[3944] : 1'b0;
  assign r_data_o[37] = (N76)? mem[37] : 
                        (N78)? mem[99] : 
                        (N80)? mem[161] : 
                        (N82)? mem[223] : 
                        (N84)? mem[285] : 
                        (N86)? mem[347] : 
                        (N88)? mem[409] : 
                        (N90)? mem[471] : 
                        (N92)? mem[533] : 
                        (N94)? mem[595] : 
                        (N96)? mem[657] : 
                        (N98)? mem[719] : 
                        (N100)? mem[781] : 
                        (N102)? mem[843] : 
                        (N104)? mem[905] : 
                        (N106)? mem[967] : 
                        (N108)? mem[1029] : 
                        (N110)? mem[1091] : 
                        (N112)? mem[1153] : 
                        (N114)? mem[1215] : 
                        (N116)? mem[1277] : 
                        (N118)? mem[1339] : 
                        (N120)? mem[1401] : 
                        (N122)? mem[1463] : 
                        (N124)? mem[1525] : 
                        (N126)? mem[1587] : 
                        (N128)? mem[1649] : 
                        (N130)? mem[1711] : 
                        (N132)? mem[1773] : 
                        (N134)? mem[1835] : 
                        (N136)? mem[1897] : 
                        (N138)? mem[1959] : 
                        (N77)? mem[2021] : 
                        (N79)? mem[2083] : 
                        (N81)? mem[2145] : 
                        (N83)? mem[2207] : 
                        (N85)? mem[2269] : 
                        (N87)? mem[2331] : 
                        (N89)? mem[2393] : 
                        (N91)? mem[2455] : 
                        (N93)? mem[2517] : 
                        (N95)? mem[2579] : 
                        (N97)? mem[2641] : 
                        (N99)? mem[2703] : 
                        (N101)? mem[2765] : 
                        (N103)? mem[2827] : 
                        (N105)? mem[2889] : 
                        (N107)? mem[2951] : 
                        (N109)? mem[3013] : 
                        (N111)? mem[3075] : 
                        (N113)? mem[3137] : 
                        (N115)? mem[3199] : 
                        (N117)? mem[3261] : 
                        (N119)? mem[3323] : 
                        (N121)? mem[3385] : 
                        (N123)? mem[3447] : 
                        (N125)? mem[3509] : 
                        (N127)? mem[3571] : 
                        (N129)? mem[3633] : 
                        (N131)? mem[3695] : 
                        (N133)? mem[3757] : 
                        (N135)? mem[3819] : 
                        (N137)? mem[3881] : 
                        (N139)? mem[3943] : 1'b0;
  assign r_data_o[36] = (N76)? mem[36] : 
                        (N78)? mem[98] : 
                        (N80)? mem[160] : 
                        (N82)? mem[222] : 
                        (N84)? mem[284] : 
                        (N86)? mem[346] : 
                        (N88)? mem[408] : 
                        (N90)? mem[470] : 
                        (N92)? mem[532] : 
                        (N94)? mem[594] : 
                        (N96)? mem[656] : 
                        (N98)? mem[718] : 
                        (N100)? mem[780] : 
                        (N102)? mem[842] : 
                        (N104)? mem[904] : 
                        (N106)? mem[966] : 
                        (N108)? mem[1028] : 
                        (N110)? mem[1090] : 
                        (N112)? mem[1152] : 
                        (N114)? mem[1214] : 
                        (N116)? mem[1276] : 
                        (N118)? mem[1338] : 
                        (N120)? mem[1400] : 
                        (N122)? mem[1462] : 
                        (N124)? mem[1524] : 
                        (N126)? mem[1586] : 
                        (N128)? mem[1648] : 
                        (N130)? mem[1710] : 
                        (N132)? mem[1772] : 
                        (N134)? mem[1834] : 
                        (N136)? mem[1896] : 
                        (N138)? mem[1958] : 
                        (N77)? mem[2020] : 
                        (N79)? mem[2082] : 
                        (N81)? mem[2144] : 
                        (N83)? mem[2206] : 
                        (N85)? mem[2268] : 
                        (N87)? mem[2330] : 
                        (N89)? mem[2392] : 
                        (N91)? mem[2454] : 
                        (N93)? mem[2516] : 
                        (N95)? mem[2578] : 
                        (N97)? mem[2640] : 
                        (N99)? mem[2702] : 
                        (N101)? mem[2764] : 
                        (N103)? mem[2826] : 
                        (N105)? mem[2888] : 
                        (N107)? mem[2950] : 
                        (N109)? mem[3012] : 
                        (N111)? mem[3074] : 
                        (N113)? mem[3136] : 
                        (N115)? mem[3198] : 
                        (N117)? mem[3260] : 
                        (N119)? mem[3322] : 
                        (N121)? mem[3384] : 
                        (N123)? mem[3446] : 
                        (N125)? mem[3508] : 
                        (N127)? mem[3570] : 
                        (N129)? mem[3632] : 
                        (N131)? mem[3694] : 
                        (N133)? mem[3756] : 
                        (N135)? mem[3818] : 
                        (N137)? mem[3880] : 
                        (N139)? mem[3942] : 1'b0;
  assign r_data_o[35] = (N76)? mem[35] : 
                        (N78)? mem[97] : 
                        (N80)? mem[159] : 
                        (N82)? mem[221] : 
                        (N84)? mem[283] : 
                        (N86)? mem[345] : 
                        (N88)? mem[407] : 
                        (N90)? mem[469] : 
                        (N92)? mem[531] : 
                        (N94)? mem[593] : 
                        (N96)? mem[655] : 
                        (N98)? mem[717] : 
                        (N100)? mem[779] : 
                        (N102)? mem[841] : 
                        (N104)? mem[903] : 
                        (N106)? mem[965] : 
                        (N108)? mem[1027] : 
                        (N110)? mem[1089] : 
                        (N112)? mem[1151] : 
                        (N114)? mem[1213] : 
                        (N116)? mem[1275] : 
                        (N118)? mem[1337] : 
                        (N120)? mem[1399] : 
                        (N122)? mem[1461] : 
                        (N124)? mem[1523] : 
                        (N126)? mem[1585] : 
                        (N128)? mem[1647] : 
                        (N130)? mem[1709] : 
                        (N132)? mem[1771] : 
                        (N134)? mem[1833] : 
                        (N136)? mem[1895] : 
                        (N138)? mem[1957] : 
                        (N77)? mem[2019] : 
                        (N79)? mem[2081] : 
                        (N81)? mem[2143] : 
                        (N83)? mem[2205] : 
                        (N85)? mem[2267] : 
                        (N87)? mem[2329] : 
                        (N89)? mem[2391] : 
                        (N91)? mem[2453] : 
                        (N93)? mem[2515] : 
                        (N95)? mem[2577] : 
                        (N97)? mem[2639] : 
                        (N99)? mem[2701] : 
                        (N101)? mem[2763] : 
                        (N103)? mem[2825] : 
                        (N105)? mem[2887] : 
                        (N107)? mem[2949] : 
                        (N109)? mem[3011] : 
                        (N111)? mem[3073] : 
                        (N113)? mem[3135] : 
                        (N115)? mem[3197] : 
                        (N117)? mem[3259] : 
                        (N119)? mem[3321] : 
                        (N121)? mem[3383] : 
                        (N123)? mem[3445] : 
                        (N125)? mem[3507] : 
                        (N127)? mem[3569] : 
                        (N129)? mem[3631] : 
                        (N131)? mem[3693] : 
                        (N133)? mem[3755] : 
                        (N135)? mem[3817] : 
                        (N137)? mem[3879] : 
                        (N139)? mem[3941] : 1'b0;
  assign r_data_o[34] = (N76)? mem[34] : 
                        (N78)? mem[96] : 
                        (N80)? mem[158] : 
                        (N82)? mem[220] : 
                        (N84)? mem[282] : 
                        (N86)? mem[344] : 
                        (N88)? mem[406] : 
                        (N90)? mem[468] : 
                        (N92)? mem[530] : 
                        (N94)? mem[592] : 
                        (N96)? mem[654] : 
                        (N98)? mem[716] : 
                        (N100)? mem[778] : 
                        (N102)? mem[840] : 
                        (N104)? mem[902] : 
                        (N106)? mem[964] : 
                        (N108)? mem[1026] : 
                        (N110)? mem[1088] : 
                        (N112)? mem[1150] : 
                        (N114)? mem[1212] : 
                        (N116)? mem[1274] : 
                        (N118)? mem[1336] : 
                        (N120)? mem[1398] : 
                        (N122)? mem[1460] : 
                        (N124)? mem[1522] : 
                        (N126)? mem[1584] : 
                        (N128)? mem[1646] : 
                        (N130)? mem[1708] : 
                        (N132)? mem[1770] : 
                        (N134)? mem[1832] : 
                        (N136)? mem[1894] : 
                        (N138)? mem[1956] : 
                        (N77)? mem[2018] : 
                        (N79)? mem[2080] : 
                        (N81)? mem[2142] : 
                        (N83)? mem[2204] : 
                        (N85)? mem[2266] : 
                        (N87)? mem[2328] : 
                        (N89)? mem[2390] : 
                        (N91)? mem[2452] : 
                        (N93)? mem[2514] : 
                        (N95)? mem[2576] : 
                        (N97)? mem[2638] : 
                        (N99)? mem[2700] : 
                        (N101)? mem[2762] : 
                        (N103)? mem[2824] : 
                        (N105)? mem[2886] : 
                        (N107)? mem[2948] : 
                        (N109)? mem[3010] : 
                        (N111)? mem[3072] : 
                        (N113)? mem[3134] : 
                        (N115)? mem[3196] : 
                        (N117)? mem[3258] : 
                        (N119)? mem[3320] : 
                        (N121)? mem[3382] : 
                        (N123)? mem[3444] : 
                        (N125)? mem[3506] : 
                        (N127)? mem[3568] : 
                        (N129)? mem[3630] : 
                        (N131)? mem[3692] : 
                        (N133)? mem[3754] : 
                        (N135)? mem[3816] : 
                        (N137)? mem[3878] : 
                        (N139)? mem[3940] : 1'b0;
  assign r_data_o[33] = (N76)? mem[33] : 
                        (N78)? mem[95] : 
                        (N80)? mem[157] : 
                        (N82)? mem[219] : 
                        (N84)? mem[281] : 
                        (N86)? mem[343] : 
                        (N88)? mem[405] : 
                        (N90)? mem[467] : 
                        (N92)? mem[529] : 
                        (N94)? mem[591] : 
                        (N96)? mem[653] : 
                        (N98)? mem[715] : 
                        (N100)? mem[777] : 
                        (N102)? mem[839] : 
                        (N104)? mem[901] : 
                        (N106)? mem[963] : 
                        (N108)? mem[1025] : 
                        (N110)? mem[1087] : 
                        (N112)? mem[1149] : 
                        (N114)? mem[1211] : 
                        (N116)? mem[1273] : 
                        (N118)? mem[1335] : 
                        (N120)? mem[1397] : 
                        (N122)? mem[1459] : 
                        (N124)? mem[1521] : 
                        (N126)? mem[1583] : 
                        (N128)? mem[1645] : 
                        (N130)? mem[1707] : 
                        (N132)? mem[1769] : 
                        (N134)? mem[1831] : 
                        (N136)? mem[1893] : 
                        (N138)? mem[1955] : 
                        (N77)? mem[2017] : 
                        (N79)? mem[2079] : 
                        (N81)? mem[2141] : 
                        (N83)? mem[2203] : 
                        (N85)? mem[2265] : 
                        (N87)? mem[2327] : 
                        (N89)? mem[2389] : 
                        (N91)? mem[2451] : 
                        (N93)? mem[2513] : 
                        (N95)? mem[2575] : 
                        (N97)? mem[2637] : 
                        (N99)? mem[2699] : 
                        (N101)? mem[2761] : 
                        (N103)? mem[2823] : 
                        (N105)? mem[2885] : 
                        (N107)? mem[2947] : 
                        (N109)? mem[3009] : 
                        (N111)? mem[3071] : 
                        (N113)? mem[3133] : 
                        (N115)? mem[3195] : 
                        (N117)? mem[3257] : 
                        (N119)? mem[3319] : 
                        (N121)? mem[3381] : 
                        (N123)? mem[3443] : 
                        (N125)? mem[3505] : 
                        (N127)? mem[3567] : 
                        (N129)? mem[3629] : 
                        (N131)? mem[3691] : 
                        (N133)? mem[3753] : 
                        (N135)? mem[3815] : 
                        (N137)? mem[3877] : 
                        (N139)? mem[3939] : 1'b0;
  assign r_data_o[32] = (N76)? mem[32] : 
                        (N78)? mem[94] : 
                        (N80)? mem[156] : 
                        (N82)? mem[218] : 
                        (N84)? mem[280] : 
                        (N86)? mem[342] : 
                        (N88)? mem[404] : 
                        (N90)? mem[466] : 
                        (N92)? mem[528] : 
                        (N94)? mem[590] : 
                        (N96)? mem[652] : 
                        (N98)? mem[714] : 
                        (N100)? mem[776] : 
                        (N102)? mem[838] : 
                        (N104)? mem[900] : 
                        (N106)? mem[962] : 
                        (N108)? mem[1024] : 
                        (N110)? mem[1086] : 
                        (N112)? mem[1148] : 
                        (N114)? mem[1210] : 
                        (N116)? mem[1272] : 
                        (N118)? mem[1334] : 
                        (N120)? mem[1396] : 
                        (N122)? mem[1458] : 
                        (N124)? mem[1520] : 
                        (N126)? mem[1582] : 
                        (N128)? mem[1644] : 
                        (N130)? mem[1706] : 
                        (N132)? mem[1768] : 
                        (N134)? mem[1830] : 
                        (N136)? mem[1892] : 
                        (N138)? mem[1954] : 
                        (N77)? mem[2016] : 
                        (N79)? mem[2078] : 
                        (N81)? mem[2140] : 
                        (N83)? mem[2202] : 
                        (N85)? mem[2264] : 
                        (N87)? mem[2326] : 
                        (N89)? mem[2388] : 
                        (N91)? mem[2450] : 
                        (N93)? mem[2512] : 
                        (N95)? mem[2574] : 
                        (N97)? mem[2636] : 
                        (N99)? mem[2698] : 
                        (N101)? mem[2760] : 
                        (N103)? mem[2822] : 
                        (N105)? mem[2884] : 
                        (N107)? mem[2946] : 
                        (N109)? mem[3008] : 
                        (N111)? mem[3070] : 
                        (N113)? mem[3132] : 
                        (N115)? mem[3194] : 
                        (N117)? mem[3256] : 
                        (N119)? mem[3318] : 
                        (N121)? mem[3380] : 
                        (N123)? mem[3442] : 
                        (N125)? mem[3504] : 
                        (N127)? mem[3566] : 
                        (N129)? mem[3628] : 
                        (N131)? mem[3690] : 
                        (N133)? mem[3752] : 
                        (N135)? mem[3814] : 
                        (N137)? mem[3876] : 
                        (N139)? mem[3938] : 1'b0;
  assign r_data_o[31] = (N76)? mem[31] : 
                        (N78)? mem[93] : 
                        (N80)? mem[155] : 
                        (N82)? mem[217] : 
                        (N84)? mem[279] : 
                        (N86)? mem[341] : 
                        (N88)? mem[403] : 
                        (N90)? mem[465] : 
                        (N92)? mem[527] : 
                        (N94)? mem[589] : 
                        (N96)? mem[651] : 
                        (N98)? mem[713] : 
                        (N100)? mem[775] : 
                        (N102)? mem[837] : 
                        (N104)? mem[899] : 
                        (N106)? mem[961] : 
                        (N108)? mem[1023] : 
                        (N110)? mem[1085] : 
                        (N112)? mem[1147] : 
                        (N114)? mem[1209] : 
                        (N116)? mem[1271] : 
                        (N118)? mem[1333] : 
                        (N120)? mem[1395] : 
                        (N122)? mem[1457] : 
                        (N124)? mem[1519] : 
                        (N126)? mem[1581] : 
                        (N128)? mem[1643] : 
                        (N130)? mem[1705] : 
                        (N132)? mem[1767] : 
                        (N134)? mem[1829] : 
                        (N136)? mem[1891] : 
                        (N138)? mem[1953] : 
                        (N77)? mem[2015] : 
                        (N79)? mem[2077] : 
                        (N81)? mem[2139] : 
                        (N83)? mem[2201] : 
                        (N85)? mem[2263] : 
                        (N87)? mem[2325] : 
                        (N89)? mem[2387] : 
                        (N91)? mem[2449] : 
                        (N93)? mem[2511] : 
                        (N95)? mem[2573] : 
                        (N97)? mem[2635] : 
                        (N99)? mem[2697] : 
                        (N101)? mem[2759] : 
                        (N103)? mem[2821] : 
                        (N105)? mem[2883] : 
                        (N107)? mem[2945] : 
                        (N109)? mem[3007] : 
                        (N111)? mem[3069] : 
                        (N113)? mem[3131] : 
                        (N115)? mem[3193] : 
                        (N117)? mem[3255] : 
                        (N119)? mem[3317] : 
                        (N121)? mem[3379] : 
                        (N123)? mem[3441] : 
                        (N125)? mem[3503] : 
                        (N127)? mem[3565] : 
                        (N129)? mem[3627] : 
                        (N131)? mem[3689] : 
                        (N133)? mem[3751] : 
                        (N135)? mem[3813] : 
                        (N137)? mem[3875] : 
                        (N139)? mem[3937] : 1'b0;
  assign r_data_o[30] = (N76)? mem[30] : 
                        (N78)? mem[92] : 
                        (N80)? mem[154] : 
                        (N82)? mem[216] : 
                        (N84)? mem[278] : 
                        (N86)? mem[340] : 
                        (N88)? mem[402] : 
                        (N90)? mem[464] : 
                        (N92)? mem[526] : 
                        (N94)? mem[588] : 
                        (N96)? mem[650] : 
                        (N98)? mem[712] : 
                        (N100)? mem[774] : 
                        (N102)? mem[836] : 
                        (N104)? mem[898] : 
                        (N106)? mem[960] : 
                        (N108)? mem[1022] : 
                        (N110)? mem[1084] : 
                        (N112)? mem[1146] : 
                        (N114)? mem[1208] : 
                        (N116)? mem[1270] : 
                        (N118)? mem[1332] : 
                        (N120)? mem[1394] : 
                        (N122)? mem[1456] : 
                        (N124)? mem[1518] : 
                        (N126)? mem[1580] : 
                        (N128)? mem[1642] : 
                        (N130)? mem[1704] : 
                        (N132)? mem[1766] : 
                        (N134)? mem[1828] : 
                        (N136)? mem[1890] : 
                        (N138)? mem[1952] : 
                        (N77)? mem[2014] : 
                        (N79)? mem[2076] : 
                        (N81)? mem[2138] : 
                        (N83)? mem[2200] : 
                        (N85)? mem[2262] : 
                        (N87)? mem[2324] : 
                        (N89)? mem[2386] : 
                        (N91)? mem[2448] : 
                        (N93)? mem[2510] : 
                        (N95)? mem[2572] : 
                        (N97)? mem[2634] : 
                        (N99)? mem[2696] : 
                        (N101)? mem[2758] : 
                        (N103)? mem[2820] : 
                        (N105)? mem[2882] : 
                        (N107)? mem[2944] : 
                        (N109)? mem[3006] : 
                        (N111)? mem[3068] : 
                        (N113)? mem[3130] : 
                        (N115)? mem[3192] : 
                        (N117)? mem[3254] : 
                        (N119)? mem[3316] : 
                        (N121)? mem[3378] : 
                        (N123)? mem[3440] : 
                        (N125)? mem[3502] : 
                        (N127)? mem[3564] : 
                        (N129)? mem[3626] : 
                        (N131)? mem[3688] : 
                        (N133)? mem[3750] : 
                        (N135)? mem[3812] : 
                        (N137)? mem[3874] : 
                        (N139)? mem[3936] : 1'b0;
  assign r_data_o[29] = (N76)? mem[29] : 
                        (N78)? mem[91] : 
                        (N80)? mem[153] : 
                        (N82)? mem[215] : 
                        (N84)? mem[277] : 
                        (N86)? mem[339] : 
                        (N88)? mem[401] : 
                        (N90)? mem[463] : 
                        (N92)? mem[525] : 
                        (N94)? mem[587] : 
                        (N96)? mem[649] : 
                        (N98)? mem[711] : 
                        (N100)? mem[773] : 
                        (N102)? mem[835] : 
                        (N104)? mem[897] : 
                        (N106)? mem[959] : 
                        (N108)? mem[1021] : 
                        (N110)? mem[1083] : 
                        (N112)? mem[1145] : 
                        (N114)? mem[1207] : 
                        (N116)? mem[1269] : 
                        (N118)? mem[1331] : 
                        (N120)? mem[1393] : 
                        (N122)? mem[1455] : 
                        (N124)? mem[1517] : 
                        (N126)? mem[1579] : 
                        (N128)? mem[1641] : 
                        (N130)? mem[1703] : 
                        (N132)? mem[1765] : 
                        (N134)? mem[1827] : 
                        (N136)? mem[1889] : 
                        (N138)? mem[1951] : 
                        (N77)? mem[2013] : 
                        (N79)? mem[2075] : 
                        (N81)? mem[2137] : 
                        (N83)? mem[2199] : 
                        (N85)? mem[2261] : 
                        (N87)? mem[2323] : 
                        (N89)? mem[2385] : 
                        (N91)? mem[2447] : 
                        (N93)? mem[2509] : 
                        (N95)? mem[2571] : 
                        (N97)? mem[2633] : 
                        (N99)? mem[2695] : 
                        (N101)? mem[2757] : 
                        (N103)? mem[2819] : 
                        (N105)? mem[2881] : 
                        (N107)? mem[2943] : 
                        (N109)? mem[3005] : 
                        (N111)? mem[3067] : 
                        (N113)? mem[3129] : 
                        (N115)? mem[3191] : 
                        (N117)? mem[3253] : 
                        (N119)? mem[3315] : 
                        (N121)? mem[3377] : 
                        (N123)? mem[3439] : 
                        (N125)? mem[3501] : 
                        (N127)? mem[3563] : 
                        (N129)? mem[3625] : 
                        (N131)? mem[3687] : 
                        (N133)? mem[3749] : 
                        (N135)? mem[3811] : 
                        (N137)? mem[3873] : 
                        (N139)? mem[3935] : 1'b0;
  assign r_data_o[28] = (N76)? mem[28] : 
                        (N78)? mem[90] : 
                        (N80)? mem[152] : 
                        (N82)? mem[214] : 
                        (N84)? mem[276] : 
                        (N86)? mem[338] : 
                        (N88)? mem[400] : 
                        (N90)? mem[462] : 
                        (N92)? mem[524] : 
                        (N94)? mem[586] : 
                        (N96)? mem[648] : 
                        (N98)? mem[710] : 
                        (N100)? mem[772] : 
                        (N102)? mem[834] : 
                        (N104)? mem[896] : 
                        (N106)? mem[958] : 
                        (N108)? mem[1020] : 
                        (N110)? mem[1082] : 
                        (N112)? mem[1144] : 
                        (N114)? mem[1206] : 
                        (N116)? mem[1268] : 
                        (N118)? mem[1330] : 
                        (N120)? mem[1392] : 
                        (N122)? mem[1454] : 
                        (N124)? mem[1516] : 
                        (N126)? mem[1578] : 
                        (N128)? mem[1640] : 
                        (N130)? mem[1702] : 
                        (N132)? mem[1764] : 
                        (N134)? mem[1826] : 
                        (N136)? mem[1888] : 
                        (N138)? mem[1950] : 
                        (N77)? mem[2012] : 
                        (N79)? mem[2074] : 
                        (N81)? mem[2136] : 
                        (N83)? mem[2198] : 
                        (N85)? mem[2260] : 
                        (N87)? mem[2322] : 
                        (N89)? mem[2384] : 
                        (N91)? mem[2446] : 
                        (N93)? mem[2508] : 
                        (N95)? mem[2570] : 
                        (N97)? mem[2632] : 
                        (N99)? mem[2694] : 
                        (N101)? mem[2756] : 
                        (N103)? mem[2818] : 
                        (N105)? mem[2880] : 
                        (N107)? mem[2942] : 
                        (N109)? mem[3004] : 
                        (N111)? mem[3066] : 
                        (N113)? mem[3128] : 
                        (N115)? mem[3190] : 
                        (N117)? mem[3252] : 
                        (N119)? mem[3314] : 
                        (N121)? mem[3376] : 
                        (N123)? mem[3438] : 
                        (N125)? mem[3500] : 
                        (N127)? mem[3562] : 
                        (N129)? mem[3624] : 
                        (N131)? mem[3686] : 
                        (N133)? mem[3748] : 
                        (N135)? mem[3810] : 
                        (N137)? mem[3872] : 
                        (N139)? mem[3934] : 1'b0;
  assign r_data_o[27] = (N76)? mem[27] : 
                        (N78)? mem[89] : 
                        (N80)? mem[151] : 
                        (N82)? mem[213] : 
                        (N84)? mem[275] : 
                        (N86)? mem[337] : 
                        (N88)? mem[399] : 
                        (N90)? mem[461] : 
                        (N92)? mem[523] : 
                        (N94)? mem[585] : 
                        (N96)? mem[647] : 
                        (N98)? mem[709] : 
                        (N100)? mem[771] : 
                        (N102)? mem[833] : 
                        (N104)? mem[895] : 
                        (N106)? mem[957] : 
                        (N108)? mem[1019] : 
                        (N110)? mem[1081] : 
                        (N112)? mem[1143] : 
                        (N114)? mem[1205] : 
                        (N116)? mem[1267] : 
                        (N118)? mem[1329] : 
                        (N120)? mem[1391] : 
                        (N122)? mem[1453] : 
                        (N124)? mem[1515] : 
                        (N126)? mem[1577] : 
                        (N128)? mem[1639] : 
                        (N130)? mem[1701] : 
                        (N132)? mem[1763] : 
                        (N134)? mem[1825] : 
                        (N136)? mem[1887] : 
                        (N138)? mem[1949] : 
                        (N77)? mem[2011] : 
                        (N79)? mem[2073] : 
                        (N81)? mem[2135] : 
                        (N83)? mem[2197] : 
                        (N85)? mem[2259] : 
                        (N87)? mem[2321] : 
                        (N89)? mem[2383] : 
                        (N91)? mem[2445] : 
                        (N93)? mem[2507] : 
                        (N95)? mem[2569] : 
                        (N97)? mem[2631] : 
                        (N99)? mem[2693] : 
                        (N101)? mem[2755] : 
                        (N103)? mem[2817] : 
                        (N105)? mem[2879] : 
                        (N107)? mem[2941] : 
                        (N109)? mem[3003] : 
                        (N111)? mem[3065] : 
                        (N113)? mem[3127] : 
                        (N115)? mem[3189] : 
                        (N117)? mem[3251] : 
                        (N119)? mem[3313] : 
                        (N121)? mem[3375] : 
                        (N123)? mem[3437] : 
                        (N125)? mem[3499] : 
                        (N127)? mem[3561] : 
                        (N129)? mem[3623] : 
                        (N131)? mem[3685] : 
                        (N133)? mem[3747] : 
                        (N135)? mem[3809] : 
                        (N137)? mem[3871] : 
                        (N139)? mem[3933] : 1'b0;
  assign r_data_o[26] = (N76)? mem[26] : 
                        (N78)? mem[88] : 
                        (N80)? mem[150] : 
                        (N82)? mem[212] : 
                        (N84)? mem[274] : 
                        (N86)? mem[336] : 
                        (N88)? mem[398] : 
                        (N90)? mem[460] : 
                        (N92)? mem[522] : 
                        (N94)? mem[584] : 
                        (N96)? mem[646] : 
                        (N98)? mem[708] : 
                        (N100)? mem[770] : 
                        (N102)? mem[832] : 
                        (N104)? mem[894] : 
                        (N106)? mem[956] : 
                        (N108)? mem[1018] : 
                        (N110)? mem[1080] : 
                        (N112)? mem[1142] : 
                        (N114)? mem[1204] : 
                        (N116)? mem[1266] : 
                        (N118)? mem[1328] : 
                        (N120)? mem[1390] : 
                        (N122)? mem[1452] : 
                        (N124)? mem[1514] : 
                        (N126)? mem[1576] : 
                        (N128)? mem[1638] : 
                        (N130)? mem[1700] : 
                        (N132)? mem[1762] : 
                        (N134)? mem[1824] : 
                        (N136)? mem[1886] : 
                        (N138)? mem[1948] : 
                        (N77)? mem[2010] : 
                        (N79)? mem[2072] : 
                        (N81)? mem[2134] : 
                        (N83)? mem[2196] : 
                        (N85)? mem[2258] : 
                        (N87)? mem[2320] : 
                        (N89)? mem[2382] : 
                        (N91)? mem[2444] : 
                        (N93)? mem[2506] : 
                        (N95)? mem[2568] : 
                        (N97)? mem[2630] : 
                        (N99)? mem[2692] : 
                        (N101)? mem[2754] : 
                        (N103)? mem[2816] : 
                        (N105)? mem[2878] : 
                        (N107)? mem[2940] : 
                        (N109)? mem[3002] : 
                        (N111)? mem[3064] : 
                        (N113)? mem[3126] : 
                        (N115)? mem[3188] : 
                        (N117)? mem[3250] : 
                        (N119)? mem[3312] : 
                        (N121)? mem[3374] : 
                        (N123)? mem[3436] : 
                        (N125)? mem[3498] : 
                        (N127)? mem[3560] : 
                        (N129)? mem[3622] : 
                        (N131)? mem[3684] : 
                        (N133)? mem[3746] : 
                        (N135)? mem[3808] : 
                        (N137)? mem[3870] : 
                        (N139)? mem[3932] : 1'b0;
  assign r_data_o[25] = (N76)? mem[25] : 
                        (N78)? mem[87] : 
                        (N80)? mem[149] : 
                        (N82)? mem[211] : 
                        (N84)? mem[273] : 
                        (N86)? mem[335] : 
                        (N88)? mem[397] : 
                        (N90)? mem[459] : 
                        (N92)? mem[521] : 
                        (N94)? mem[583] : 
                        (N96)? mem[645] : 
                        (N98)? mem[707] : 
                        (N100)? mem[769] : 
                        (N102)? mem[831] : 
                        (N104)? mem[893] : 
                        (N106)? mem[955] : 
                        (N108)? mem[1017] : 
                        (N110)? mem[1079] : 
                        (N112)? mem[1141] : 
                        (N114)? mem[1203] : 
                        (N116)? mem[1265] : 
                        (N118)? mem[1327] : 
                        (N120)? mem[1389] : 
                        (N122)? mem[1451] : 
                        (N124)? mem[1513] : 
                        (N126)? mem[1575] : 
                        (N128)? mem[1637] : 
                        (N130)? mem[1699] : 
                        (N132)? mem[1761] : 
                        (N134)? mem[1823] : 
                        (N136)? mem[1885] : 
                        (N138)? mem[1947] : 
                        (N77)? mem[2009] : 
                        (N79)? mem[2071] : 
                        (N81)? mem[2133] : 
                        (N83)? mem[2195] : 
                        (N85)? mem[2257] : 
                        (N87)? mem[2319] : 
                        (N89)? mem[2381] : 
                        (N91)? mem[2443] : 
                        (N93)? mem[2505] : 
                        (N95)? mem[2567] : 
                        (N97)? mem[2629] : 
                        (N99)? mem[2691] : 
                        (N101)? mem[2753] : 
                        (N103)? mem[2815] : 
                        (N105)? mem[2877] : 
                        (N107)? mem[2939] : 
                        (N109)? mem[3001] : 
                        (N111)? mem[3063] : 
                        (N113)? mem[3125] : 
                        (N115)? mem[3187] : 
                        (N117)? mem[3249] : 
                        (N119)? mem[3311] : 
                        (N121)? mem[3373] : 
                        (N123)? mem[3435] : 
                        (N125)? mem[3497] : 
                        (N127)? mem[3559] : 
                        (N129)? mem[3621] : 
                        (N131)? mem[3683] : 
                        (N133)? mem[3745] : 
                        (N135)? mem[3807] : 
                        (N137)? mem[3869] : 
                        (N139)? mem[3931] : 1'b0;
  assign r_data_o[24] = (N76)? mem[24] : 
                        (N78)? mem[86] : 
                        (N80)? mem[148] : 
                        (N82)? mem[210] : 
                        (N84)? mem[272] : 
                        (N86)? mem[334] : 
                        (N88)? mem[396] : 
                        (N90)? mem[458] : 
                        (N92)? mem[520] : 
                        (N94)? mem[582] : 
                        (N96)? mem[644] : 
                        (N98)? mem[706] : 
                        (N100)? mem[768] : 
                        (N102)? mem[830] : 
                        (N104)? mem[892] : 
                        (N106)? mem[954] : 
                        (N108)? mem[1016] : 
                        (N110)? mem[1078] : 
                        (N112)? mem[1140] : 
                        (N114)? mem[1202] : 
                        (N116)? mem[1264] : 
                        (N118)? mem[1326] : 
                        (N120)? mem[1388] : 
                        (N122)? mem[1450] : 
                        (N124)? mem[1512] : 
                        (N126)? mem[1574] : 
                        (N128)? mem[1636] : 
                        (N130)? mem[1698] : 
                        (N132)? mem[1760] : 
                        (N134)? mem[1822] : 
                        (N136)? mem[1884] : 
                        (N138)? mem[1946] : 
                        (N77)? mem[2008] : 
                        (N79)? mem[2070] : 
                        (N81)? mem[2132] : 
                        (N83)? mem[2194] : 
                        (N85)? mem[2256] : 
                        (N87)? mem[2318] : 
                        (N89)? mem[2380] : 
                        (N91)? mem[2442] : 
                        (N93)? mem[2504] : 
                        (N95)? mem[2566] : 
                        (N97)? mem[2628] : 
                        (N99)? mem[2690] : 
                        (N101)? mem[2752] : 
                        (N103)? mem[2814] : 
                        (N105)? mem[2876] : 
                        (N107)? mem[2938] : 
                        (N109)? mem[3000] : 
                        (N111)? mem[3062] : 
                        (N113)? mem[3124] : 
                        (N115)? mem[3186] : 
                        (N117)? mem[3248] : 
                        (N119)? mem[3310] : 
                        (N121)? mem[3372] : 
                        (N123)? mem[3434] : 
                        (N125)? mem[3496] : 
                        (N127)? mem[3558] : 
                        (N129)? mem[3620] : 
                        (N131)? mem[3682] : 
                        (N133)? mem[3744] : 
                        (N135)? mem[3806] : 
                        (N137)? mem[3868] : 
                        (N139)? mem[3930] : 1'b0;
  assign r_data_o[23] = (N76)? mem[23] : 
                        (N78)? mem[85] : 
                        (N80)? mem[147] : 
                        (N82)? mem[209] : 
                        (N84)? mem[271] : 
                        (N86)? mem[333] : 
                        (N88)? mem[395] : 
                        (N90)? mem[457] : 
                        (N92)? mem[519] : 
                        (N94)? mem[581] : 
                        (N96)? mem[643] : 
                        (N98)? mem[705] : 
                        (N100)? mem[767] : 
                        (N102)? mem[829] : 
                        (N104)? mem[891] : 
                        (N106)? mem[953] : 
                        (N108)? mem[1015] : 
                        (N110)? mem[1077] : 
                        (N112)? mem[1139] : 
                        (N114)? mem[1201] : 
                        (N116)? mem[1263] : 
                        (N118)? mem[1325] : 
                        (N120)? mem[1387] : 
                        (N122)? mem[1449] : 
                        (N124)? mem[1511] : 
                        (N126)? mem[1573] : 
                        (N128)? mem[1635] : 
                        (N130)? mem[1697] : 
                        (N132)? mem[1759] : 
                        (N134)? mem[1821] : 
                        (N136)? mem[1883] : 
                        (N138)? mem[1945] : 
                        (N77)? mem[2007] : 
                        (N79)? mem[2069] : 
                        (N81)? mem[2131] : 
                        (N83)? mem[2193] : 
                        (N85)? mem[2255] : 
                        (N87)? mem[2317] : 
                        (N89)? mem[2379] : 
                        (N91)? mem[2441] : 
                        (N93)? mem[2503] : 
                        (N95)? mem[2565] : 
                        (N97)? mem[2627] : 
                        (N99)? mem[2689] : 
                        (N101)? mem[2751] : 
                        (N103)? mem[2813] : 
                        (N105)? mem[2875] : 
                        (N107)? mem[2937] : 
                        (N109)? mem[2999] : 
                        (N111)? mem[3061] : 
                        (N113)? mem[3123] : 
                        (N115)? mem[3185] : 
                        (N117)? mem[3247] : 
                        (N119)? mem[3309] : 
                        (N121)? mem[3371] : 
                        (N123)? mem[3433] : 
                        (N125)? mem[3495] : 
                        (N127)? mem[3557] : 
                        (N129)? mem[3619] : 
                        (N131)? mem[3681] : 
                        (N133)? mem[3743] : 
                        (N135)? mem[3805] : 
                        (N137)? mem[3867] : 
                        (N139)? mem[3929] : 1'b0;
  assign r_data_o[22] = (N76)? mem[22] : 
                        (N78)? mem[84] : 
                        (N80)? mem[146] : 
                        (N82)? mem[208] : 
                        (N84)? mem[270] : 
                        (N86)? mem[332] : 
                        (N88)? mem[394] : 
                        (N90)? mem[456] : 
                        (N92)? mem[518] : 
                        (N94)? mem[580] : 
                        (N96)? mem[642] : 
                        (N98)? mem[704] : 
                        (N100)? mem[766] : 
                        (N102)? mem[828] : 
                        (N104)? mem[890] : 
                        (N106)? mem[952] : 
                        (N108)? mem[1014] : 
                        (N110)? mem[1076] : 
                        (N112)? mem[1138] : 
                        (N114)? mem[1200] : 
                        (N116)? mem[1262] : 
                        (N118)? mem[1324] : 
                        (N120)? mem[1386] : 
                        (N122)? mem[1448] : 
                        (N124)? mem[1510] : 
                        (N126)? mem[1572] : 
                        (N128)? mem[1634] : 
                        (N130)? mem[1696] : 
                        (N132)? mem[1758] : 
                        (N134)? mem[1820] : 
                        (N136)? mem[1882] : 
                        (N138)? mem[1944] : 
                        (N77)? mem[2006] : 
                        (N79)? mem[2068] : 
                        (N81)? mem[2130] : 
                        (N83)? mem[2192] : 
                        (N85)? mem[2254] : 
                        (N87)? mem[2316] : 
                        (N89)? mem[2378] : 
                        (N91)? mem[2440] : 
                        (N93)? mem[2502] : 
                        (N95)? mem[2564] : 
                        (N97)? mem[2626] : 
                        (N99)? mem[2688] : 
                        (N101)? mem[2750] : 
                        (N103)? mem[2812] : 
                        (N105)? mem[2874] : 
                        (N107)? mem[2936] : 
                        (N109)? mem[2998] : 
                        (N111)? mem[3060] : 
                        (N113)? mem[3122] : 
                        (N115)? mem[3184] : 
                        (N117)? mem[3246] : 
                        (N119)? mem[3308] : 
                        (N121)? mem[3370] : 
                        (N123)? mem[3432] : 
                        (N125)? mem[3494] : 
                        (N127)? mem[3556] : 
                        (N129)? mem[3618] : 
                        (N131)? mem[3680] : 
                        (N133)? mem[3742] : 
                        (N135)? mem[3804] : 
                        (N137)? mem[3866] : 
                        (N139)? mem[3928] : 1'b0;
  assign r_data_o[21] = (N76)? mem[21] : 
                        (N78)? mem[83] : 
                        (N80)? mem[145] : 
                        (N82)? mem[207] : 
                        (N84)? mem[269] : 
                        (N86)? mem[331] : 
                        (N88)? mem[393] : 
                        (N90)? mem[455] : 
                        (N92)? mem[517] : 
                        (N94)? mem[579] : 
                        (N96)? mem[641] : 
                        (N98)? mem[703] : 
                        (N100)? mem[765] : 
                        (N102)? mem[827] : 
                        (N104)? mem[889] : 
                        (N106)? mem[951] : 
                        (N108)? mem[1013] : 
                        (N110)? mem[1075] : 
                        (N112)? mem[1137] : 
                        (N114)? mem[1199] : 
                        (N116)? mem[1261] : 
                        (N118)? mem[1323] : 
                        (N120)? mem[1385] : 
                        (N122)? mem[1447] : 
                        (N124)? mem[1509] : 
                        (N126)? mem[1571] : 
                        (N128)? mem[1633] : 
                        (N130)? mem[1695] : 
                        (N132)? mem[1757] : 
                        (N134)? mem[1819] : 
                        (N136)? mem[1881] : 
                        (N138)? mem[1943] : 
                        (N77)? mem[2005] : 
                        (N79)? mem[2067] : 
                        (N81)? mem[2129] : 
                        (N83)? mem[2191] : 
                        (N85)? mem[2253] : 
                        (N87)? mem[2315] : 
                        (N89)? mem[2377] : 
                        (N91)? mem[2439] : 
                        (N93)? mem[2501] : 
                        (N95)? mem[2563] : 
                        (N97)? mem[2625] : 
                        (N99)? mem[2687] : 
                        (N101)? mem[2749] : 
                        (N103)? mem[2811] : 
                        (N105)? mem[2873] : 
                        (N107)? mem[2935] : 
                        (N109)? mem[2997] : 
                        (N111)? mem[3059] : 
                        (N113)? mem[3121] : 
                        (N115)? mem[3183] : 
                        (N117)? mem[3245] : 
                        (N119)? mem[3307] : 
                        (N121)? mem[3369] : 
                        (N123)? mem[3431] : 
                        (N125)? mem[3493] : 
                        (N127)? mem[3555] : 
                        (N129)? mem[3617] : 
                        (N131)? mem[3679] : 
                        (N133)? mem[3741] : 
                        (N135)? mem[3803] : 
                        (N137)? mem[3865] : 
                        (N139)? mem[3927] : 1'b0;
  assign r_data_o[20] = (N76)? mem[20] : 
                        (N78)? mem[82] : 
                        (N80)? mem[144] : 
                        (N82)? mem[206] : 
                        (N84)? mem[268] : 
                        (N86)? mem[330] : 
                        (N88)? mem[392] : 
                        (N90)? mem[454] : 
                        (N92)? mem[516] : 
                        (N94)? mem[578] : 
                        (N96)? mem[640] : 
                        (N98)? mem[702] : 
                        (N100)? mem[764] : 
                        (N102)? mem[826] : 
                        (N104)? mem[888] : 
                        (N106)? mem[950] : 
                        (N108)? mem[1012] : 
                        (N110)? mem[1074] : 
                        (N112)? mem[1136] : 
                        (N114)? mem[1198] : 
                        (N116)? mem[1260] : 
                        (N118)? mem[1322] : 
                        (N120)? mem[1384] : 
                        (N122)? mem[1446] : 
                        (N124)? mem[1508] : 
                        (N126)? mem[1570] : 
                        (N128)? mem[1632] : 
                        (N130)? mem[1694] : 
                        (N132)? mem[1756] : 
                        (N134)? mem[1818] : 
                        (N136)? mem[1880] : 
                        (N138)? mem[1942] : 
                        (N77)? mem[2004] : 
                        (N79)? mem[2066] : 
                        (N81)? mem[2128] : 
                        (N83)? mem[2190] : 
                        (N85)? mem[2252] : 
                        (N87)? mem[2314] : 
                        (N89)? mem[2376] : 
                        (N91)? mem[2438] : 
                        (N93)? mem[2500] : 
                        (N95)? mem[2562] : 
                        (N97)? mem[2624] : 
                        (N99)? mem[2686] : 
                        (N101)? mem[2748] : 
                        (N103)? mem[2810] : 
                        (N105)? mem[2872] : 
                        (N107)? mem[2934] : 
                        (N109)? mem[2996] : 
                        (N111)? mem[3058] : 
                        (N113)? mem[3120] : 
                        (N115)? mem[3182] : 
                        (N117)? mem[3244] : 
                        (N119)? mem[3306] : 
                        (N121)? mem[3368] : 
                        (N123)? mem[3430] : 
                        (N125)? mem[3492] : 
                        (N127)? mem[3554] : 
                        (N129)? mem[3616] : 
                        (N131)? mem[3678] : 
                        (N133)? mem[3740] : 
                        (N135)? mem[3802] : 
                        (N137)? mem[3864] : 
                        (N139)? mem[3926] : 1'b0;
  assign r_data_o[19] = (N76)? mem[19] : 
                        (N78)? mem[81] : 
                        (N80)? mem[143] : 
                        (N82)? mem[205] : 
                        (N84)? mem[267] : 
                        (N86)? mem[329] : 
                        (N88)? mem[391] : 
                        (N90)? mem[453] : 
                        (N92)? mem[515] : 
                        (N94)? mem[577] : 
                        (N96)? mem[639] : 
                        (N98)? mem[701] : 
                        (N100)? mem[763] : 
                        (N102)? mem[825] : 
                        (N104)? mem[887] : 
                        (N106)? mem[949] : 
                        (N108)? mem[1011] : 
                        (N110)? mem[1073] : 
                        (N112)? mem[1135] : 
                        (N114)? mem[1197] : 
                        (N116)? mem[1259] : 
                        (N118)? mem[1321] : 
                        (N120)? mem[1383] : 
                        (N122)? mem[1445] : 
                        (N124)? mem[1507] : 
                        (N126)? mem[1569] : 
                        (N128)? mem[1631] : 
                        (N130)? mem[1693] : 
                        (N132)? mem[1755] : 
                        (N134)? mem[1817] : 
                        (N136)? mem[1879] : 
                        (N138)? mem[1941] : 
                        (N77)? mem[2003] : 
                        (N79)? mem[2065] : 
                        (N81)? mem[2127] : 
                        (N83)? mem[2189] : 
                        (N85)? mem[2251] : 
                        (N87)? mem[2313] : 
                        (N89)? mem[2375] : 
                        (N91)? mem[2437] : 
                        (N93)? mem[2499] : 
                        (N95)? mem[2561] : 
                        (N97)? mem[2623] : 
                        (N99)? mem[2685] : 
                        (N101)? mem[2747] : 
                        (N103)? mem[2809] : 
                        (N105)? mem[2871] : 
                        (N107)? mem[2933] : 
                        (N109)? mem[2995] : 
                        (N111)? mem[3057] : 
                        (N113)? mem[3119] : 
                        (N115)? mem[3181] : 
                        (N117)? mem[3243] : 
                        (N119)? mem[3305] : 
                        (N121)? mem[3367] : 
                        (N123)? mem[3429] : 
                        (N125)? mem[3491] : 
                        (N127)? mem[3553] : 
                        (N129)? mem[3615] : 
                        (N131)? mem[3677] : 
                        (N133)? mem[3739] : 
                        (N135)? mem[3801] : 
                        (N137)? mem[3863] : 
                        (N139)? mem[3925] : 1'b0;
  assign r_data_o[18] = (N76)? mem[18] : 
                        (N78)? mem[80] : 
                        (N80)? mem[142] : 
                        (N82)? mem[204] : 
                        (N84)? mem[266] : 
                        (N86)? mem[328] : 
                        (N88)? mem[390] : 
                        (N90)? mem[452] : 
                        (N92)? mem[514] : 
                        (N94)? mem[576] : 
                        (N96)? mem[638] : 
                        (N98)? mem[700] : 
                        (N100)? mem[762] : 
                        (N102)? mem[824] : 
                        (N104)? mem[886] : 
                        (N106)? mem[948] : 
                        (N108)? mem[1010] : 
                        (N110)? mem[1072] : 
                        (N112)? mem[1134] : 
                        (N114)? mem[1196] : 
                        (N116)? mem[1258] : 
                        (N118)? mem[1320] : 
                        (N120)? mem[1382] : 
                        (N122)? mem[1444] : 
                        (N124)? mem[1506] : 
                        (N126)? mem[1568] : 
                        (N128)? mem[1630] : 
                        (N130)? mem[1692] : 
                        (N132)? mem[1754] : 
                        (N134)? mem[1816] : 
                        (N136)? mem[1878] : 
                        (N138)? mem[1940] : 
                        (N77)? mem[2002] : 
                        (N79)? mem[2064] : 
                        (N81)? mem[2126] : 
                        (N83)? mem[2188] : 
                        (N85)? mem[2250] : 
                        (N87)? mem[2312] : 
                        (N89)? mem[2374] : 
                        (N91)? mem[2436] : 
                        (N93)? mem[2498] : 
                        (N95)? mem[2560] : 
                        (N97)? mem[2622] : 
                        (N99)? mem[2684] : 
                        (N101)? mem[2746] : 
                        (N103)? mem[2808] : 
                        (N105)? mem[2870] : 
                        (N107)? mem[2932] : 
                        (N109)? mem[2994] : 
                        (N111)? mem[3056] : 
                        (N113)? mem[3118] : 
                        (N115)? mem[3180] : 
                        (N117)? mem[3242] : 
                        (N119)? mem[3304] : 
                        (N121)? mem[3366] : 
                        (N123)? mem[3428] : 
                        (N125)? mem[3490] : 
                        (N127)? mem[3552] : 
                        (N129)? mem[3614] : 
                        (N131)? mem[3676] : 
                        (N133)? mem[3738] : 
                        (N135)? mem[3800] : 
                        (N137)? mem[3862] : 
                        (N139)? mem[3924] : 1'b0;
  assign r_data_o[17] = (N76)? mem[17] : 
                        (N78)? mem[79] : 
                        (N80)? mem[141] : 
                        (N82)? mem[203] : 
                        (N84)? mem[265] : 
                        (N86)? mem[327] : 
                        (N88)? mem[389] : 
                        (N90)? mem[451] : 
                        (N92)? mem[513] : 
                        (N94)? mem[575] : 
                        (N96)? mem[637] : 
                        (N98)? mem[699] : 
                        (N100)? mem[761] : 
                        (N102)? mem[823] : 
                        (N104)? mem[885] : 
                        (N106)? mem[947] : 
                        (N108)? mem[1009] : 
                        (N110)? mem[1071] : 
                        (N112)? mem[1133] : 
                        (N114)? mem[1195] : 
                        (N116)? mem[1257] : 
                        (N118)? mem[1319] : 
                        (N120)? mem[1381] : 
                        (N122)? mem[1443] : 
                        (N124)? mem[1505] : 
                        (N126)? mem[1567] : 
                        (N128)? mem[1629] : 
                        (N130)? mem[1691] : 
                        (N132)? mem[1753] : 
                        (N134)? mem[1815] : 
                        (N136)? mem[1877] : 
                        (N138)? mem[1939] : 
                        (N77)? mem[2001] : 
                        (N79)? mem[2063] : 
                        (N81)? mem[2125] : 
                        (N83)? mem[2187] : 
                        (N85)? mem[2249] : 
                        (N87)? mem[2311] : 
                        (N89)? mem[2373] : 
                        (N91)? mem[2435] : 
                        (N93)? mem[2497] : 
                        (N95)? mem[2559] : 
                        (N97)? mem[2621] : 
                        (N99)? mem[2683] : 
                        (N101)? mem[2745] : 
                        (N103)? mem[2807] : 
                        (N105)? mem[2869] : 
                        (N107)? mem[2931] : 
                        (N109)? mem[2993] : 
                        (N111)? mem[3055] : 
                        (N113)? mem[3117] : 
                        (N115)? mem[3179] : 
                        (N117)? mem[3241] : 
                        (N119)? mem[3303] : 
                        (N121)? mem[3365] : 
                        (N123)? mem[3427] : 
                        (N125)? mem[3489] : 
                        (N127)? mem[3551] : 
                        (N129)? mem[3613] : 
                        (N131)? mem[3675] : 
                        (N133)? mem[3737] : 
                        (N135)? mem[3799] : 
                        (N137)? mem[3861] : 
                        (N139)? mem[3923] : 1'b0;
  assign r_data_o[16] = (N76)? mem[16] : 
                        (N78)? mem[78] : 
                        (N80)? mem[140] : 
                        (N82)? mem[202] : 
                        (N84)? mem[264] : 
                        (N86)? mem[326] : 
                        (N88)? mem[388] : 
                        (N90)? mem[450] : 
                        (N92)? mem[512] : 
                        (N94)? mem[574] : 
                        (N96)? mem[636] : 
                        (N98)? mem[698] : 
                        (N100)? mem[760] : 
                        (N102)? mem[822] : 
                        (N104)? mem[884] : 
                        (N106)? mem[946] : 
                        (N108)? mem[1008] : 
                        (N110)? mem[1070] : 
                        (N112)? mem[1132] : 
                        (N114)? mem[1194] : 
                        (N116)? mem[1256] : 
                        (N118)? mem[1318] : 
                        (N120)? mem[1380] : 
                        (N122)? mem[1442] : 
                        (N124)? mem[1504] : 
                        (N126)? mem[1566] : 
                        (N128)? mem[1628] : 
                        (N130)? mem[1690] : 
                        (N132)? mem[1752] : 
                        (N134)? mem[1814] : 
                        (N136)? mem[1876] : 
                        (N138)? mem[1938] : 
                        (N77)? mem[2000] : 
                        (N79)? mem[2062] : 
                        (N81)? mem[2124] : 
                        (N83)? mem[2186] : 
                        (N85)? mem[2248] : 
                        (N87)? mem[2310] : 
                        (N89)? mem[2372] : 
                        (N91)? mem[2434] : 
                        (N93)? mem[2496] : 
                        (N95)? mem[2558] : 
                        (N97)? mem[2620] : 
                        (N99)? mem[2682] : 
                        (N101)? mem[2744] : 
                        (N103)? mem[2806] : 
                        (N105)? mem[2868] : 
                        (N107)? mem[2930] : 
                        (N109)? mem[2992] : 
                        (N111)? mem[3054] : 
                        (N113)? mem[3116] : 
                        (N115)? mem[3178] : 
                        (N117)? mem[3240] : 
                        (N119)? mem[3302] : 
                        (N121)? mem[3364] : 
                        (N123)? mem[3426] : 
                        (N125)? mem[3488] : 
                        (N127)? mem[3550] : 
                        (N129)? mem[3612] : 
                        (N131)? mem[3674] : 
                        (N133)? mem[3736] : 
                        (N135)? mem[3798] : 
                        (N137)? mem[3860] : 
                        (N139)? mem[3922] : 1'b0;
  assign r_data_o[15] = (N76)? mem[15] : 
                        (N78)? mem[77] : 
                        (N80)? mem[139] : 
                        (N82)? mem[201] : 
                        (N84)? mem[263] : 
                        (N86)? mem[325] : 
                        (N88)? mem[387] : 
                        (N90)? mem[449] : 
                        (N92)? mem[511] : 
                        (N94)? mem[573] : 
                        (N96)? mem[635] : 
                        (N98)? mem[697] : 
                        (N100)? mem[759] : 
                        (N102)? mem[821] : 
                        (N104)? mem[883] : 
                        (N106)? mem[945] : 
                        (N108)? mem[1007] : 
                        (N110)? mem[1069] : 
                        (N112)? mem[1131] : 
                        (N114)? mem[1193] : 
                        (N116)? mem[1255] : 
                        (N118)? mem[1317] : 
                        (N120)? mem[1379] : 
                        (N122)? mem[1441] : 
                        (N124)? mem[1503] : 
                        (N126)? mem[1565] : 
                        (N128)? mem[1627] : 
                        (N130)? mem[1689] : 
                        (N132)? mem[1751] : 
                        (N134)? mem[1813] : 
                        (N136)? mem[1875] : 
                        (N138)? mem[1937] : 
                        (N77)? mem[1999] : 
                        (N79)? mem[2061] : 
                        (N81)? mem[2123] : 
                        (N83)? mem[2185] : 
                        (N85)? mem[2247] : 
                        (N87)? mem[2309] : 
                        (N89)? mem[2371] : 
                        (N91)? mem[2433] : 
                        (N93)? mem[2495] : 
                        (N95)? mem[2557] : 
                        (N97)? mem[2619] : 
                        (N99)? mem[2681] : 
                        (N101)? mem[2743] : 
                        (N103)? mem[2805] : 
                        (N105)? mem[2867] : 
                        (N107)? mem[2929] : 
                        (N109)? mem[2991] : 
                        (N111)? mem[3053] : 
                        (N113)? mem[3115] : 
                        (N115)? mem[3177] : 
                        (N117)? mem[3239] : 
                        (N119)? mem[3301] : 
                        (N121)? mem[3363] : 
                        (N123)? mem[3425] : 
                        (N125)? mem[3487] : 
                        (N127)? mem[3549] : 
                        (N129)? mem[3611] : 
                        (N131)? mem[3673] : 
                        (N133)? mem[3735] : 
                        (N135)? mem[3797] : 
                        (N137)? mem[3859] : 
                        (N139)? mem[3921] : 1'b0;
  assign r_data_o[14] = (N76)? mem[14] : 
                        (N78)? mem[76] : 
                        (N80)? mem[138] : 
                        (N82)? mem[200] : 
                        (N84)? mem[262] : 
                        (N86)? mem[324] : 
                        (N88)? mem[386] : 
                        (N90)? mem[448] : 
                        (N92)? mem[510] : 
                        (N94)? mem[572] : 
                        (N96)? mem[634] : 
                        (N98)? mem[696] : 
                        (N100)? mem[758] : 
                        (N102)? mem[820] : 
                        (N104)? mem[882] : 
                        (N106)? mem[944] : 
                        (N108)? mem[1006] : 
                        (N110)? mem[1068] : 
                        (N112)? mem[1130] : 
                        (N114)? mem[1192] : 
                        (N116)? mem[1254] : 
                        (N118)? mem[1316] : 
                        (N120)? mem[1378] : 
                        (N122)? mem[1440] : 
                        (N124)? mem[1502] : 
                        (N126)? mem[1564] : 
                        (N128)? mem[1626] : 
                        (N130)? mem[1688] : 
                        (N132)? mem[1750] : 
                        (N134)? mem[1812] : 
                        (N136)? mem[1874] : 
                        (N138)? mem[1936] : 
                        (N77)? mem[1998] : 
                        (N79)? mem[2060] : 
                        (N81)? mem[2122] : 
                        (N83)? mem[2184] : 
                        (N85)? mem[2246] : 
                        (N87)? mem[2308] : 
                        (N89)? mem[2370] : 
                        (N91)? mem[2432] : 
                        (N93)? mem[2494] : 
                        (N95)? mem[2556] : 
                        (N97)? mem[2618] : 
                        (N99)? mem[2680] : 
                        (N101)? mem[2742] : 
                        (N103)? mem[2804] : 
                        (N105)? mem[2866] : 
                        (N107)? mem[2928] : 
                        (N109)? mem[2990] : 
                        (N111)? mem[3052] : 
                        (N113)? mem[3114] : 
                        (N115)? mem[3176] : 
                        (N117)? mem[3238] : 
                        (N119)? mem[3300] : 
                        (N121)? mem[3362] : 
                        (N123)? mem[3424] : 
                        (N125)? mem[3486] : 
                        (N127)? mem[3548] : 
                        (N129)? mem[3610] : 
                        (N131)? mem[3672] : 
                        (N133)? mem[3734] : 
                        (N135)? mem[3796] : 
                        (N137)? mem[3858] : 
                        (N139)? mem[3920] : 1'b0;
  assign r_data_o[13] = (N76)? mem[13] : 
                        (N78)? mem[75] : 
                        (N80)? mem[137] : 
                        (N82)? mem[199] : 
                        (N84)? mem[261] : 
                        (N86)? mem[323] : 
                        (N88)? mem[385] : 
                        (N90)? mem[447] : 
                        (N92)? mem[509] : 
                        (N94)? mem[571] : 
                        (N96)? mem[633] : 
                        (N98)? mem[695] : 
                        (N100)? mem[757] : 
                        (N102)? mem[819] : 
                        (N104)? mem[881] : 
                        (N106)? mem[943] : 
                        (N108)? mem[1005] : 
                        (N110)? mem[1067] : 
                        (N112)? mem[1129] : 
                        (N114)? mem[1191] : 
                        (N116)? mem[1253] : 
                        (N118)? mem[1315] : 
                        (N120)? mem[1377] : 
                        (N122)? mem[1439] : 
                        (N124)? mem[1501] : 
                        (N126)? mem[1563] : 
                        (N128)? mem[1625] : 
                        (N130)? mem[1687] : 
                        (N132)? mem[1749] : 
                        (N134)? mem[1811] : 
                        (N136)? mem[1873] : 
                        (N138)? mem[1935] : 
                        (N77)? mem[1997] : 
                        (N79)? mem[2059] : 
                        (N81)? mem[2121] : 
                        (N83)? mem[2183] : 
                        (N85)? mem[2245] : 
                        (N87)? mem[2307] : 
                        (N89)? mem[2369] : 
                        (N91)? mem[2431] : 
                        (N93)? mem[2493] : 
                        (N95)? mem[2555] : 
                        (N97)? mem[2617] : 
                        (N99)? mem[2679] : 
                        (N101)? mem[2741] : 
                        (N103)? mem[2803] : 
                        (N105)? mem[2865] : 
                        (N107)? mem[2927] : 
                        (N109)? mem[2989] : 
                        (N111)? mem[3051] : 
                        (N113)? mem[3113] : 
                        (N115)? mem[3175] : 
                        (N117)? mem[3237] : 
                        (N119)? mem[3299] : 
                        (N121)? mem[3361] : 
                        (N123)? mem[3423] : 
                        (N125)? mem[3485] : 
                        (N127)? mem[3547] : 
                        (N129)? mem[3609] : 
                        (N131)? mem[3671] : 
                        (N133)? mem[3733] : 
                        (N135)? mem[3795] : 
                        (N137)? mem[3857] : 
                        (N139)? mem[3919] : 1'b0;
  assign r_data_o[12] = (N76)? mem[12] : 
                        (N78)? mem[74] : 
                        (N80)? mem[136] : 
                        (N82)? mem[198] : 
                        (N84)? mem[260] : 
                        (N86)? mem[322] : 
                        (N88)? mem[384] : 
                        (N90)? mem[446] : 
                        (N92)? mem[508] : 
                        (N94)? mem[570] : 
                        (N96)? mem[632] : 
                        (N98)? mem[694] : 
                        (N100)? mem[756] : 
                        (N102)? mem[818] : 
                        (N104)? mem[880] : 
                        (N106)? mem[942] : 
                        (N108)? mem[1004] : 
                        (N110)? mem[1066] : 
                        (N112)? mem[1128] : 
                        (N114)? mem[1190] : 
                        (N116)? mem[1252] : 
                        (N118)? mem[1314] : 
                        (N120)? mem[1376] : 
                        (N122)? mem[1438] : 
                        (N124)? mem[1500] : 
                        (N126)? mem[1562] : 
                        (N128)? mem[1624] : 
                        (N130)? mem[1686] : 
                        (N132)? mem[1748] : 
                        (N134)? mem[1810] : 
                        (N136)? mem[1872] : 
                        (N138)? mem[1934] : 
                        (N77)? mem[1996] : 
                        (N79)? mem[2058] : 
                        (N81)? mem[2120] : 
                        (N83)? mem[2182] : 
                        (N85)? mem[2244] : 
                        (N87)? mem[2306] : 
                        (N89)? mem[2368] : 
                        (N91)? mem[2430] : 
                        (N93)? mem[2492] : 
                        (N95)? mem[2554] : 
                        (N97)? mem[2616] : 
                        (N99)? mem[2678] : 
                        (N101)? mem[2740] : 
                        (N103)? mem[2802] : 
                        (N105)? mem[2864] : 
                        (N107)? mem[2926] : 
                        (N109)? mem[2988] : 
                        (N111)? mem[3050] : 
                        (N113)? mem[3112] : 
                        (N115)? mem[3174] : 
                        (N117)? mem[3236] : 
                        (N119)? mem[3298] : 
                        (N121)? mem[3360] : 
                        (N123)? mem[3422] : 
                        (N125)? mem[3484] : 
                        (N127)? mem[3546] : 
                        (N129)? mem[3608] : 
                        (N131)? mem[3670] : 
                        (N133)? mem[3732] : 
                        (N135)? mem[3794] : 
                        (N137)? mem[3856] : 
                        (N139)? mem[3918] : 1'b0;
  assign r_data_o[11] = (N76)? mem[11] : 
                        (N78)? mem[73] : 
                        (N80)? mem[135] : 
                        (N82)? mem[197] : 
                        (N84)? mem[259] : 
                        (N86)? mem[321] : 
                        (N88)? mem[383] : 
                        (N90)? mem[445] : 
                        (N92)? mem[507] : 
                        (N94)? mem[569] : 
                        (N96)? mem[631] : 
                        (N98)? mem[693] : 
                        (N100)? mem[755] : 
                        (N102)? mem[817] : 
                        (N104)? mem[879] : 
                        (N106)? mem[941] : 
                        (N108)? mem[1003] : 
                        (N110)? mem[1065] : 
                        (N112)? mem[1127] : 
                        (N114)? mem[1189] : 
                        (N116)? mem[1251] : 
                        (N118)? mem[1313] : 
                        (N120)? mem[1375] : 
                        (N122)? mem[1437] : 
                        (N124)? mem[1499] : 
                        (N126)? mem[1561] : 
                        (N128)? mem[1623] : 
                        (N130)? mem[1685] : 
                        (N132)? mem[1747] : 
                        (N134)? mem[1809] : 
                        (N136)? mem[1871] : 
                        (N138)? mem[1933] : 
                        (N77)? mem[1995] : 
                        (N79)? mem[2057] : 
                        (N81)? mem[2119] : 
                        (N83)? mem[2181] : 
                        (N85)? mem[2243] : 
                        (N87)? mem[2305] : 
                        (N89)? mem[2367] : 
                        (N91)? mem[2429] : 
                        (N93)? mem[2491] : 
                        (N95)? mem[2553] : 
                        (N97)? mem[2615] : 
                        (N99)? mem[2677] : 
                        (N101)? mem[2739] : 
                        (N103)? mem[2801] : 
                        (N105)? mem[2863] : 
                        (N107)? mem[2925] : 
                        (N109)? mem[2987] : 
                        (N111)? mem[3049] : 
                        (N113)? mem[3111] : 
                        (N115)? mem[3173] : 
                        (N117)? mem[3235] : 
                        (N119)? mem[3297] : 
                        (N121)? mem[3359] : 
                        (N123)? mem[3421] : 
                        (N125)? mem[3483] : 
                        (N127)? mem[3545] : 
                        (N129)? mem[3607] : 
                        (N131)? mem[3669] : 
                        (N133)? mem[3731] : 
                        (N135)? mem[3793] : 
                        (N137)? mem[3855] : 
                        (N139)? mem[3917] : 1'b0;
  assign r_data_o[10] = (N76)? mem[10] : 
                        (N78)? mem[72] : 
                        (N80)? mem[134] : 
                        (N82)? mem[196] : 
                        (N84)? mem[258] : 
                        (N86)? mem[320] : 
                        (N88)? mem[382] : 
                        (N90)? mem[444] : 
                        (N92)? mem[506] : 
                        (N94)? mem[568] : 
                        (N96)? mem[630] : 
                        (N98)? mem[692] : 
                        (N100)? mem[754] : 
                        (N102)? mem[816] : 
                        (N104)? mem[878] : 
                        (N106)? mem[940] : 
                        (N108)? mem[1002] : 
                        (N110)? mem[1064] : 
                        (N112)? mem[1126] : 
                        (N114)? mem[1188] : 
                        (N116)? mem[1250] : 
                        (N118)? mem[1312] : 
                        (N120)? mem[1374] : 
                        (N122)? mem[1436] : 
                        (N124)? mem[1498] : 
                        (N126)? mem[1560] : 
                        (N128)? mem[1622] : 
                        (N130)? mem[1684] : 
                        (N132)? mem[1746] : 
                        (N134)? mem[1808] : 
                        (N136)? mem[1870] : 
                        (N138)? mem[1932] : 
                        (N77)? mem[1994] : 
                        (N79)? mem[2056] : 
                        (N81)? mem[2118] : 
                        (N83)? mem[2180] : 
                        (N85)? mem[2242] : 
                        (N87)? mem[2304] : 
                        (N89)? mem[2366] : 
                        (N91)? mem[2428] : 
                        (N93)? mem[2490] : 
                        (N95)? mem[2552] : 
                        (N97)? mem[2614] : 
                        (N99)? mem[2676] : 
                        (N101)? mem[2738] : 
                        (N103)? mem[2800] : 
                        (N105)? mem[2862] : 
                        (N107)? mem[2924] : 
                        (N109)? mem[2986] : 
                        (N111)? mem[3048] : 
                        (N113)? mem[3110] : 
                        (N115)? mem[3172] : 
                        (N117)? mem[3234] : 
                        (N119)? mem[3296] : 
                        (N121)? mem[3358] : 
                        (N123)? mem[3420] : 
                        (N125)? mem[3482] : 
                        (N127)? mem[3544] : 
                        (N129)? mem[3606] : 
                        (N131)? mem[3668] : 
                        (N133)? mem[3730] : 
                        (N135)? mem[3792] : 
                        (N137)? mem[3854] : 
                        (N139)? mem[3916] : 1'b0;
  assign r_data_o[9] = (N76)? mem[9] : 
                       (N78)? mem[71] : 
                       (N80)? mem[133] : 
                       (N82)? mem[195] : 
                       (N84)? mem[257] : 
                       (N86)? mem[319] : 
                       (N88)? mem[381] : 
                       (N90)? mem[443] : 
                       (N92)? mem[505] : 
                       (N94)? mem[567] : 
                       (N96)? mem[629] : 
                       (N98)? mem[691] : 
                       (N100)? mem[753] : 
                       (N102)? mem[815] : 
                       (N104)? mem[877] : 
                       (N106)? mem[939] : 
                       (N108)? mem[1001] : 
                       (N110)? mem[1063] : 
                       (N112)? mem[1125] : 
                       (N114)? mem[1187] : 
                       (N116)? mem[1249] : 
                       (N118)? mem[1311] : 
                       (N120)? mem[1373] : 
                       (N122)? mem[1435] : 
                       (N124)? mem[1497] : 
                       (N126)? mem[1559] : 
                       (N128)? mem[1621] : 
                       (N130)? mem[1683] : 
                       (N132)? mem[1745] : 
                       (N134)? mem[1807] : 
                       (N136)? mem[1869] : 
                       (N138)? mem[1931] : 
                       (N77)? mem[1993] : 
                       (N79)? mem[2055] : 
                       (N81)? mem[2117] : 
                       (N83)? mem[2179] : 
                       (N85)? mem[2241] : 
                       (N87)? mem[2303] : 
                       (N89)? mem[2365] : 
                       (N91)? mem[2427] : 
                       (N93)? mem[2489] : 
                       (N95)? mem[2551] : 
                       (N97)? mem[2613] : 
                       (N99)? mem[2675] : 
                       (N101)? mem[2737] : 
                       (N103)? mem[2799] : 
                       (N105)? mem[2861] : 
                       (N107)? mem[2923] : 
                       (N109)? mem[2985] : 
                       (N111)? mem[3047] : 
                       (N113)? mem[3109] : 
                       (N115)? mem[3171] : 
                       (N117)? mem[3233] : 
                       (N119)? mem[3295] : 
                       (N121)? mem[3357] : 
                       (N123)? mem[3419] : 
                       (N125)? mem[3481] : 
                       (N127)? mem[3543] : 
                       (N129)? mem[3605] : 
                       (N131)? mem[3667] : 
                       (N133)? mem[3729] : 
                       (N135)? mem[3791] : 
                       (N137)? mem[3853] : 
                       (N139)? mem[3915] : 1'b0;
  assign r_data_o[8] = (N76)? mem[8] : 
                       (N78)? mem[70] : 
                       (N80)? mem[132] : 
                       (N82)? mem[194] : 
                       (N84)? mem[256] : 
                       (N86)? mem[318] : 
                       (N88)? mem[380] : 
                       (N90)? mem[442] : 
                       (N92)? mem[504] : 
                       (N94)? mem[566] : 
                       (N96)? mem[628] : 
                       (N98)? mem[690] : 
                       (N100)? mem[752] : 
                       (N102)? mem[814] : 
                       (N104)? mem[876] : 
                       (N106)? mem[938] : 
                       (N108)? mem[1000] : 
                       (N110)? mem[1062] : 
                       (N112)? mem[1124] : 
                       (N114)? mem[1186] : 
                       (N116)? mem[1248] : 
                       (N118)? mem[1310] : 
                       (N120)? mem[1372] : 
                       (N122)? mem[1434] : 
                       (N124)? mem[1496] : 
                       (N126)? mem[1558] : 
                       (N128)? mem[1620] : 
                       (N130)? mem[1682] : 
                       (N132)? mem[1744] : 
                       (N134)? mem[1806] : 
                       (N136)? mem[1868] : 
                       (N138)? mem[1930] : 
                       (N77)? mem[1992] : 
                       (N79)? mem[2054] : 
                       (N81)? mem[2116] : 
                       (N83)? mem[2178] : 
                       (N85)? mem[2240] : 
                       (N87)? mem[2302] : 
                       (N89)? mem[2364] : 
                       (N91)? mem[2426] : 
                       (N93)? mem[2488] : 
                       (N95)? mem[2550] : 
                       (N97)? mem[2612] : 
                       (N99)? mem[2674] : 
                       (N101)? mem[2736] : 
                       (N103)? mem[2798] : 
                       (N105)? mem[2860] : 
                       (N107)? mem[2922] : 
                       (N109)? mem[2984] : 
                       (N111)? mem[3046] : 
                       (N113)? mem[3108] : 
                       (N115)? mem[3170] : 
                       (N117)? mem[3232] : 
                       (N119)? mem[3294] : 
                       (N121)? mem[3356] : 
                       (N123)? mem[3418] : 
                       (N125)? mem[3480] : 
                       (N127)? mem[3542] : 
                       (N129)? mem[3604] : 
                       (N131)? mem[3666] : 
                       (N133)? mem[3728] : 
                       (N135)? mem[3790] : 
                       (N137)? mem[3852] : 
                       (N139)? mem[3914] : 1'b0;
  assign r_data_o[7] = (N76)? mem[7] : 
                       (N78)? mem[69] : 
                       (N80)? mem[131] : 
                       (N82)? mem[193] : 
                       (N84)? mem[255] : 
                       (N86)? mem[317] : 
                       (N88)? mem[379] : 
                       (N90)? mem[441] : 
                       (N92)? mem[503] : 
                       (N94)? mem[565] : 
                       (N96)? mem[627] : 
                       (N98)? mem[689] : 
                       (N100)? mem[751] : 
                       (N102)? mem[813] : 
                       (N104)? mem[875] : 
                       (N106)? mem[937] : 
                       (N108)? mem[999] : 
                       (N110)? mem[1061] : 
                       (N112)? mem[1123] : 
                       (N114)? mem[1185] : 
                       (N116)? mem[1247] : 
                       (N118)? mem[1309] : 
                       (N120)? mem[1371] : 
                       (N122)? mem[1433] : 
                       (N124)? mem[1495] : 
                       (N126)? mem[1557] : 
                       (N128)? mem[1619] : 
                       (N130)? mem[1681] : 
                       (N132)? mem[1743] : 
                       (N134)? mem[1805] : 
                       (N136)? mem[1867] : 
                       (N138)? mem[1929] : 
                       (N77)? mem[1991] : 
                       (N79)? mem[2053] : 
                       (N81)? mem[2115] : 
                       (N83)? mem[2177] : 
                       (N85)? mem[2239] : 
                       (N87)? mem[2301] : 
                       (N89)? mem[2363] : 
                       (N91)? mem[2425] : 
                       (N93)? mem[2487] : 
                       (N95)? mem[2549] : 
                       (N97)? mem[2611] : 
                       (N99)? mem[2673] : 
                       (N101)? mem[2735] : 
                       (N103)? mem[2797] : 
                       (N105)? mem[2859] : 
                       (N107)? mem[2921] : 
                       (N109)? mem[2983] : 
                       (N111)? mem[3045] : 
                       (N113)? mem[3107] : 
                       (N115)? mem[3169] : 
                       (N117)? mem[3231] : 
                       (N119)? mem[3293] : 
                       (N121)? mem[3355] : 
                       (N123)? mem[3417] : 
                       (N125)? mem[3479] : 
                       (N127)? mem[3541] : 
                       (N129)? mem[3603] : 
                       (N131)? mem[3665] : 
                       (N133)? mem[3727] : 
                       (N135)? mem[3789] : 
                       (N137)? mem[3851] : 
                       (N139)? mem[3913] : 1'b0;
  assign r_data_o[6] = (N76)? mem[6] : 
                       (N78)? mem[68] : 
                       (N80)? mem[130] : 
                       (N82)? mem[192] : 
                       (N84)? mem[254] : 
                       (N86)? mem[316] : 
                       (N88)? mem[378] : 
                       (N90)? mem[440] : 
                       (N92)? mem[502] : 
                       (N94)? mem[564] : 
                       (N96)? mem[626] : 
                       (N98)? mem[688] : 
                       (N100)? mem[750] : 
                       (N102)? mem[812] : 
                       (N104)? mem[874] : 
                       (N106)? mem[936] : 
                       (N108)? mem[998] : 
                       (N110)? mem[1060] : 
                       (N112)? mem[1122] : 
                       (N114)? mem[1184] : 
                       (N116)? mem[1246] : 
                       (N118)? mem[1308] : 
                       (N120)? mem[1370] : 
                       (N122)? mem[1432] : 
                       (N124)? mem[1494] : 
                       (N126)? mem[1556] : 
                       (N128)? mem[1618] : 
                       (N130)? mem[1680] : 
                       (N132)? mem[1742] : 
                       (N134)? mem[1804] : 
                       (N136)? mem[1866] : 
                       (N138)? mem[1928] : 
                       (N77)? mem[1990] : 
                       (N79)? mem[2052] : 
                       (N81)? mem[2114] : 
                       (N83)? mem[2176] : 
                       (N85)? mem[2238] : 
                       (N87)? mem[2300] : 
                       (N89)? mem[2362] : 
                       (N91)? mem[2424] : 
                       (N93)? mem[2486] : 
                       (N95)? mem[2548] : 
                       (N97)? mem[2610] : 
                       (N99)? mem[2672] : 
                       (N101)? mem[2734] : 
                       (N103)? mem[2796] : 
                       (N105)? mem[2858] : 
                       (N107)? mem[2920] : 
                       (N109)? mem[2982] : 
                       (N111)? mem[3044] : 
                       (N113)? mem[3106] : 
                       (N115)? mem[3168] : 
                       (N117)? mem[3230] : 
                       (N119)? mem[3292] : 
                       (N121)? mem[3354] : 
                       (N123)? mem[3416] : 
                       (N125)? mem[3478] : 
                       (N127)? mem[3540] : 
                       (N129)? mem[3602] : 
                       (N131)? mem[3664] : 
                       (N133)? mem[3726] : 
                       (N135)? mem[3788] : 
                       (N137)? mem[3850] : 
                       (N139)? mem[3912] : 1'b0;
  assign r_data_o[5] = (N76)? mem[5] : 
                       (N78)? mem[67] : 
                       (N80)? mem[129] : 
                       (N82)? mem[191] : 
                       (N84)? mem[253] : 
                       (N86)? mem[315] : 
                       (N88)? mem[377] : 
                       (N90)? mem[439] : 
                       (N92)? mem[501] : 
                       (N94)? mem[563] : 
                       (N96)? mem[625] : 
                       (N98)? mem[687] : 
                       (N100)? mem[749] : 
                       (N102)? mem[811] : 
                       (N104)? mem[873] : 
                       (N106)? mem[935] : 
                       (N108)? mem[997] : 
                       (N110)? mem[1059] : 
                       (N112)? mem[1121] : 
                       (N114)? mem[1183] : 
                       (N116)? mem[1245] : 
                       (N118)? mem[1307] : 
                       (N120)? mem[1369] : 
                       (N122)? mem[1431] : 
                       (N124)? mem[1493] : 
                       (N126)? mem[1555] : 
                       (N128)? mem[1617] : 
                       (N130)? mem[1679] : 
                       (N132)? mem[1741] : 
                       (N134)? mem[1803] : 
                       (N136)? mem[1865] : 
                       (N138)? mem[1927] : 
                       (N77)? mem[1989] : 
                       (N79)? mem[2051] : 
                       (N81)? mem[2113] : 
                       (N83)? mem[2175] : 
                       (N85)? mem[2237] : 
                       (N87)? mem[2299] : 
                       (N89)? mem[2361] : 
                       (N91)? mem[2423] : 
                       (N93)? mem[2485] : 
                       (N95)? mem[2547] : 
                       (N97)? mem[2609] : 
                       (N99)? mem[2671] : 
                       (N101)? mem[2733] : 
                       (N103)? mem[2795] : 
                       (N105)? mem[2857] : 
                       (N107)? mem[2919] : 
                       (N109)? mem[2981] : 
                       (N111)? mem[3043] : 
                       (N113)? mem[3105] : 
                       (N115)? mem[3167] : 
                       (N117)? mem[3229] : 
                       (N119)? mem[3291] : 
                       (N121)? mem[3353] : 
                       (N123)? mem[3415] : 
                       (N125)? mem[3477] : 
                       (N127)? mem[3539] : 
                       (N129)? mem[3601] : 
                       (N131)? mem[3663] : 
                       (N133)? mem[3725] : 
                       (N135)? mem[3787] : 
                       (N137)? mem[3849] : 
                       (N139)? mem[3911] : 1'b0;
  assign r_data_o[4] = (N76)? mem[4] : 
                       (N78)? mem[66] : 
                       (N80)? mem[128] : 
                       (N82)? mem[190] : 
                       (N84)? mem[252] : 
                       (N86)? mem[314] : 
                       (N88)? mem[376] : 
                       (N90)? mem[438] : 
                       (N92)? mem[500] : 
                       (N94)? mem[562] : 
                       (N96)? mem[624] : 
                       (N98)? mem[686] : 
                       (N100)? mem[748] : 
                       (N102)? mem[810] : 
                       (N104)? mem[872] : 
                       (N106)? mem[934] : 
                       (N108)? mem[996] : 
                       (N110)? mem[1058] : 
                       (N112)? mem[1120] : 
                       (N114)? mem[1182] : 
                       (N116)? mem[1244] : 
                       (N118)? mem[1306] : 
                       (N120)? mem[1368] : 
                       (N122)? mem[1430] : 
                       (N124)? mem[1492] : 
                       (N126)? mem[1554] : 
                       (N128)? mem[1616] : 
                       (N130)? mem[1678] : 
                       (N132)? mem[1740] : 
                       (N134)? mem[1802] : 
                       (N136)? mem[1864] : 
                       (N138)? mem[1926] : 
                       (N77)? mem[1988] : 
                       (N79)? mem[2050] : 
                       (N81)? mem[2112] : 
                       (N83)? mem[2174] : 
                       (N85)? mem[2236] : 
                       (N87)? mem[2298] : 
                       (N89)? mem[2360] : 
                       (N91)? mem[2422] : 
                       (N93)? mem[2484] : 
                       (N95)? mem[2546] : 
                       (N97)? mem[2608] : 
                       (N99)? mem[2670] : 
                       (N101)? mem[2732] : 
                       (N103)? mem[2794] : 
                       (N105)? mem[2856] : 
                       (N107)? mem[2918] : 
                       (N109)? mem[2980] : 
                       (N111)? mem[3042] : 
                       (N113)? mem[3104] : 
                       (N115)? mem[3166] : 
                       (N117)? mem[3228] : 
                       (N119)? mem[3290] : 
                       (N121)? mem[3352] : 
                       (N123)? mem[3414] : 
                       (N125)? mem[3476] : 
                       (N127)? mem[3538] : 
                       (N129)? mem[3600] : 
                       (N131)? mem[3662] : 
                       (N133)? mem[3724] : 
                       (N135)? mem[3786] : 
                       (N137)? mem[3848] : 
                       (N139)? mem[3910] : 1'b0;
  assign r_data_o[3] = (N76)? mem[3] : 
                       (N78)? mem[65] : 
                       (N80)? mem[127] : 
                       (N82)? mem[189] : 
                       (N84)? mem[251] : 
                       (N86)? mem[313] : 
                       (N88)? mem[375] : 
                       (N90)? mem[437] : 
                       (N92)? mem[499] : 
                       (N94)? mem[561] : 
                       (N96)? mem[623] : 
                       (N98)? mem[685] : 
                       (N100)? mem[747] : 
                       (N102)? mem[809] : 
                       (N104)? mem[871] : 
                       (N106)? mem[933] : 
                       (N108)? mem[995] : 
                       (N110)? mem[1057] : 
                       (N112)? mem[1119] : 
                       (N114)? mem[1181] : 
                       (N116)? mem[1243] : 
                       (N118)? mem[1305] : 
                       (N120)? mem[1367] : 
                       (N122)? mem[1429] : 
                       (N124)? mem[1491] : 
                       (N126)? mem[1553] : 
                       (N128)? mem[1615] : 
                       (N130)? mem[1677] : 
                       (N132)? mem[1739] : 
                       (N134)? mem[1801] : 
                       (N136)? mem[1863] : 
                       (N138)? mem[1925] : 
                       (N77)? mem[1987] : 
                       (N79)? mem[2049] : 
                       (N81)? mem[2111] : 
                       (N83)? mem[2173] : 
                       (N85)? mem[2235] : 
                       (N87)? mem[2297] : 
                       (N89)? mem[2359] : 
                       (N91)? mem[2421] : 
                       (N93)? mem[2483] : 
                       (N95)? mem[2545] : 
                       (N97)? mem[2607] : 
                       (N99)? mem[2669] : 
                       (N101)? mem[2731] : 
                       (N103)? mem[2793] : 
                       (N105)? mem[2855] : 
                       (N107)? mem[2917] : 
                       (N109)? mem[2979] : 
                       (N111)? mem[3041] : 
                       (N113)? mem[3103] : 
                       (N115)? mem[3165] : 
                       (N117)? mem[3227] : 
                       (N119)? mem[3289] : 
                       (N121)? mem[3351] : 
                       (N123)? mem[3413] : 
                       (N125)? mem[3475] : 
                       (N127)? mem[3537] : 
                       (N129)? mem[3599] : 
                       (N131)? mem[3661] : 
                       (N133)? mem[3723] : 
                       (N135)? mem[3785] : 
                       (N137)? mem[3847] : 
                       (N139)? mem[3909] : 1'b0;
  assign r_data_o[2] = (N76)? mem[2] : 
                       (N78)? mem[64] : 
                       (N80)? mem[126] : 
                       (N82)? mem[188] : 
                       (N84)? mem[250] : 
                       (N86)? mem[312] : 
                       (N88)? mem[374] : 
                       (N90)? mem[436] : 
                       (N92)? mem[498] : 
                       (N94)? mem[560] : 
                       (N96)? mem[622] : 
                       (N98)? mem[684] : 
                       (N100)? mem[746] : 
                       (N102)? mem[808] : 
                       (N104)? mem[870] : 
                       (N106)? mem[932] : 
                       (N108)? mem[994] : 
                       (N110)? mem[1056] : 
                       (N112)? mem[1118] : 
                       (N114)? mem[1180] : 
                       (N116)? mem[1242] : 
                       (N118)? mem[1304] : 
                       (N120)? mem[1366] : 
                       (N122)? mem[1428] : 
                       (N124)? mem[1490] : 
                       (N126)? mem[1552] : 
                       (N128)? mem[1614] : 
                       (N130)? mem[1676] : 
                       (N132)? mem[1738] : 
                       (N134)? mem[1800] : 
                       (N136)? mem[1862] : 
                       (N138)? mem[1924] : 
                       (N77)? mem[1986] : 
                       (N79)? mem[2048] : 
                       (N81)? mem[2110] : 
                       (N83)? mem[2172] : 
                       (N85)? mem[2234] : 
                       (N87)? mem[2296] : 
                       (N89)? mem[2358] : 
                       (N91)? mem[2420] : 
                       (N93)? mem[2482] : 
                       (N95)? mem[2544] : 
                       (N97)? mem[2606] : 
                       (N99)? mem[2668] : 
                       (N101)? mem[2730] : 
                       (N103)? mem[2792] : 
                       (N105)? mem[2854] : 
                       (N107)? mem[2916] : 
                       (N109)? mem[2978] : 
                       (N111)? mem[3040] : 
                       (N113)? mem[3102] : 
                       (N115)? mem[3164] : 
                       (N117)? mem[3226] : 
                       (N119)? mem[3288] : 
                       (N121)? mem[3350] : 
                       (N123)? mem[3412] : 
                       (N125)? mem[3474] : 
                       (N127)? mem[3536] : 
                       (N129)? mem[3598] : 
                       (N131)? mem[3660] : 
                       (N133)? mem[3722] : 
                       (N135)? mem[3784] : 
                       (N137)? mem[3846] : 
                       (N139)? mem[3908] : 1'b0;
  assign r_data_o[1] = (N76)? mem[1] : 
                       (N78)? mem[63] : 
                       (N80)? mem[125] : 
                       (N82)? mem[187] : 
                       (N84)? mem[249] : 
                       (N86)? mem[311] : 
                       (N88)? mem[373] : 
                       (N90)? mem[435] : 
                       (N92)? mem[497] : 
                       (N94)? mem[559] : 
                       (N96)? mem[621] : 
                       (N98)? mem[683] : 
                       (N100)? mem[745] : 
                       (N102)? mem[807] : 
                       (N104)? mem[869] : 
                       (N106)? mem[931] : 
                       (N108)? mem[993] : 
                       (N110)? mem[1055] : 
                       (N112)? mem[1117] : 
                       (N114)? mem[1179] : 
                       (N116)? mem[1241] : 
                       (N118)? mem[1303] : 
                       (N120)? mem[1365] : 
                       (N122)? mem[1427] : 
                       (N124)? mem[1489] : 
                       (N126)? mem[1551] : 
                       (N128)? mem[1613] : 
                       (N130)? mem[1675] : 
                       (N132)? mem[1737] : 
                       (N134)? mem[1799] : 
                       (N136)? mem[1861] : 
                       (N138)? mem[1923] : 
                       (N77)? mem[1985] : 
                       (N79)? mem[2047] : 
                       (N81)? mem[2109] : 
                       (N83)? mem[2171] : 
                       (N85)? mem[2233] : 
                       (N87)? mem[2295] : 
                       (N89)? mem[2357] : 
                       (N91)? mem[2419] : 
                       (N93)? mem[2481] : 
                       (N95)? mem[2543] : 
                       (N97)? mem[2605] : 
                       (N99)? mem[2667] : 
                       (N101)? mem[2729] : 
                       (N103)? mem[2791] : 
                       (N105)? mem[2853] : 
                       (N107)? mem[2915] : 
                       (N109)? mem[2977] : 
                       (N111)? mem[3039] : 
                       (N113)? mem[3101] : 
                       (N115)? mem[3163] : 
                       (N117)? mem[3225] : 
                       (N119)? mem[3287] : 
                       (N121)? mem[3349] : 
                       (N123)? mem[3411] : 
                       (N125)? mem[3473] : 
                       (N127)? mem[3535] : 
                       (N129)? mem[3597] : 
                       (N131)? mem[3659] : 
                       (N133)? mem[3721] : 
                       (N135)? mem[3783] : 
                       (N137)? mem[3845] : 
                       (N139)? mem[3907] : 1'b0;
  assign r_data_o[0] = (N76)? mem[0] : 
                       (N78)? mem[62] : 
                       (N80)? mem[124] : 
                       (N82)? mem[186] : 
                       (N84)? mem[248] : 
                       (N86)? mem[310] : 
                       (N88)? mem[372] : 
                       (N90)? mem[434] : 
                       (N92)? mem[496] : 
                       (N94)? mem[558] : 
                       (N96)? mem[620] : 
                       (N98)? mem[682] : 
                       (N100)? mem[744] : 
                       (N102)? mem[806] : 
                       (N104)? mem[868] : 
                       (N106)? mem[930] : 
                       (N108)? mem[992] : 
                       (N110)? mem[1054] : 
                       (N112)? mem[1116] : 
                       (N114)? mem[1178] : 
                       (N116)? mem[1240] : 
                       (N118)? mem[1302] : 
                       (N120)? mem[1364] : 
                       (N122)? mem[1426] : 
                       (N124)? mem[1488] : 
                       (N126)? mem[1550] : 
                       (N128)? mem[1612] : 
                       (N130)? mem[1674] : 
                       (N132)? mem[1736] : 
                       (N134)? mem[1798] : 
                       (N136)? mem[1860] : 
                       (N138)? mem[1922] : 
                       (N77)? mem[1984] : 
                       (N79)? mem[2046] : 
                       (N81)? mem[2108] : 
                       (N83)? mem[2170] : 
                       (N85)? mem[2232] : 
                       (N87)? mem[2294] : 
                       (N89)? mem[2356] : 
                       (N91)? mem[2418] : 
                       (N93)? mem[2480] : 
                       (N95)? mem[2542] : 
                       (N97)? mem[2604] : 
                       (N99)? mem[2666] : 
                       (N101)? mem[2728] : 
                       (N103)? mem[2790] : 
                       (N105)? mem[2852] : 
                       (N107)? mem[2914] : 
                       (N109)? mem[2976] : 
                       (N111)? mem[3038] : 
                       (N113)? mem[3100] : 
                       (N115)? mem[3162] : 
                       (N117)? mem[3224] : 
                       (N119)? mem[3286] : 
                       (N121)? mem[3348] : 
                       (N123)? mem[3410] : 
                       (N125)? mem[3472] : 
                       (N127)? mem[3534] : 
                       (N129)? mem[3596] : 
                       (N131)? mem[3658] : 
                       (N133)? mem[3720] : 
                       (N135)? mem[3782] : 
                       (N137)? mem[3844] : 
                       (N139)? mem[3906] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3967_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3966_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3965_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3964_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3963_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3962_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3961_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3960_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3959_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3958_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3957_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3956_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3955_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3954_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3953_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3952_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3951_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3950_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3949_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3948_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3947_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3946_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3945_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3944_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3943_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3942_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3941_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3940_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3939_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3938_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3937_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3936_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3935_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3934_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3933_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3932_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3931_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3930_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3929_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3928_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3927_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3926_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3925_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3924_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3923_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3922_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3921_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3920_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3919_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3918_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3917_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3916_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3915_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3914_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3913_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3912_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3911_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3910_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3909_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3908_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3907_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N268) begin
      mem_3906_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3905_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3904_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3903_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3902_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3901_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3900_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3899_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3898_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3897_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3896_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3895_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3894_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3893_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3892_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3891_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3890_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3889_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3888_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3887_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3886_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3885_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3884_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3883_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3882_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3881_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3880_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3879_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3878_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3877_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3876_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3875_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3874_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3873_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3872_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3871_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3870_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3869_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3868_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3867_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3866_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3865_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3864_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3863_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3862_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3861_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3860_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3859_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3858_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3857_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3856_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3855_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3854_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3853_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3852_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3851_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3850_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3849_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3848_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3847_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3846_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3845_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N267) begin
      mem_3844_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3843_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3842_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3841_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3840_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3839_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3838_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3837_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3836_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3835_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3834_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3833_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3832_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3831_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3830_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3829_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3828_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3827_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3826_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3825_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3824_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3823_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3822_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3821_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3820_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3819_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3818_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3817_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3816_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3815_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3814_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3813_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3812_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3811_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3810_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3809_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3808_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3807_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3806_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3805_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3804_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3803_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3802_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3801_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3800_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3799_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3798_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3797_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3796_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3795_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3794_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3793_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3792_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3791_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3790_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3789_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3788_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3787_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3786_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3785_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3784_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3783_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N266) begin
      mem_3782_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3781_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3780_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3779_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3778_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3777_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3776_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3775_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3774_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3773_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3772_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3771_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3770_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3769_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3768_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3767_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3766_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3765_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3764_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3763_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3762_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3761_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3760_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3759_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3758_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3757_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3756_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3755_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3754_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3753_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3752_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3751_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3750_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3749_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3748_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3747_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3746_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3745_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3744_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3743_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3742_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3741_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3740_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3739_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3738_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3737_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3736_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3735_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3734_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3733_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3732_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3731_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3730_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3729_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3728_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3727_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3726_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3725_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3724_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3723_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3722_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3721_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N265) begin
      mem_3720_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3719_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3718_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3717_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3716_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3715_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3714_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3713_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3712_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3711_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3710_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3709_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3708_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3707_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3706_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3705_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3704_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3703_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3702_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3701_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3700_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3699_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3698_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3697_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3696_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3695_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3694_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3693_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3692_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3691_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3690_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3689_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3688_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3687_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3686_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3685_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3684_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3683_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3682_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3681_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3680_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3679_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3678_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3677_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3676_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3675_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3674_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3673_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3672_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3671_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3670_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3669_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3668_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3667_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3666_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3665_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3664_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3663_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3662_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3661_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3660_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3659_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N264) begin
      mem_3658_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3657_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3656_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3655_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3654_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3653_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3652_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3651_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3650_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3649_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3648_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3647_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3646_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3645_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3644_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3643_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3642_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3641_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3640_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3639_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3638_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3637_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3636_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3635_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3634_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3633_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3632_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3631_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3630_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3629_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3628_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3627_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3626_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3625_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3624_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3623_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3622_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3621_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3620_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3619_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3618_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3617_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3616_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3615_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3614_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3613_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3612_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3611_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3610_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3609_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3608_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3607_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3606_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3605_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3604_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3603_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3602_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3601_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3600_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3599_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3598_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3597_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N263) begin
      mem_3596_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3595_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3594_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3593_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3592_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3591_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3590_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3589_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3588_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3587_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3586_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3585_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3584_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3583_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3582_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3581_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3580_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3579_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3578_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3577_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3576_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3575_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3574_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3573_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3572_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3571_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3570_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3569_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3568_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3567_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3566_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3565_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3564_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3563_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3562_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3561_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3560_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3559_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3558_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3557_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3556_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3555_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3554_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3553_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3552_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3551_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3550_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3549_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3548_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3547_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3546_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3545_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3544_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3543_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3542_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3541_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3540_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3539_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3538_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3537_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3536_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3535_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N262) begin
      mem_3534_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3533_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3532_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3531_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3530_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3529_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3528_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3527_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3526_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3525_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3524_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3523_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3522_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3521_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3520_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3519_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3518_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3517_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3516_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3515_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3514_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3513_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3512_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3511_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3510_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3509_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3508_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3507_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3506_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3505_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3504_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3503_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3502_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3501_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3500_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3499_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3498_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3497_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3496_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3495_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3494_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3493_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3492_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3491_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3490_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3489_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3488_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3487_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3486_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3485_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3484_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3483_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3482_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3481_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3480_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3479_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3478_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3477_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3476_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3475_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3474_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3473_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N261) begin
      mem_3472_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3471_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3470_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3469_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3468_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3467_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3466_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3465_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3464_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3463_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3462_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3461_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3460_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3459_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3458_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3457_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3456_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3455_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3454_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3453_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3452_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3451_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3450_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3449_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3448_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3447_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3446_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3445_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3444_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3443_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3442_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3441_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3440_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3439_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3438_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3437_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3436_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3435_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3434_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3433_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3432_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3431_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3430_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3429_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3428_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3427_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3426_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3425_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3424_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3423_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3422_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3421_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3420_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3419_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3418_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3417_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3416_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3415_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3414_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3413_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3412_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3411_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N260) begin
      mem_3410_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3409_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3408_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3407_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3406_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3405_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3404_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3403_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3402_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3401_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3400_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3399_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3398_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3397_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3396_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3395_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3394_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3393_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3392_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3391_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3390_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3389_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3388_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3387_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3386_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3385_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3384_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3383_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3382_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3381_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3380_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3379_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3378_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3377_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3376_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3375_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3374_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3373_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3372_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3371_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3370_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3369_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3368_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3367_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3366_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3365_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3364_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3363_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3362_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3361_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3360_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3359_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3358_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3357_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3356_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3355_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3354_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3353_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3352_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3351_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3350_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3349_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N259) begin
      mem_3348_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3347_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3346_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3345_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3344_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3343_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3342_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3341_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3340_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3339_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3338_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3337_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3336_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3335_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3334_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3333_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3332_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3331_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3330_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3329_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3328_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3327_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3326_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3325_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3324_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3323_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3322_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3321_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3320_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3319_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3318_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3317_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3316_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3315_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3314_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3313_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3312_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3311_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3310_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3309_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3308_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3307_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3306_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3305_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3304_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3303_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3302_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3301_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3300_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3299_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3298_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3297_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3296_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3295_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3294_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3293_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3292_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3291_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3290_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3289_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3288_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3287_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N258) begin
      mem_3286_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3285_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3284_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3283_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3282_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3281_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3280_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3279_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3278_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3277_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3276_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3275_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3274_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3273_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3272_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3271_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3270_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3269_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3268_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3267_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3266_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3265_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3264_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3263_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3262_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3261_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3260_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3259_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3258_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3257_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3256_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3255_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3254_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3253_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3252_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3251_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3250_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3249_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3248_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3247_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3246_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3245_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3244_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3243_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3242_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3241_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3240_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3239_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3238_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3237_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3236_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3235_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3234_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3233_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3232_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3231_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3230_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3229_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3228_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3227_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3226_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3225_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N257) begin
      mem_3224_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3223_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3222_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3221_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3220_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3219_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3218_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3217_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3216_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3215_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3214_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3213_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3212_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3211_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3210_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3209_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3208_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3207_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3206_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3205_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3204_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3203_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3202_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3201_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3200_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3199_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3198_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3197_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3196_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3195_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3194_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3193_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3192_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3191_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3190_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3189_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3188_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3187_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3186_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3185_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3184_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3183_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3182_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3181_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3180_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3179_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3178_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3177_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3176_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3175_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3174_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3173_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3172_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3171_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3170_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3169_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3168_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3167_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3166_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3165_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3164_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3163_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N256) begin
      mem_3162_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3161_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3160_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3159_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3158_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3157_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3156_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3155_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3154_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3153_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3152_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3151_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3150_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3149_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3148_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3147_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3146_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3145_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3144_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3143_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3142_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3141_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3140_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3139_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3138_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3137_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3136_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3135_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3134_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3133_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3132_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3131_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3130_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3129_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3128_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3127_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3126_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3125_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3124_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3123_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3122_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3121_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3120_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3119_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3118_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3117_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3116_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3115_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3114_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3113_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3112_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3111_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3110_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3109_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3108_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3107_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3106_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3105_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3104_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3103_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3102_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3101_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N255) begin
      mem_3100_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3099_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3098_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3097_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3096_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3095_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3094_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3093_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3092_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3091_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3090_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3089_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3088_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3087_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3086_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3085_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3084_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3083_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3082_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3081_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3080_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3079_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3078_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3077_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3076_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3075_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3074_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3073_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3072_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3071_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3070_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3069_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3068_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3067_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3066_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3065_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3064_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3063_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3062_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3061_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3060_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3059_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3058_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3057_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3056_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3055_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3054_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3053_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3052_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3051_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3050_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3049_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3048_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3047_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3046_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3045_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3044_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3043_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3042_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3041_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3040_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3039_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N254) begin
      mem_3038_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3037_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3036_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3035_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3034_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3033_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3032_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3031_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3030_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3029_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3028_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3027_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3026_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3025_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3024_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3023_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3022_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3021_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3020_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3019_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3018_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3017_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3016_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3015_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3014_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3013_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3012_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3011_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3010_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3009_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3008_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3007_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3006_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3005_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3004_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3003_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3002_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3001_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_3000_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2999_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2998_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2997_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2996_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2995_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2994_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2993_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2992_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2991_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2990_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2989_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2988_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2987_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2986_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2985_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2984_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2983_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2982_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2981_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2980_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2979_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2978_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2977_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N253) begin
      mem_2976_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2975_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2974_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2973_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2972_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2971_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2970_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2969_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2968_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2967_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2966_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2965_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2964_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2963_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2962_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2961_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2960_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2959_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2958_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2957_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2956_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2955_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2954_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2953_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2952_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2951_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2950_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2949_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2948_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2947_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2946_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2945_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2944_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2943_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2942_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2941_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2940_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2939_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2938_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2937_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2936_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2935_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2934_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2933_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2932_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2931_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2930_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2929_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2928_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2927_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2926_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2925_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2924_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2923_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2922_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2921_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2920_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2919_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2918_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2917_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2916_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2915_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N252) begin
      mem_2914_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2913_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2912_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2911_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2910_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2909_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2908_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2907_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2906_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2905_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2904_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2903_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2902_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2901_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2900_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2899_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2898_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2897_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2896_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2895_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2894_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2893_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2892_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2891_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2890_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2889_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2888_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2887_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2886_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2885_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2884_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2883_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2882_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2881_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2880_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2879_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2878_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2877_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2876_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2875_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2874_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2873_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2872_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2871_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2870_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2869_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2868_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2867_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2866_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2865_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2864_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2863_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2862_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2861_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2860_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2859_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2858_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2857_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2856_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2855_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2854_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2853_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N251) begin
      mem_2852_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2851_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2850_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2849_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2848_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2847_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2846_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2845_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2844_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2843_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2842_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2841_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2840_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2839_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2838_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2837_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2836_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2835_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2834_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2833_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2832_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2831_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2830_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2829_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2828_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2827_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2826_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2825_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2824_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2823_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2822_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2821_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2820_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2819_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2818_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2817_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2816_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2815_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2814_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2813_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2812_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2811_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2810_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2809_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2808_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2807_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2806_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2805_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2804_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2803_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2802_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2801_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2800_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2799_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2798_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2797_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2796_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2795_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2794_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2793_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2792_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2791_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N250) begin
      mem_2790_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2789_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2788_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2787_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2786_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2785_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2784_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2783_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2782_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2781_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2780_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2779_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2778_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2777_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2776_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2775_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2774_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2773_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2772_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2771_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2770_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2769_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2768_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2767_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2766_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2765_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2764_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2763_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2762_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2761_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2760_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2759_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2758_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2757_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2756_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2755_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2754_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2753_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2752_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2751_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2750_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2749_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2748_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2747_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2746_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2745_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2744_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2743_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2742_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2741_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2740_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2739_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2738_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2737_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2736_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2735_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2734_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2733_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2732_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2731_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2730_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2729_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N249) begin
      mem_2728_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2727_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2726_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2725_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2724_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2723_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2722_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2721_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2720_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2719_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2718_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2717_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2716_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2715_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2714_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2713_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2712_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2711_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2710_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2709_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2708_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2707_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2706_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2705_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2704_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2703_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2702_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2701_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2700_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2699_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2698_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2697_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2696_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2695_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2694_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2693_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2692_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2691_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2690_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2689_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2688_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2687_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2686_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2685_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2684_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2683_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2682_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2681_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2680_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2679_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2678_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2677_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2676_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2675_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2674_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2673_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2672_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2671_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2670_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2669_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2668_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2667_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N248) begin
      mem_2666_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2665_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2664_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2663_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2662_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2661_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2660_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2659_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2658_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2657_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2656_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2655_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2654_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2653_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2652_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2651_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2650_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2649_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2648_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2647_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2646_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2645_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2644_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2643_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2642_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2641_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2640_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2639_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2638_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2637_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2636_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2635_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2634_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2633_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2632_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2631_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2630_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2629_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2628_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2627_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2626_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2625_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2624_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2623_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2622_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2621_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2620_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2619_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2618_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2617_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2616_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2615_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2614_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2613_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2612_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2611_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2610_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2609_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2608_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2607_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2606_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2605_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N247) begin
      mem_2604_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2603_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2602_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2601_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2600_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2599_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2598_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2597_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2596_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2595_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2594_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2593_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2592_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2591_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2590_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2589_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2588_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2587_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2586_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2585_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2584_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2583_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2582_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2581_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2580_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2579_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2578_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2577_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2576_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2575_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2574_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2573_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2572_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2571_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2570_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2569_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2568_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2567_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2566_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2565_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2564_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2563_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2562_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2561_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2560_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2559_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2558_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2557_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2556_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2555_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2554_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2553_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2552_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2551_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2550_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2549_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2548_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2547_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2546_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2545_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2544_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2543_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N246) begin
      mem_2542_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2541_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2540_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2539_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2538_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2537_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2536_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2535_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2534_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2533_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2532_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2531_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2530_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2529_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2528_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2527_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2526_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2525_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2524_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2523_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2522_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2521_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2520_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2519_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2518_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2517_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2516_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2515_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2514_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2513_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2512_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2511_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2510_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2509_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2508_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2507_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2506_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2505_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2504_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2503_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2502_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2501_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2500_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2499_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2498_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2497_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2496_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2495_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2494_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2493_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2492_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2491_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2490_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2489_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2488_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2487_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2486_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2485_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2484_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2483_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2482_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2481_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N245) begin
      mem_2480_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2479_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2478_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2477_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2476_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2475_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2474_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2473_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2472_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2471_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2470_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2469_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2468_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2467_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2466_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2465_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2464_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2463_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2462_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2461_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2460_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2459_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2458_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2457_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2456_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2455_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2454_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2453_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2452_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2451_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2450_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2449_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2448_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2447_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2446_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2445_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2444_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2443_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2442_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2441_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2440_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2439_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2438_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2437_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2436_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2435_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2434_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2433_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2432_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2431_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2430_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2429_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2428_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2427_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2426_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2425_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2424_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2423_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2422_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2421_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2420_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2419_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N244) begin
      mem_2418_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2417_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2416_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2415_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2414_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2413_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2412_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2411_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2410_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2409_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2408_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2407_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2406_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2405_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2404_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2403_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2402_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2401_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2400_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2399_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2398_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2397_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2396_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2395_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2394_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2393_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2392_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2391_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2390_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2389_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2388_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2387_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2386_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2385_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2384_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2383_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2382_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2381_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2380_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2379_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2378_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2377_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2376_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2375_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2374_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2373_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2372_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2371_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2370_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2369_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2368_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2367_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2366_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2365_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2364_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2363_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2362_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2361_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2360_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2359_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2358_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2357_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N243) begin
      mem_2356_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2355_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2354_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2353_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2352_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2351_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2350_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2349_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2348_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2347_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2346_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2345_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2344_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2343_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2342_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2341_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2340_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2339_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2338_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2337_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2336_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2335_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2334_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2333_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2332_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2331_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2330_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2329_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2328_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2327_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2326_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2325_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2324_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2323_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2322_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2321_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2320_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2319_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2318_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2317_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2316_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2315_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2314_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2313_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2312_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2311_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2310_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2309_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2308_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2307_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2306_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2305_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2304_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2303_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2302_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2301_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2300_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2299_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2298_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2297_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2296_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2295_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N242) begin
      mem_2294_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2293_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2292_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2291_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2290_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2289_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2288_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2287_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2286_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2285_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2284_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2283_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2282_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2281_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2280_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2279_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2278_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2277_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2276_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2275_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2274_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2273_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2272_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2271_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2270_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2269_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2268_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2267_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2266_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2265_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2264_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2263_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2262_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2261_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2260_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2259_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2258_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2257_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2256_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2255_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2254_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2253_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2252_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2251_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2250_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2249_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2248_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2247_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2246_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2245_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2244_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2243_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2242_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2241_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2240_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2239_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2238_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2237_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2236_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2235_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2234_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2233_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N241) begin
      mem_2232_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2231_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2230_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2229_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2228_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2227_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2226_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2225_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2224_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2223_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2222_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2221_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2220_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2219_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2218_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2217_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2216_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2215_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2214_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2213_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2212_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2211_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2210_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2209_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2208_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2207_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2206_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2205_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2204_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2203_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2202_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2201_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2200_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2199_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2198_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2197_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2196_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2195_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2194_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2193_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2192_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2191_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2190_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2189_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2188_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2187_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2186_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2185_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2184_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2183_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2182_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2181_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2180_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2179_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2178_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2177_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2176_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2175_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2174_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2173_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2172_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2171_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N240) begin
      mem_2170_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2169_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2168_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2167_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2166_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2165_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2164_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2163_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2162_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2161_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2160_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2159_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2158_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2157_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2156_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2155_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2154_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2153_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2152_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2151_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2150_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2149_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2148_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2147_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2146_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2145_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2144_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2143_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2142_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2141_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2140_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2139_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2138_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2137_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2136_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2135_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2134_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2133_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2132_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2131_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2130_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2129_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2128_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2127_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2126_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2125_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2124_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2123_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2122_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2121_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2120_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2119_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2118_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2117_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2116_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2115_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2114_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2113_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2112_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2111_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2110_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2109_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N239) begin
      mem_2108_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2107_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2106_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2105_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2104_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2103_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2102_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2101_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2100_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2099_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2098_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2097_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2096_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2095_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2094_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2093_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2092_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2091_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2090_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2089_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2088_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2087_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2086_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2085_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2084_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2083_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2082_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2081_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2080_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2079_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2078_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2077_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2076_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2075_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2074_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2073_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2072_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2071_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2070_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2069_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2068_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2067_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2066_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2065_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2064_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2063_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2062_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2061_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2060_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2059_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2058_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2057_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2056_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2055_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2054_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2053_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2052_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2051_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2050_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2049_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2048_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2047_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N238) begin
      mem_2046_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2045_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2044_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2043_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2042_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2041_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2040_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2039_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2038_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2037_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2036_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2035_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2034_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2033_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2032_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2031_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2030_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2029_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2028_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2027_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2026_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2025_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2024_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2023_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2022_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2021_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2020_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2019_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2018_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2017_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2016_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2015_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2014_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2013_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2012_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2011_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2010_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2009_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2008_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2007_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2006_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2005_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2004_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2003_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2002_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2001_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_2000_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1999_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1998_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1997_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1996_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1995_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1994_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1993_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1992_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1991_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1990_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1989_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1988_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1987_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1986_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1985_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N237) begin
      mem_1984_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1983_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1982_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1981_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1980_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1979_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1978_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1977_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1976_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1975_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1974_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1973_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1972_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1971_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1970_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1969_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1968_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1967_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1966_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1965_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1964_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1963_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1962_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1961_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1960_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1959_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1958_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1957_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1956_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1955_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1954_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1953_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1952_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1951_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1950_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1949_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1948_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1947_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1946_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1945_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1944_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1943_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1942_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1941_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1940_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1939_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1938_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1937_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1936_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1935_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1934_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1933_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1932_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1931_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1930_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1929_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1928_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1927_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1926_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1925_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1924_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1923_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N236) begin
      mem_1922_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1921_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1920_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1919_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1918_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1917_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1916_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1915_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1914_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1913_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1912_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1911_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1910_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1909_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1908_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1907_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1906_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1905_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1904_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1903_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1902_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1901_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1900_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1899_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1898_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1897_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1896_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1895_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1894_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1893_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1892_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1891_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1890_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1889_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1888_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1887_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1886_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1885_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1884_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1883_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1882_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1881_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1880_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1879_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1878_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1877_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1876_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1875_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1874_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1873_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1872_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1871_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1870_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1869_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1868_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1867_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1866_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1865_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1864_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1863_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1862_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1861_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N235) begin
      mem_1860_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1859_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1858_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1857_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1856_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1855_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1854_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1853_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1852_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1851_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1850_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1849_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1848_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1847_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1846_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1845_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1844_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1843_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1842_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1841_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1840_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1839_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1838_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1837_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1836_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1835_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1834_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1833_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1832_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1831_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1830_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1829_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1828_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1827_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1826_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1825_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1824_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1823_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1822_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1821_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1820_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1819_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1818_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1817_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1816_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1815_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1814_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1813_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1812_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1811_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1810_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1809_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1808_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1807_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1806_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1805_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1804_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1803_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1802_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1801_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1800_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1799_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N234) begin
      mem_1798_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1797_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1796_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1795_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1794_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1793_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1792_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1791_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1790_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1789_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1788_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1787_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1786_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1785_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1784_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1783_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1782_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1781_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1780_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1779_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1778_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1777_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1776_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1775_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1774_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1773_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1772_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1771_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1770_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1769_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1768_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1767_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1766_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1765_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1764_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1763_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1762_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1761_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1760_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1759_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1758_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1757_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1756_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1755_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1754_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1753_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1752_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1751_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1750_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1749_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1748_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1747_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1746_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1745_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1744_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1743_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1742_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1741_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1740_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1739_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1738_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1737_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N233) begin
      mem_1736_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1735_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1734_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1733_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1732_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1731_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1730_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1729_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1728_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1727_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1726_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1725_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1724_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1723_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1722_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1721_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1720_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1719_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1718_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1717_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1716_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1715_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1714_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1713_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1712_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1711_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1710_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1709_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1708_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1707_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1706_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1705_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1704_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1703_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1702_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1701_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1700_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1699_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1698_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1697_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1696_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1695_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1694_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1693_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1692_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1691_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1690_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1689_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1688_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1687_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1686_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1685_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1684_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1683_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1682_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1681_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1680_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1679_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1678_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1677_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1676_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1675_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N232) begin
      mem_1674_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1673_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1672_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1671_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1670_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1669_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1668_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1667_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1666_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1665_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1664_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1663_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1662_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1661_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1660_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1659_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1658_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1657_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1656_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1655_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1654_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1653_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1652_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1651_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1650_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1649_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1648_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1647_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1646_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1645_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1644_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1643_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1642_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1641_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1640_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1639_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1638_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1637_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1636_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1635_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1634_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1633_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1632_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1631_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1630_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1629_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1628_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1627_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1626_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1625_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1624_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1623_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1622_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1621_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1620_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1619_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1618_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1617_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1616_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1615_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1614_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1613_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N231) begin
      mem_1612_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1611_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1610_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1609_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1608_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1607_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1606_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1605_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1604_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1603_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1602_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1601_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1600_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1599_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1598_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1597_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1596_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1595_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1594_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1593_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1592_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1591_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1590_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1589_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1588_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1587_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1586_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1585_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1584_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1583_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1582_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1581_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1580_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1579_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1578_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1577_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1576_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1575_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1574_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1573_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1572_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1571_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1570_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1569_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1568_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1567_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1566_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1565_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1564_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1563_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1562_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1561_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1560_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1559_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1558_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1557_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1556_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1555_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1554_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1553_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1552_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1551_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N230) begin
      mem_1550_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1549_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1548_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1547_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1546_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1545_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1544_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1543_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1542_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1541_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1540_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1539_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1538_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1537_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1536_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1535_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1534_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1533_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1532_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1531_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1530_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1529_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1528_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1527_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1526_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1525_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1524_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1523_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1522_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1521_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1520_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1519_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1518_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1517_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1516_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1515_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1514_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1513_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1512_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1511_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1510_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1509_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1508_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1507_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1506_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1505_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1504_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1503_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1502_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1501_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1500_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1499_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1498_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1497_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1496_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1495_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1494_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1493_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1492_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1491_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1490_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1489_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N229) begin
      mem_1488_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1487_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1486_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1485_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1484_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1483_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1482_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1481_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1480_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1479_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1478_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1477_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1476_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1475_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1474_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1473_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1472_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1471_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1470_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1469_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1468_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1467_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1466_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1465_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1464_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1463_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1462_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1461_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1460_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1459_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1458_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1457_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1456_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1455_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1454_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1453_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1452_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1451_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1450_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1449_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1448_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1447_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1446_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1445_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1444_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1443_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1442_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1441_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1440_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1439_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1438_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1437_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1436_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1435_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1434_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1433_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1432_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1431_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1430_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1429_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1428_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1427_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N228) begin
      mem_1426_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1425_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1424_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1423_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1422_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1421_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1420_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1419_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1418_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1417_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1416_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1415_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1414_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1413_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1412_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1411_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1410_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1409_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1408_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1407_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1406_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1405_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1404_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1403_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1402_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1401_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1400_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1399_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1398_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1397_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1396_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1395_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1394_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1393_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1392_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1391_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1390_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1389_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1388_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1387_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1386_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1385_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1384_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1383_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1382_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1381_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1380_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1379_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1378_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1377_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1376_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1375_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1374_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1373_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1372_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1371_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1370_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1369_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1368_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1367_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1366_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1365_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N227) begin
      mem_1364_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1363_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1362_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1361_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1360_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1359_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1358_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1357_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1356_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1355_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1354_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1353_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1352_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1351_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1350_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1349_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1348_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1347_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1346_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1345_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1344_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1343_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1342_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1341_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1340_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1339_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1338_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1337_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1336_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1335_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1334_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1333_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1332_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1331_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1330_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1329_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1328_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1327_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1326_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1325_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1324_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1323_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1322_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1321_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1320_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1319_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1318_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1317_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1316_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1315_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1314_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1313_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1312_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1311_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1310_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1309_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1308_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1307_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1306_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1305_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1304_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1303_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N226) begin
      mem_1302_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1301_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1300_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1299_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1298_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1297_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1296_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1295_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1294_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1293_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1292_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1291_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1290_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1289_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1288_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1287_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1286_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1285_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1284_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1283_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1282_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1281_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1280_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1279_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1278_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1277_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1276_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1275_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1274_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1273_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1272_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1271_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1270_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1269_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1268_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1267_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1266_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1265_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1264_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1263_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1262_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1261_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1260_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1259_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1258_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1257_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1256_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1255_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1254_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1253_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1252_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1251_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1250_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1249_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1248_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1247_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1246_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1245_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1244_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1243_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1242_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1241_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N225) begin
      mem_1240_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1239_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1238_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1237_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1236_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1235_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1234_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1233_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1232_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1231_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1230_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1229_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1228_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1227_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1226_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1225_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1224_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1223_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1222_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1221_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1220_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1219_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1218_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1217_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1216_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1215_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1214_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1213_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1212_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1211_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1210_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1209_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1208_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1207_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1206_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1205_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1204_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1203_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1202_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1201_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1200_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1199_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1198_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1197_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1196_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1195_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1194_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1193_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1192_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1191_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1190_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1189_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1188_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1187_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1186_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1185_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1184_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1183_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1182_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1181_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1180_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1179_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N224) begin
      mem_1178_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1177_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1176_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1175_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1174_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1173_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1172_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1171_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1170_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1169_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1168_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1167_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1166_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1165_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1164_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1163_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1162_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1161_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1160_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1159_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1158_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1157_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1156_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1155_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1154_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1153_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1152_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1151_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1150_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1149_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1148_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1147_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1146_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1145_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1144_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1143_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1142_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1141_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1140_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1139_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1138_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1137_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1136_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1135_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1134_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1133_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1132_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1131_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1130_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1129_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1128_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1127_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1126_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1125_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1124_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1123_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1122_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1121_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1120_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1119_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1118_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1117_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N223) begin
      mem_1116_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1115_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1114_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1113_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1112_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1111_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1110_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1109_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1108_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1107_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1106_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1105_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1104_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1103_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1102_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1101_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1100_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1099_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1098_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1097_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1096_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1095_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1094_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1093_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1092_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1091_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1090_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1089_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1088_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1087_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1086_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1085_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1084_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1083_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1082_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1081_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1080_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1079_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1078_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1077_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1076_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1075_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1074_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1073_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1072_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1071_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1070_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1069_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1068_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1067_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1066_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1065_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1064_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1063_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1062_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1061_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1060_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1059_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1058_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1057_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1056_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1055_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N222) begin
      mem_1054_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1053_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1052_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1051_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1050_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1049_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1048_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1047_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1046_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1045_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1044_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1043_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1042_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1041_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1040_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1039_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1038_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1037_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1036_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1035_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1034_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1033_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1032_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1031_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1030_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1029_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1028_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1027_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1026_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1025_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1024_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1023_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1022_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1021_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1020_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1019_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1018_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1017_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1016_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1015_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1014_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1013_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1012_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1011_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1010_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1009_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1008_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1007_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1006_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1005_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1004_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1003_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1002_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1001_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_1000_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_999_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_998_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_997_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_996_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_995_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_994_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_993_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N221) begin
      mem_992_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_991_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_990_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_989_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_988_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_987_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_986_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_985_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_984_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_983_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_982_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_981_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_980_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_979_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_978_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_977_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_976_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_975_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_974_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_973_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_972_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_971_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_970_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_969_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_968_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_967_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_966_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_965_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_964_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_963_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_962_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_961_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_960_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_959_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_958_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_957_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_956_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_955_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_954_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_953_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_952_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_951_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_950_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_949_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_948_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_947_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_946_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_945_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_944_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_943_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_942_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_941_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_940_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_939_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_938_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_937_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_936_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_935_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_934_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_933_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_932_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_931_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N220) begin
      mem_930_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_929_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_928_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_927_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_926_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_925_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_924_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_923_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_922_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_921_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_920_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_919_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_918_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_917_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_916_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_915_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_914_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_913_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_912_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_911_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_910_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_909_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_908_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_907_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_906_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_905_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_904_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_903_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_902_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_901_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_900_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_899_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_898_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_897_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_896_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_895_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_894_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_893_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_892_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_891_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_890_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_889_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_888_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_887_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_886_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_885_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_884_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_883_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_882_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_881_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_880_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_879_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_878_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_877_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_876_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_875_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_874_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_873_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_872_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_871_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_870_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_869_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N219) begin
      mem_868_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_867_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_866_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_865_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_864_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_863_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_862_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_861_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_860_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_859_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_858_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_857_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_856_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_855_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_854_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_853_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_852_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_851_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_850_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_849_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_848_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_847_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_846_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_845_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_844_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_843_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_842_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_841_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_840_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_839_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_838_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_837_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_836_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_835_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_834_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_833_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_832_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_831_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_830_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_829_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_828_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_827_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_826_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_825_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_824_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_823_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_822_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_821_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_820_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_819_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_818_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_817_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_816_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_815_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_814_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_813_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_812_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_811_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_810_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_809_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_808_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_807_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N218) begin
      mem_806_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_805_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_804_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_803_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_802_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_801_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_800_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_799_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_798_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_797_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_796_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_795_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_794_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_793_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_792_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_791_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_790_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_789_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_788_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_787_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_786_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_785_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_784_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_783_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_782_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_781_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_780_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_779_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_778_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_777_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_776_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_775_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_774_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_773_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_772_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_771_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_770_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_769_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_768_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_767_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_766_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_765_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_764_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_763_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_762_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_761_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_760_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_759_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_758_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_757_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_756_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_755_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_754_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_753_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_752_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_751_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_750_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_749_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_748_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_747_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_746_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_745_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N217) begin
      mem_744_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_743_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_742_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_741_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_740_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_739_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_738_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_737_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_736_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_735_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_734_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_733_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_732_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_731_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_730_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_729_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_728_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_727_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_726_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_725_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_724_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_723_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_722_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_721_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_720_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_719_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_718_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_717_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_716_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_715_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_714_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_713_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_712_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_711_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_710_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_709_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_708_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_707_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_706_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_705_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_704_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_703_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_702_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_701_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_700_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_699_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_698_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_697_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_696_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_695_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_694_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_693_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_692_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_691_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_690_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_689_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_688_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_687_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_686_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_685_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_684_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_683_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N216) begin
      mem_682_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_681_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_680_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_679_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_678_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_677_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_676_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_675_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_674_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_673_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_672_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_671_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_670_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_669_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_668_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_667_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_666_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_665_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_664_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_663_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_662_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_661_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_660_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_659_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_658_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_657_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_656_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_655_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_654_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_653_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_652_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_651_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_650_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_649_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_648_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_647_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_646_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_645_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_644_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_643_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_642_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_641_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_640_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_639_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_638_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_637_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_636_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_635_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_634_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_633_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_632_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_631_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_630_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_629_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_628_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_627_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_626_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_625_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_624_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_623_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_622_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_621_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N215) begin
      mem_620_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_619_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_618_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_617_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_616_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_615_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_614_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_613_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_612_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_611_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_610_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_609_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_608_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_607_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_606_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_605_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_604_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_603_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_602_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_601_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_600_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_599_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_598_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_597_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_596_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_595_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_594_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_593_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_592_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_591_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_590_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_589_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_588_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_587_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_586_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_585_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_584_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_583_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_582_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_581_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_580_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_579_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_578_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_577_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_576_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_575_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_574_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_573_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_572_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_571_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_570_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_569_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_568_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_567_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_566_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_565_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_564_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_563_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_562_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_561_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_560_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_559_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N214) begin
      mem_558_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_557_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_556_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_555_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_554_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_553_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_552_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_551_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_550_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_549_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_548_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_547_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_546_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_545_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_544_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_543_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_542_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_541_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_540_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_539_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_538_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_537_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_536_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_535_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_534_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_533_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_532_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_531_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_530_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_529_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_528_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_527_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_526_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_525_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_524_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_523_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_522_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_521_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_520_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_519_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_518_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_517_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_516_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_515_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_514_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_513_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_512_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_511_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_510_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_509_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_508_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_507_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_506_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_505_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_504_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_503_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_502_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_501_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_500_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_499_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_498_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_497_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N213) begin
      mem_496_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_495_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_494_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_493_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_492_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_491_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_490_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_489_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_488_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_487_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_486_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_485_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_484_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_483_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_482_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_481_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_480_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_479_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_478_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_477_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_476_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_475_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_474_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_473_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_472_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_471_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_470_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_469_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_468_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_467_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_466_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_465_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_464_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_463_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_462_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_461_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_460_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_459_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_458_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_457_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_456_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_455_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_454_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_453_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_452_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_451_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_450_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_449_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_448_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_447_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_446_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_445_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_444_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_443_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_442_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_441_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_440_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_439_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_438_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_437_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_436_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_435_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N212) begin
      mem_434_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_433_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_432_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_431_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_430_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_429_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_428_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_427_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_426_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_425_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_424_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_423_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_422_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_421_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_420_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_419_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_418_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_417_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_416_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_415_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_414_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_413_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_412_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_411_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_410_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_409_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_408_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_407_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_406_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_405_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_404_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_403_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_402_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_401_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_400_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_399_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_398_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_397_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_396_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_395_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_394_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_393_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_392_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_391_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_390_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_389_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_388_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_387_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_386_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_385_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_384_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_383_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_382_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_381_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_380_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_379_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_378_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_377_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_376_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_375_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_374_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_373_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N211) begin
      mem_372_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_371_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_370_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_369_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_368_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_367_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_366_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_365_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_364_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_363_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_362_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_361_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_360_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_359_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_358_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_357_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_356_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_355_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_354_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_353_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_352_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_351_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_350_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_349_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_348_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_347_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_346_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_345_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_344_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_343_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_342_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_341_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_340_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_339_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_338_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_337_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_336_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_335_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_334_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_333_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_332_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_331_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_330_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_329_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_328_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_327_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_326_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_325_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_324_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_323_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_322_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_321_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_320_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_319_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_318_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_317_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_316_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_315_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_314_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_313_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_312_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_311_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N210) begin
      mem_310_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_309_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_308_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_307_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_306_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_305_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_304_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_303_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_302_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_301_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_300_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_299_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_298_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_297_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_296_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_295_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_294_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_293_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_292_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_291_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_290_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_289_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_288_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_287_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_286_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_285_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_284_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_283_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_282_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_281_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_280_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_279_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_278_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_277_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_276_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_275_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_274_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_273_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_272_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_271_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_270_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_269_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_268_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_267_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_266_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_265_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_264_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_263_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_262_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_261_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_260_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_259_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_258_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_257_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_256_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_255_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_254_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_253_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_252_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_251_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_250_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_249_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N209) begin
      mem_248_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_247_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_246_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_245_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_244_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_243_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_242_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_241_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_240_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_239_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_238_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_237_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_236_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_235_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_234_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_233_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_232_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_231_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_230_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_229_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_228_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_227_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_226_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_225_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_224_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_223_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_222_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_221_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_220_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_219_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_218_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_217_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_216_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_215_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_214_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_213_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_212_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_211_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_210_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_209_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_208_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_207_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_206_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_205_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_204_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_203_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_202_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_201_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_200_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_199_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_198_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_197_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_196_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_195_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_194_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_193_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_192_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_191_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_190_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_189_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_188_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_187_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N208) begin
      mem_186_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_185_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_184_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_183_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_182_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_181_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_180_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_179_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_178_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_177_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_176_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_175_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_174_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_173_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_172_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_171_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_170_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_169_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_168_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_167_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_166_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_165_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_164_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_163_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_162_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_161_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_160_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_159_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_158_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_157_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_156_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_155_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_154_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_153_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_152_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_151_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_150_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_149_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_148_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_147_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_146_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_145_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_144_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_143_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_142_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_141_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_140_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_139_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_138_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_137_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_136_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_135_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_134_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_133_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_132_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_131_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_130_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_129_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_128_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_127_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_126_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_125_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N207) begin
      mem_124_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_123_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_122_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_121_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_120_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_119_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_118_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_117_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_116_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_115_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_114_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_113_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_112_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_111_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_110_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_109_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_108_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_107_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_106_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_105_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_104_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_103_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_102_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_101_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_100_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_99_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_98_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_97_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_96_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_95_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_94_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_93_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_92_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_91_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_90_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_89_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_88_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_87_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_86_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_85_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_84_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_83_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_82_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_81_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_80_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_79_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_78_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_77_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_76_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_75_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_74_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_73_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_72_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_71_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_70_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_69_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_68_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_67_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_66_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_65_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_64_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_63_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N206) begin
      mem_62_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_61_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_60_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_59_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_58_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_57_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_56_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_55_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_54_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_53_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_52_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_51_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_50_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_49_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_48_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_47_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_46_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_45_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_44_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_43_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_42_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_41_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_40_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_39_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_38_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_37_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_36_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_35_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_34_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_33_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_32_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_31_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_30_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_29_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_28_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_27_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_26_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_25_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_24_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_23_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_22_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_21_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_20_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_19_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_18_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_17_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_16_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_15_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_14_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_13_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_12_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_11_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_10_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_9_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_8_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_7_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_6_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_5_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_4_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_3_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_2_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_1_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N205) begin
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end

  assign N269 = ~w_addr_i[5];
  assign N270 = w_addr_i[3] & w_addr_i[4];
  assign N271 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N272 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N273 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N274 = w_addr_i[5] & N270;
  assign N275 = w_addr_i[5] & N271;
  assign N276 = w_addr_i[5] & N272;
  assign N277 = w_addr_i[5] & N273;
  assign N278 = N269 & N270;
  assign N279 = N269 & N271;
  assign N280 = N269 & N272;
  assign N281 = N269 & N273;
  assign N282 = ~w_addr_i[2];
  assign N283 = w_addr_i[0] & w_addr_i[1];
  assign N284 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N285 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N286 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N287 = w_addr_i[2] & N283;
  assign N288 = w_addr_i[2] & N284;
  assign N289 = w_addr_i[2] & N285;
  assign N290 = w_addr_i[2] & N286;
  assign N291 = N282 & N283;
  assign N292 = N282 & N284;
  assign N293 = N282 & N285;
  assign N294 = N282 & N286;
  assign N204 = N274 & N287;
  assign N203 = N274 & N288;
  assign N202 = N274 & N289;
  assign N201 = N274 & N290;
  assign N200 = N274 & N291;
  assign N199 = N274 & N292;
  assign N198 = N274 & N293;
  assign N197 = N274 & N294;
  assign N196 = N275 & N287;
  assign N195 = N275 & N288;
  assign N194 = N275 & N289;
  assign N193 = N275 & N290;
  assign N192 = N275 & N291;
  assign N191 = N275 & N292;
  assign N190 = N275 & N293;
  assign N189 = N275 & N294;
  assign N188 = N276 & N287;
  assign N187 = N276 & N288;
  assign N186 = N276 & N289;
  assign N185 = N276 & N290;
  assign N184 = N276 & N291;
  assign N183 = N276 & N292;
  assign N182 = N276 & N293;
  assign N181 = N276 & N294;
  assign N180 = N277 & N287;
  assign N179 = N277 & N288;
  assign N178 = N277 & N289;
  assign N177 = N277 & N290;
  assign N176 = N277 & N291;
  assign N175 = N277 & N292;
  assign N174 = N277 & N293;
  assign N173 = N277 & N294;
  assign N172 = N278 & N287;
  assign N171 = N278 & N288;
  assign N170 = N278 & N289;
  assign N169 = N278 & N290;
  assign N168 = N278 & N291;
  assign N167 = N278 & N292;
  assign N166 = N278 & N293;
  assign N165 = N278 & N294;
  assign N164 = N279 & N287;
  assign N163 = N279 & N288;
  assign N162 = N279 & N289;
  assign N161 = N279 & N290;
  assign N160 = N279 & N291;
  assign N159 = N279 & N292;
  assign N158 = N279 & N293;
  assign N157 = N279 & N294;
  assign N156 = N280 & N287;
  assign N155 = N280 & N288;
  assign N154 = N280 & N289;
  assign N153 = N280 & N290;
  assign N152 = N280 & N291;
  assign N151 = N280 & N292;
  assign N150 = N280 & N293;
  assign N149 = N280 & N294;
  assign N148 = N281 & N287;
  assign N147 = N281 & N288;
  assign N146 = N281 & N289;
  assign N145 = N281 & N290;
  assign N144 = N281 & N291;
  assign N143 = N281 & N292;
  assign N142 = N281 & N293;
  assign N141 = N281 & N294;
  assign { N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205 } = (N8)? { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~r_addr_i[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_i[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_i[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_i[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_i[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = ~r_addr_i[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r_addr_i[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r_addr_i[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r_addr_i[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r_addr_i[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r_addr_i[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r_addr_i[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r_addr_i[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r_addr_i[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r_addr_i[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r_addr_i[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r_addr_i[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r_addr_i[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r_addr_i[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r_addr_i[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r_addr_i[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r_addr_i[4];
  assign N75 = ~r_addr_i[5];
  assign N76 = N43 & N75;
  assign N77 = N43 & r_addr_i[5];
  assign N78 = N45 & N75;
  assign N79 = N45 & r_addr_i[5];
  assign N80 = N47 & N75;
  assign N81 = N47 & r_addr_i[5];
  assign N82 = N49 & N75;
  assign N83 = N49 & r_addr_i[5];
  assign N84 = N51 & N75;
  assign N85 = N51 & r_addr_i[5];
  assign N86 = N53 & N75;
  assign N87 = N53 & r_addr_i[5];
  assign N88 = N55 & N75;
  assign N89 = N55 & r_addr_i[5];
  assign N90 = N57 & N75;
  assign N91 = N57 & r_addr_i[5];
  assign N92 = N59 & N75;
  assign N93 = N59 & r_addr_i[5];
  assign N94 = N61 & N75;
  assign N95 = N61 & r_addr_i[5];
  assign N96 = N63 & N75;
  assign N97 = N63 & r_addr_i[5];
  assign N98 = N65 & N75;
  assign N99 = N65 & r_addr_i[5];
  assign N100 = N67 & N75;
  assign N101 = N67 & r_addr_i[5];
  assign N102 = N69 & N75;
  assign N103 = N69 & r_addr_i[5];
  assign N104 = N71 & N75;
  assign N105 = N71 & r_addr_i[5];
  assign N106 = N73 & N75;
  assign N107 = N73 & r_addr_i[5];
  assign N108 = N44 & N75;
  assign N109 = N44 & r_addr_i[5];
  assign N110 = N46 & N75;
  assign N111 = N46 & r_addr_i[5];
  assign N112 = N48 & N75;
  assign N113 = N48 & r_addr_i[5];
  assign N114 = N50 & N75;
  assign N115 = N50 & r_addr_i[5];
  assign N116 = N52 & N75;
  assign N117 = N52 & r_addr_i[5];
  assign N118 = N54 & N75;
  assign N119 = N54 & r_addr_i[5];
  assign N120 = N56 & N75;
  assign N121 = N56 & r_addr_i[5];
  assign N122 = N58 & N75;
  assign N123 = N58 & r_addr_i[5];
  assign N124 = N60 & N75;
  assign N125 = N60 & r_addr_i[5];
  assign N126 = N62 & N75;
  assign N127 = N62 & r_addr_i[5];
  assign N128 = N64 & N75;
  assign N129 = N64 & r_addr_i[5];
  assign N130 = N66 & N75;
  assign N131 = N66 & r_addr_i[5];
  assign N132 = N68 & N75;
  assign N133 = N68 & r_addr_i[5];
  assign N134 = N70 & N75;
  assign N135 = N70 & r_addr_i[5];
  assign N136 = N72 & N75;
  assign N137 = N72 & r_addr_i[5];
  assign N138 = N74 & N75;
  assign N139 = N74 & r_addr_i[5];
  assign N140 = ~w_v_i;

endmodule