module RecFNToRecFN
(
  io_in,
  io_roundingMode,
  io_out,
  io_exceptionFlags
);

  input [32:0] io_in;
  input [1:0] io_roundingMode;
  output [64:0] io_out;
  output [4:0] io_exceptionFlags;
  wire [64:0] io_out;
  wire [4:0] io_exceptionFlags;
  wire N0,N1,outRawFloat_isNaN,T1,N2,outRawFloat_isInf,T24,T29,T42,N3,N4,N5,N6;
  wire [11:0] T20,T26,T33,T27,T36,T34;
  wire [11:11] T19,T21,T35,T46;
  wire [9:9] T28;
  assign io_out[28] = 1'b0;
  assign io_out[27] = 1'b0;
  assign io_out[26] = 1'b0;
  assign io_out[25] = 1'b0;
  assign io_out[24] = 1'b0;
  assign io_out[23] = 1'b0;
  assign io_out[22] = 1'b0;
  assign io_out[21] = 1'b0;
  assign io_out[20] = 1'b0;
  assign io_out[19] = 1'b0;
  assign io_out[18] = 1'b0;
  assign io_out[17] = 1'b0;
  assign io_out[16] = 1'b0;
  assign io_out[15] = 1'b0;
  assign io_out[14] = 1'b0;
  assign io_out[13] = 1'b0;
  assign io_out[12] = 1'b0;
  assign io_out[11] = 1'b0;
  assign io_out[10] = 1'b0;
  assign io_out[9] = 1'b0;
  assign io_out[8] = 1'b0;
  assign io_out[7] = 1'b0;
  assign io_out[6] = 1'b0;
  assign io_out[5] = 1'b0;
  assign io_out[4] = 1'b0;
  assign io_out[3] = 1'b0;
  assign io_out[2] = 1'b0;
  assign io_out[1] = 1'b0;
  assign io_out[0] = 1'b0;
  assign io_exceptionFlags[0] = 1'b0;
  assign io_exceptionFlags[1] = 1'b0;
  assign io_exceptionFlags[2] = 1'b0;
  assign io_exceptionFlags[3] = 1'b0;
  assign N3 = io_in[30] | io_in[31];
  assign N4 = io_in[29] | N3;
  assign N5 = ~N4;
  assign N6 = io_in[30] & io_in[31];
  assign T36 = { T46[11:11], T46[11:11], 1'b0, io_in[31:23] } + { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign io_out[51:29] = (N0)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N1)? io_in[22:0] : 1'b0;
  assign N0 = outRawFloat_isNaN;
  assign N1 = N2;
  assign io_exceptionFlags[4] = outRawFloat_isNaN & T1;
  assign T1 = ~io_in[22];
  assign outRawFloat_isNaN = N6 & io_in[29];
  assign N2 = ~outRawFloat_isNaN;
  assign io_out[63] = T20[11] | T19[11];
  assign io_out[62] = T20[10] | T19[11];
  assign io_out[61] = T20[9] | T19[11];
  assign io_out[60] = T20[8] | 1'b0;
  assign io_out[59] = T20[7] | 1'b0;
  assign io_out[58] = T20[6] | 1'b0;
  assign io_out[57] = T20[5] | 1'b0;
  assign io_out[56] = T20[4] | 1'b0;
  assign io_out[55] = T20[3] | 1'b0;
  assign io_out[54] = T20[2] | 1'b0;
  assign io_out[53] = T20[1] | 1'b0;
  assign io_out[52] = T20[0] | 1'b0;
  assign T19[11] = outRawFloat_isNaN;
  assign T20[11] = T26[11] | T21[11];
  assign T20[10] = T26[10] | T21[11];
  assign T20[9] = T26[9] | 1'b0;
  assign T20[8] = T26[8] | 1'b0;
  assign T20[7] = T26[7] | 1'b0;
  assign T20[6] = T26[6] | 1'b0;
  assign T20[5] = T26[5] | 1'b0;
  assign T20[4] = T26[4] | 1'b0;
  assign T20[3] = T26[3] | 1'b0;
  assign T20[2] = T26[2] | 1'b0;
  assign T20[1] = T26[1] | 1'b0;
  assign T20[0] = T26[0] | 1'b0;
  assign T21[11] = outRawFloat_isInf;
  assign outRawFloat_isInf = N6 & T24;
  assign T24 = ~io_in[29];
  assign T26[11] = T33[11] & T27[11];
  assign T26[10] = T33[10] & T27[10];
  assign T26[9] = T33[9] & T27[9];
  assign T26[8] = T33[8] & T27[8];
  assign T26[7] = T33[7] & T27[7];
  assign T26[6] = T33[6] & T27[6];
  assign T26[5] = T33[5] & T27[5];
  assign T26[4] = T33[4] & T27[4];
  assign T26[3] = T33[3] & T27[3];
  assign T26[2] = T33[2] & T27[2];
  assign T26[1] = T33[1] & T27[1];
  assign T26[0] = T33[0] & T27[0];
  assign T27[11] = ~1'b0;
  assign T27[10] = ~1'b0;
  assign T27[9] = ~T28[9];
  assign T27[8] = ~1'b0;
  assign T27[7] = ~1'b0;
  assign T27[6] = ~1'b0;
  assign T27[5] = ~1'b0;
  assign T27[4] = ~1'b0;
  assign T27[3] = ~1'b0;
  assign T27[2] = ~1'b0;
  assign T27[1] = ~1'b0;
  assign T27[0] = ~1'b0;
  assign T28[9] = T29;
  assign T29 = N5 | outRawFloat_isInf;
  assign T33[11] = T36[11] & T34[11];
  assign T33[10] = T36[10] & T34[10];
  assign T33[9] = T36[9] & T34[9];
  assign T33[8] = T36[8] & T34[8];
  assign T33[7] = T36[7] & T34[7];
  assign T33[6] = T36[6] & T34[6];
  assign T33[5] = T36[5] & T34[5];
  assign T33[4] = T36[4] & T34[4];
  assign T33[3] = T36[3] & T34[3];
  assign T33[2] = T36[2] & T34[2];
  assign T33[1] = T36[1] & T34[1];
  assign T33[0] = T36[0] & T34[0];
  assign T34[11] = ~T35[11];
  assign T34[10] = ~T35[11];
  assign T34[9] = ~1'b0;
  assign T34[8] = ~1'b0;
  assign T34[7] = ~1'b0;
  assign T34[6] = ~1'b0;
  assign T34[5] = ~1'b0;
  assign T34[4] = ~1'b0;
  assign T34[3] = ~1'b0;
  assign T34[2] = ~1'b0;
  assign T34[1] = ~1'b0;
  assign T34[0] = ~1'b0;
  assign T35[11] = N5;
  assign T46[11] = 1'b0;
  assign io_out[64] = io_in[32] & T42;
  assign T42 = ~outRawFloat_isNaN;

endmodule