module bsg_mem_1r1w_synth_width_p134_els_p16_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [3:0] w_addr_i;
  input [133:0] w_data_i;
  input [3:0] r_addr_i;
  output [133:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [133:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98;
  reg [2143:0] mem;
  assign r_data_o[133] = (N26)? mem[133] :
                         (N28)? mem[267] :
                         (N30)? mem[401] :
                         (N32)? mem[535] :
                         (N34)? mem[669] :
                         (N36)? mem[803] :
                         (N38)? mem[937] :
                         (N40)? mem[1071] :
                         (N27)? mem[1205] :
                         (N29)? mem[1339] :
                         (N31)? mem[1473] :
                         (N33)? mem[1607] :
                         (N35)? mem[1741] :
                         (N37)? mem[1875] :
                         (N39)? mem[2009] :
                         (N41)? mem[2143] : 1'b0;
  assign r_data_o[132] = (N26)? mem[132] :
                         (N28)? mem[266] :
                         (N30)? mem[400] :
                         (N32)? mem[534] :
                         (N34)? mem[668] :
                         (N36)? mem[802] :
                         (N38)? mem[936] :
                         (N40)? mem[1070] :
                         (N27)? mem[1204] :
                         (N29)? mem[1338] :
                         (N31)? mem[1472] :
                         (N33)? mem[1606] :
                         (N35)? mem[1740] :
                         (N37)? mem[1874] :
                         (N39)? mem[2008] :
                         (N41)? mem[2142] : 1'b0;
  assign r_data_o[131] = (N26)? mem[131] :
                         (N28)? mem[265] :
                         (N30)? mem[399] :
                         (N32)? mem[533] :
                         (N34)? mem[667] :
                         (N36)? mem[801] :
                         (N38)? mem[935] :
                         (N40)? mem[1069] :
                         (N27)? mem[1203] :
                         (N29)? mem[1337] :
                         (N31)? mem[1471] :
                         (N33)? mem[1605] :
                         (N35)? mem[1739] :
                         (N37)? mem[1873] :
                         (N39)? mem[2007] :
                         (N41)? mem[2141] : 1'b0;
  assign r_data_o[130] = (N26)? mem[130] :
                         (N28)? mem[264] :
                         (N30)? mem[398] :
                         (N32)? mem[532] :
                         (N34)? mem[666] :
                         (N36)? mem[800] :
                         (N38)? mem[934] :
                         (N40)? mem[1068] :
                         (N27)? mem[1202] :
                         (N29)? mem[1336] :
                         (N31)? mem[1470] :
                         (N33)? mem[1604] :
                         (N35)? mem[1738] :
                         (N37)? mem[1872] :
                         (N39)? mem[2006] :
                         (N41)? mem[2140] : 1'b0;
  assign r_data_o[129] = (N26)? mem[129] :
                         (N28)? mem[263] :
                         (N30)? mem[397] :
                         (N32)? mem[531] :
                         (N34)? mem[665] :
                         (N36)? mem[799] :
                         (N38)? mem[933] :
                         (N40)? mem[1067] :
                         (N27)? mem[1201] :
                         (N29)? mem[1335] :
                         (N31)? mem[1469] :
                         (N33)? mem[1603] :
                         (N35)? mem[1737] :
                         (N37)? mem[1871] :
                         (N39)? mem[2005] :
                         (N41)? mem[2139] : 1'b0;
  assign r_data_o[128] = (N26)? mem[128] :
                         (N28)? mem[262] :
                         (N30)? mem[396] :
                         (N32)? mem[530] :
                         (N34)? mem[664] :
                         (N36)? mem[798] :
                         (N38)? mem[932] :
                         (N40)? mem[1066] :
                         (N27)? mem[1200] :
                         (N29)? mem[1334] :
                         (N31)? mem[1468] :
                         (N33)? mem[1602] :
                         (N35)? mem[1736] :
                         (N37)? mem[1870] :
                         (N39)? mem[2004] :
                         (N41)? mem[2138] : 1'b0;
  assign r_data_o[127] = (N26)? mem[127] :
                         (N28)? mem[261] :
                         (N30)? mem[395] :
                         (N32)? mem[529] :
                         (N34)? mem[663] :
                         (N36)? mem[797] :
                         (N38)? mem[931] :
                         (N40)? mem[1065] :
                         (N27)? mem[1199] :
                         (N29)? mem[1333] :
                         (N31)? mem[1467] :
                         (N33)? mem[1601] :
                         (N35)? mem[1735] :
                         (N37)? mem[1869] :
                         (N39)? mem[2003] :
                         (N41)? mem[2137] : 1'b0;
  assign r_data_o[126] = (N26)? mem[126] :
                         (N28)? mem[260] :
                         (N30)? mem[394] :
                         (N32)? mem[528] :
                         (N34)? mem[662] :
                         (N36)? mem[796] :
                         (N38)? mem[930] :
                         (N40)? mem[1064] :
                         (N27)? mem[1198] :
                         (N29)? mem[1332] :
                         (N31)? mem[1466] :
                         (N33)? mem[1600] :
                         (N35)? mem[1734] :
                         (N37)? mem[1868] :
                         (N39)? mem[2002] :
                         (N41)? mem[2136] : 1'b0;
  assign r_data_o[125] = (N26)? mem[125] :
                         (N28)? mem[259] :
                         (N30)? mem[393] :
                         (N32)? mem[527] :
                         (N34)? mem[661] :
                         (N36)? mem[795] :
                         (N38)? mem[929] :
                         (N40)? mem[1063] :
                         (N27)? mem[1197] :
                         (N29)? mem[1331] :
                         (N31)? mem[1465] :
                         (N33)? mem[1599] :
                         (N35)? mem[1733] :
                         (N37)? mem[1867] :
                         (N39)? mem[2001] :
                         (N41)? mem[2135] : 1'b0;
  assign r_data_o[124] = (N26)? mem[124] :
                         (N28)? mem[258] :
                         (N30)? mem[392] :
                         (N32)? mem[526] :
                         (N34)? mem[660] :
                         (N36)? mem[794] :
                         (N38)? mem[928] :
                         (N40)? mem[1062] :
                         (N27)? mem[1196] :
                         (N29)? mem[1330] :
                         (N31)? mem[1464] :
                         (N33)? mem[1598] :
                         (N35)? mem[1732] :
                         (N37)? mem[1866] :
                         (N39)? mem[2000] :
                         (N41)? mem[2134] : 1'b0;
  assign r_data_o[123] = (N26)? mem[123] :
                         (N28)? mem[257] :
                         (N30)? mem[391] :
                         (N32)? mem[525] :
                         (N34)? mem[659] :
                         (N36)? mem[793] :
                         (N38)? mem[927] :
                         (N40)? mem[1061] :
                         (N27)? mem[1195] :
                         (N29)? mem[1329] :
                         (N31)? mem[1463] :
                         (N33)? mem[1597] :
                         (N35)? mem[1731] :
                         (N37)? mem[1865] :
                         (N39)? mem[1999] :
                         (N41)? mem[2133] : 1'b0;
  assign r_data_o[122] = (N26)? mem[122] :
                         (N28)? mem[256] :
                         (N30)? mem[390] :
                         (N32)? mem[524] :
                         (N34)? mem[658] :
                         (N36)? mem[792] :
                         (N38)? mem[926] :
                         (N40)? mem[1060] :
                         (N27)? mem[1194] :
                         (N29)? mem[1328] :
                         (N31)? mem[1462] :
                         (N33)? mem[1596] :
                         (N35)? mem[1730] :
                         (N37)? mem[1864] :
                         (N39)? mem[1998] :
                         (N41)? mem[2132] : 1'b0;
  assign r_data_o[121] = (N26)? mem[121] :
                         (N28)? mem[255] :
                         (N30)? mem[389] :
                         (N32)? mem[523] :
                         (N34)? mem[657] :
                         (N36)? mem[791] :
                         (N38)? mem[925] :
                         (N40)? mem[1059] :
                         (N27)? mem[1193] :
                         (N29)? mem[1327] :
                         (N31)? mem[1461] :
                         (N33)? mem[1595] :
                         (N35)? mem[1729] :
                         (N37)? mem[1863] :
                         (N39)? mem[1997] :
                         (N41)? mem[2131] : 1'b0;
  assign r_data_o[120] = (N26)? mem[120] :
                         (N28)? mem[254] :
                         (N30)? mem[388] :
                         (N32)? mem[522] :
                         (N34)? mem[656] :
                         (N36)? mem[790] :
                         (N38)? mem[924] :
                         (N40)? mem[1058] :
                         (N27)? mem[1192] :
                         (N29)? mem[1326] :
                         (N31)? mem[1460] :
                         (N33)? mem[1594] :
                         (N35)? mem[1728] :
                         (N37)? mem[1862] :
                         (N39)? mem[1996] :
                         (N41)? mem[2130] : 1'b0;
  assign r_data_o[119] = (N26)? mem[119] :
                         (N28)? mem[253] :
                         (N30)? mem[387] :
                         (N32)? mem[521] :
                         (N34)? mem[655] :
                         (N36)? mem[789] :
                         (N38)? mem[923] :
                         (N40)? mem[1057] :
                         (N27)? mem[1191] :
                         (N29)? mem[1325] :
                         (N31)? mem[1459] :
                         (N33)? mem[1593] :
                         (N35)? mem[1727] :
                         (N37)? mem[1861] :
                         (N39)? mem[1995] :
                         (N41)? mem[2129] : 1'b0;
  assign r_data_o[118] = (N26)? mem[118] :
                         (N28)? mem[252] :
                         (N30)? mem[386] :
                         (N32)? mem[520] :
                         (N34)? mem[654] :
                         (N36)? mem[788] :
                         (N38)? mem[922] :
                         (N40)? mem[1056] :
                         (N27)? mem[1190] :
                         (N29)? mem[1324] :
                         (N31)? mem[1458] :
                         (N33)? mem[1592] :
                         (N35)? mem[1726] :
                         (N37)? mem[1860] :
                         (N39)? mem[1994] :
                         (N41)? mem[2128] : 1'b0;
  assign r_data_o[117] = (N26)? mem[117] :
                         (N28)? mem[251] :
                         (N30)? mem[385] :
                         (N32)? mem[519] :
                         (N34)? mem[653] :
                         (N36)? mem[787] :
                         (N38)? mem[921] :
                         (N40)? mem[1055] :
                         (N27)? mem[1189] :
                         (N29)? mem[1323] :
                         (N31)? mem[1457] :
                         (N33)? mem[1591] :
                         (N35)? mem[1725] :
                         (N37)? mem[1859] :
                         (N39)? mem[1993] :
                         (N41)? mem[2127] : 1'b0;
  assign r_data_o[116] = (N26)? mem[116] :
                         (N28)? mem[250] :
                         (N30)? mem[384] :
                         (N32)? mem[518] :
                         (N34)? mem[652] :
                         (N36)? mem[786] :
                         (N38)? mem[920] :
                         (N40)? mem[1054] :
                         (N27)? mem[1188] :
                         (N29)? mem[1322] :
                         (N31)? mem[1456] :
                         (N33)? mem[1590] :
                         (N35)? mem[1724] :
                         (N37)? mem[1858] :
                         (N39)? mem[1992] :
                         (N41)? mem[2126] : 1'b0;
  assign r_data_o[115] = (N26)? mem[115] :
                         (N28)? mem[249] :
                         (N30)? mem[383] :
                         (N32)? mem[517] :
                         (N34)? mem[651] :
                         (N36)? mem[785] :
                         (N38)? mem[919] :
                         (N40)? mem[1053] :
                         (N27)? mem[1187] :
                         (N29)? mem[1321] :
                         (N31)? mem[1455] :
                         (N33)? mem[1589] :
                         (N35)? mem[1723] :
                         (N37)? mem[1857] :
                         (N39)? mem[1991] :
                         (N41)? mem[2125] : 1'b0;
  assign r_data_o[114] = (N26)? mem[114] :
                         (N28)? mem[248] :
                         (N30)? mem[382] :
                         (N32)? mem[516] :
                         (N34)? mem[650] :
                         (N36)? mem[784] :
                         (N38)? mem[918] :
                         (N40)? mem[1052] :
                         (N27)? mem[1186] :
                         (N29)? mem[1320] :
                         (N31)? mem[1454] :
                         (N33)? mem[1588] :
                         (N35)? mem[1722] :
                         (N37)? mem[1856] :
                         (N39)? mem[1990] :
                         (N41)? mem[2124] : 1'b0;
  assign r_data_o[113] = (N26)? mem[113] :
                         (N28)? mem[247] :
                         (N30)? mem[381] :
                         (N32)? mem[515] :
                         (N34)? mem[649] :
                         (N36)? mem[783] :
                         (N38)? mem[917] :
                         (N40)? mem[1051] :
                         (N27)? mem[1185] :
                         (N29)? mem[1319] :
                         (N31)? mem[1453] :
                         (N33)? mem[1587] :
                         (N35)? mem[1721] :
                         (N37)? mem[1855] :
                         (N39)? mem[1989] :
                         (N41)? mem[2123] : 1'b0;
  assign r_data_o[112] = (N26)? mem[112] :
                         (N28)? mem[246] :
                         (N30)? mem[380] :
                         (N32)? mem[514] :
                         (N34)? mem[648] :
                         (N36)? mem[782] :
                         (N38)? mem[916] :
                         (N40)? mem[1050] :
                         (N27)? mem[1184] :
                         (N29)? mem[1318] :
                         (N31)? mem[1452] :
                         (N33)? mem[1586] :
                         (N35)? mem[1720] :
                         (N37)? mem[1854] :
                         (N39)? mem[1988] :
                         (N41)? mem[2122] : 1'b0;
  assign r_data_o[111] = (N26)? mem[111] :
                         (N28)? mem[245] :
                         (N30)? mem[379] :
                         (N32)? mem[513] :
                         (N34)? mem[647] :
                         (N36)? mem[781] :
                         (N38)? mem[915] :
                         (N40)? mem[1049] :
                         (N27)? mem[1183] :
                         (N29)? mem[1317] :
                         (N31)? mem[1451] :
                         (N33)? mem[1585] :
                         (N35)? mem[1719] :
                         (N37)? mem[1853] :
                         (N39)? mem[1987] :
                         (N41)? mem[2121] : 1'b0;
  assign r_data_o[110] = (N26)? mem[110] :
                         (N28)? mem[244] :
                         (N30)? mem[378] :
                         (N32)? mem[512] :
                         (N34)? mem[646] :
                         (N36)? mem[780] :
                         (N38)? mem[914] :
                         (N40)? mem[1048] :
                         (N27)? mem[1182] :
                         (N29)? mem[1316] :
                         (N31)? mem[1450] :
                         (N33)? mem[1584] :
                         (N35)? mem[1718] :
                         (N37)? mem[1852] :
                         (N39)? mem[1986] :
                         (N41)? mem[2120] : 1'b0;
  assign r_data_o[109] = (N26)? mem[109] :
                         (N28)? mem[243] :
                         (N30)? mem[377] :
                         (N32)? mem[511] :
                         (N34)? mem[645] :
                         (N36)? mem[779] :
                         (N38)? mem[913] :
                         (N40)? mem[1047] :
                         (N27)? mem[1181] :
                         (N29)? mem[1315] :
                         (N31)? mem[1449] :
                         (N33)? mem[1583] :
                         (N35)? mem[1717] :
                         (N37)? mem[1851] :
                         (N39)? mem[1985] :
                         (N41)? mem[2119] : 1'b0;
  assign r_data_o[108] = (N26)? mem[108] :
                         (N28)? mem[242] :
                         (N30)? mem[376] :
                         (N32)? mem[510] :
                         (N34)? mem[644] :
                         (N36)? mem[778] :
                         (N38)? mem[912] :
                         (N40)? mem[1046] :
                         (N27)? mem[1180] :
                         (N29)? mem[1314] :
                         (N31)? mem[1448] :
                         (N33)? mem[1582] :
                         (N35)? mem[1716] :
                         (N37)? mem[1850] :
                         (N39)? mem[1984] :
                         (N41)? mem[2118] : 1'b0;
  assign r_data_o[107] = (N26)? mem[107] :
                         (N28)? mem[241] :
                         (N30)? mem[375] :
                         (N32)? mem[509] :
                         (N34)? mem[643] :
                         (N36)? mem[777] :
                         (N38)? mem[911] :
                         (N40)? mem[1045] :
                         (N27)? mem[1179] :
                         (N29)? mem[1313] :
                         (N31)? mem[1447] :
                         (N33)? mem[1581] :
                         (N35)? mem[1715] :
                         (N37)? mem[1849] :
                         (N39)? mem[1983] :
                         (N41)? mem[2117] : 1'b0;
  assign r_data_o[106] = (N26)? mem[106] :
                         (N28)? mem[240] :
                         (N30)? mem[374] :
                         (N32)? mem[508] :
                         (N34)? mem[642] :
                         (N36)? mem[776] :
                         (N38)? mem[910] :
                         (N40)? mem[1044] :
                         (N27)? mem[1178] :
                         (N29)? mem[1312] :
                         (N31)? mem[1446] :
                         (N33)? mem[1580] :
                         (N35)? mem[1714] :
                         (N37)? mem[1848] :
                         (N39)? mem[1982] :
                         (N41)? mem[2116] : 1'b0;
  assign r_data_o[105] = (N26)? mem[105] :
                         (N28)? mem[239] :
                         (N30)? mem[373] :
                         (N32)? mem[507] :
                         (N34)? mem[641] :
                         (N36)? mem[775] :
                         (N38)? mem[909] :
                         (N40)? mem[1043] :
                         (N27)? mem[1177] :
                         (N29)? mem[1311] :
                         (N31)? mem[1445] :
                         (N33)? mem[1579] :
                         (N35)? mem[1713] :
                         (N37)? mem[1847] :
                         (N39)? mem[1981] :
                         (N41)? mem[2115] : 1'b0;
  assign r_data_o[104] = (N26)? mem[104] :
                         (N28)? mem[238] :
                         (N30)? mem[372] :
                         (N32)? mem[506] :
                         (N34)? mem[640] :
                         (N36)? mem[774] :
                         (N38)? mem[908] :
                         (N40)? mem[1042] :
                         (N27)? mem[1176] :
                         (N29)? mem[1310] :
                         (N31)? mem[1444] :
                         (N33)? mem[1578] :
                         (N35)? mem[1712] :
                         (N37)? mem[1846] :
                         (N39)? mem[1980] :
                         (N41)? mem[2114] : 1'b0;
  assign r_data_o[103] = (N26)? mem[103] :
                         (N28)? mem[237] :
                         (N30)? mem[371] :
                         (N32)? mem[505] :
                         (N34)? mem[639] :
                         (N36)? mem[773] :
                         (N38)? mem[907] :
                         (N40)? mem[1041] :
                         (N27)? mem[1175] :
                         (N29)? mem[1309] :
                         (N31)? mem[1443] :
                         (N33)? mem[1577] :
                         (N35)? mem[1711] :
                         (N37)? mem[1845] :
                         (N39)? mem[1979] :
                         (N41)? mem[2113] : 1'b0;
  assign r_data_o[102] = (N26)? mem[102] :
                         (N28)? mem[236] :
                         (N30)? mem[370] :
                         (N32)? mem[504] :
                         (N34)? mem[638] :
                         (N36)? mem[772] :
                         (N38)? mem[906] :
                         (N40)? mem[1040] :
                         (N27)? mem[1174] :
                         (N29)? mem[1308] :
                         (N31)? mem[1442] :
                         (N33)? mem[1576] :
                         (N35)? mem[1710] :
                         (N37)? mem[1844] :
                         (N39)? mem[1978] :
                         (N41)? mem[2112] : 1'b0;
  assign r_data_o[101] = (N26)? mem[101] :
                         (N28)? mem[235] :
                         (N30)? mem[369] :
                         (N32)? mem[503] :
                         (N34)? mem[637] :
                         (N36)? mem[771] :
                         (N38)? mem[905] :
                         (N40)? mem[1039] :
                         (N27)? mem[1173] :
                         (N29)? mem[1307] :
                         (N31)? mem[1441] :
                         (N33)? mem[1575] :
                         (N35)? mem[1709] :
                         (N37)? mem[1843] :
                         (N39)? mem[1977] :
                         (N41)? mem[2111] : 1'b0;
  assign r_data_o[100] = (N26)? mem[100] :
                         (N28)? mem[234] :
                         (N30)? mem[368] :
                         (N32)? mem[502] :
                         (N34)? mem[636] :
                         (N36)? mem[770] :
                         (N38)? mem[904] :
                         (N40)? mem[1038] :
                         (N27)? mem[1172] :
                         (N29)? mem[1306] :
                         (N31)? mem[1440] :
                         (N33)? mem[1574] :
                         (N35)? mem[1708] :
                         (N37)? mem[1842] :
                         (N39)? mem[1976] :
                         (N41)? mem[2110] : 1'b0;
  assign r_data_o[99] = (N26)? mem[99] :
                        (N28)? mem[233] :
                        (N30)? mem[367] :
                        (N32)? mem[501] :
                        (N34)? mem[635] :
                        (N36)? mem[769] :
                        (N38)? mem[903] :
                        (N40)? mem[1037] :
                        (N27)? mem[1171] :
                        (N29)? mem[1305] :
                        (N31)? mem[1439] :
                        (N33)? mem[1573] :
                        (N35)? mem[1707] :
                        (N37)? mem[1841] :
                        (N39)? mem[1975] :
                        (N41)? mem[2109] : 1'b0;
  assign r_data_o[98] = (N26)? mem[98] :
                        (N28)? mem[232] :
                        (N30)? mem[366] :
                        (N32)? mem[500] :
                        (N34)? mem[634] :
                        (N36)? mem[768] :
                        (N38)? mem[902] :
                        (N40)? mem[1036] :
                        (N27)? mem[1170] :
                        (N29)? mem[1304] :
                        (N31)? mem[1438] :
                        (N33)? mem[1572] :
                        (N35)? mem[1706] :
                        (N37)? mem[1840] :
                        (N39)? mem[1974] :
                        (N41)? mem[2108] : 1'b0;
  assign r_data_o[97] = (N26)? mem[97] :
                        (N28)? mem[231] :
                        (N30)? mem[365] :
                        (N32)? mem[499] :
                        (N34)? mem[633] :
                        (N36)? mem[767] :
                        (N38)? mem[901] :
                        (N40)? mem[1035] :
                        (N27)? mem[1169] :
                        (N29)? mem[1303] :
                        (N31)? mem[1437] :
                        (N33)? mem[1571] :
                        (N35)? mem[1705] :
                        (N37)? mem[1839] :
                        (N39)? mem[1973] :
                        (N41)? mem[2107] : 1'b0;
  assign r_data_o[96] = (N26)? mem[96] :
                        (N28)? mem[230] :
                        (N30)? mem[364] :
                        (N32)? mem[498] :
                        (N34)? mem[632] :
                        (N36)? mem[766] :
                        (N38)? mem[900] :
                        (N40)? mem[1034] :
                        (N27)? mem[1168] :
                        (N29)? mem[1302] :
                        (N31)? mem[1436] :
                        (N33)? mem[1570] :
                        (N35)? mem[1704] :
                        (N37)? mem[1838] :
                        (N39)? mem[1972] :
                        (N41)? mem[2106] : 1'b0;
  assign r_data_o[95] = (N26)? mem[95] :
                        (N28)? mem[229] :
                        (N30)? mem[363] :
                        (N32)? mem[497] :
                        (N34)? mem[631] :
                        (N36)? mem[765] :
                        (N38)? mem[899] :
                        (N40)? mem[1033] :
                        (N27)? mem[1167] :
                        (N29)? mem[1301] :
                        (N31)? mem[1435] :
                        (N33)? mem[1569] :
                        (N35)? mem[1703] :
                        (N37)? mem[1837] :
                        (N39)? mem[1971] :
                        (N41)? mem[2105] : 1'b0;
  assign r_data_o[94] = (N26)? mem[94] :
                        (N28)? mem[228] :
                        (N30)? mem[362] :
                        (N32)? mem[496] :
                        (N34)? mem[630] :
                        (N36)? mem[764] :
                        (N38)? mem[898] :
                        (N40)? mem[1032] :
                        (N27)? mem[1166] :
                        (N29)? mem[1300] :
                        (N31)? mem[1434] :
                        (N33)? mem[1568] :
                        (N35)? mem[1702] :
                        (N37)? mem[1836] :
                        (N39)? mem[1970] :
                        (N41)? mem[2104] : 1'b0;
  assign r_data_o[93] = (N26)? mem[93] :
                        (N28)? mem[227] :
                        (N30)? mem[361] :
                        (N32)? mem[495] :
                        (N34)? mem[629] :
                        (N36)? mem[763] :
                        (N38)? mem[897] :
                        (N40)? mem[1031] :
                        (N27)? mem[1165] :
                        (N29)? mem[1299] :
                        (N31)? mem[1433] :
                        (N33)? mem[1567] :
                        (N35)? mem[1701] :
                        (N37)? mem[1835] :
                        (N39)? mem[1969] :
                        (N41)? mem[2103] : 1'b0;
  assign r_data_o[92] = (N26)? mem[92] :
                        (N28)? mem[226] :
                        (N30)? mem[360] :
                        (N32)? mem[494] :
                        (N34)? mem[628] :
                        (N36)? mem[762] :
                        (N38)? mem[896] :
                        (N40)? mem[1030] :
                        (N27)? mem[1164] :
                        (N29)? mem[1298] :
                        (N31)? mem[1432] :
                        (N33)? mem[1566] :
                        (N35)? mem[1700] :
                        (N37)? mem[1834] :
                        (N39)? mem[1968] :
                        (N41)? mem[2102] : 1'b0;
  assign r_data_o[91] = (N26)? mem[91] :
                        (N28)? mem[225] :
                        (N30)? mem[359] :
                        (N32)? mem[493] :
                        (N34)? mem[627] :
                        (N36)? mem[761] :
                        (N38)? mem[895] :
                        (N40)? mem[1029] :
                        (N27)? mem[1163] :
                        (N29)? mem[1297] :
                        (N31)? mem[1431] :
                        (N33)? mem[1565] :
                        (N35)? mem[1699] :
                        (N37)? mem[1833] :
                        (N39)? mem[1967] :
                        (N41)? mem[2101] : 1'b0;
  assign r_data_o[90] = (N26)? mem[90] :
                        (N28)? mem[224] :
                        (N30)? mem[358] :
                        (N32)? mem[492] :
                        (N34)? mem[626] :
                        (N36)? mem[760] :
                        (N38)? mem[894] :
                        (N40)? mem[1028] :
                        (N27)? mem[1162] :
                        (N29)? mem[1296] :
                        (N31)? mem[1430] :
                        (N33)? mem[1564] :
                        (N35)? mem[1698] :
                        (N37)? mem[1832] :
                        (N39)? mem[1966] :
                        (N41)? mem[2100] : 1'b0;
  assign r_data_o[89] = (N26)? mem[89] :
                        (N28)? mem[223] :
                        (N30)? mem[357] :
                        (N32)? mem[491] :
                        (N34)? mem[625] :
                        (N36)? mem[759] :
                        (N38)? mem[893] :
                        (N40)? mem[1027] :
                        (N27)? mem[1161] :
                        (N29)? mem[1295] :
                        (N31)? mem[1429] :
                        (N33)? mem[1563] :
                        (N35)? mem[1697] :
                        (N37)? mem[1831] :
                        (N39)? mem[1965] :
                        (N41)? mem[2099] : 1'b0;
  assign r_data_o[88] = (N26)? mem[88] :
                        (N28)? mem[222] :
                        (N30)? mem[356] :
                        (N32)? mem[490] :
                        (N34)? mem[624] :
                        (N36)? mem[758] :
                        (N38)? mem[892] :
                        (N40)? mem[1026] :
                        (N27)? mem[1160] :
                        (N29)? mem[1294] :
                        (N31)? mem[1428] :
                        (N33)? mem[1562] :
                        (N35)? mem[1696] :
                        (N37)? mem[1830] :
                        (N39)? mem[1964] :
                        (N41)? mem[2098] : 1'b0;
  assign r_data_o[87] = (N26)? mem[87] :
                        (N28)? mem[221] :
                        (N30)? mem[355] :
                        (N32)? mem[489] :
                        (N34)? mem[623] :
                        (N36)? mem[757] :
                        (N38)? mem[891] :
                        (N40)? mem[1025] :
                        (N27)? mem[1159] :
                        (N29)? mem[1293] :
                        (N31)? mem[1427] :
                        (N33)? mem[1561] :
                        (N35)? mem[1695] :
                        (N37)? mem[1829] :
                        (N39)? mem[1963] :
                        (N41)? mem[2097] : 1'b0;
  assign r_data_o[86] = (N26)? mem[86] :
                        (N28)? mem[220] :
                        (N30)? mem[354] :
                        (N32)? mem[488] :
                        (N34)? mem[622] :
                        (N36)? mem[756] :
                        (N38)? mem[890] :
                        (N40)? mem[1024] :
                        (N27)? mem[1158] :
                        (N29)? mem[1292] :
                        (N31)? mem[1426] :
                        (N33)? mem[1560] :
                        (N35)? mem[1694] :
                        (N37)? mem[1828] :
                        (N39)? mem[1962] :
                        (N41)? mem[2096] : 1'b0;
  assign r_data_o[85] = (N26)? mem[85] :
                        (N28)? mem[219] :
                        (N30)? mem[353] :
                        (N32)? mem[487] :
                        (N34)? mem[621] :
                        (N36)? mem[755] :
                        (N38)? mem[889] :
                        (N40)? mem[1023] :
                        (N27)? mem[1157] :
                        (N29)? mem[1291] :
                        (N31)? mem[1425] :
                        (N33)? mem[1559] :
                        (N35)? mem[1693] :
                        (N37)? mem[1827] :
                        (N39)? mem[1961] :
                        (N41)? mem[2095] : 1'b0;
  assign r_data_o[84] = (N26)? mem[84] :
                        (N28)? mem[218] :
                        (N30)? mem[352] :
                        (N32)? mem[486] :
                        (N34)? mem[620] :
                        (N36)? mem[754] :
                        (N38)? mem[888] :
                        (N40)? mem[1022] :
                        (N27)? mem[1156] :
                        (N29)? mem[1290] :
                        (N31)? mem[1424] :
                        (N33)? mem[1558] :
                        (N35)? mem[1692] :
                        (N37)? mem[1826] :
                        (N39)? mem[1960] :
                        (N41)? mem[2094] : 1'b0;
  assign r_data_o[83] = (N26)? mem[83] :
                        (N28)? mem[217] :
                        (N30)? mem[351] :
                        (N32)? mem[485] :
                        (N34)? mem[619] :
                        (N36)? mem[753] :
                        (N38)? mem[887] :
                        (N40)? mem[1021] :
                        (N27)? mem[1155] :
                        (N29)? mem[1289] :
                        (N31)? mem[1423] :
                        (N33)? mem[1557] :
                        (N35)? mem[1691] :
                        (N37)? mem[1825] :
                        (N39)? mem[1959] :
                        (N41)? mem[2093] : 1'b0;
  assign r_data_o[82] = (N26)? mem[82] :
                        (N28)? mem[216] :
                        (N30)? mem[350] :
                        (N32)? mem[484] :
                        (N34)? mem[618] :
                        (N36)? mem[752] :
                        (N38)? mem[886] :
                        (N40)? mem[1020] :
                        (N27)? mem[1154] :
                        (N29)? mem[1288] :
                        (N31)? mem[1422] :
                        (N33)? mem[1556] :
                        (N35)? mem[1690] :
                        (N37)? mem[1824] :
                        (N39)? mem[1958] :
                        (N41)? mem[2092] : 1'b0;
  assign r_data_o[81] = (N26)? mem[81] :
                        (N28)? mem[215] :
                        (N30)? mem[349] :
                        (N32)? mem[483] :
                        (N34)? mem[617] :
                        (N36)? mem[751] :
                        (N38)? mem[885] :
                        (N40)? mem[1019] :
                        (N27)? mem[1153] :
                        (N29)? mem[1287] :
                        (N31)? mem[1421] :
                        (N33)? mem[1555] :
                        (N35)? mem[1689] :
                        (N37)? mem[1823] :
                        (N39)? mem[1957] :
                        (N41)? mem[2091] : 1'b0;
  assign r_data_o[80] = (N26)? mem[80] :
                        (N28)? mem[214] :
                        (N30)? mem[348] :
                        (N32)? mem[482] :
                        (N34)? mem[616] :
                        (N36)? mem[750] :
                        (N38)? mem[884] :
                        (N40)? mem[1018] :
                        (N27)? mem[1152] :
                        (N29)? mem[1286] :
                        (N31)? mem[1420] :
                        (N33)? mem[1554] :
                        (N35)? mem[1688] :
                        (N37)? mem[1822] :
                        (N39)? mem[1956] :
                        (N41)? mem[2090] : 1'b0;
  assign r_data_o[79] = (N26)? mem[79] :
                        (N28)? mem[213] :
                        (N30)? mem[347] :
                        (N32)? mem[481] :
                        (N34)? mem[615] :
                        (N36)? mem[749] :
                        (N38)? mem[883] :
                        (N40)? mem[1017] :
                        (N27)? mem[1151] :
                        (N29)? mem[1285] :
                        (N31)? mem[1419] :
                        (N33)? mem[1553] :
                        (N35)? mem[1687] :
                        (N37)? mem[1821] :
                        (N39)? mem[1955] :
                        (N41)? mem[2089] : 1'b0;
  assign r_data_o[78] = (N26)? mem[78] :
                        (N28)? mem[212] :
                        (N30)? mem[346] :
                        (N32)? mem[480] :
                        (N34)? mem[614] :
                        (N36)? mem[748] :
                        (N38)? mem[882] :
                        (N40)? mem[1016] :
                        (N27)? mem[1150] :
                        (N29)? mem[1284] :
                        (N31)? mem[1418] :
                        (N33)? mem[1552] :
                        (N35)? mem[1686] :
                        (N37)? mem[1820] :
                        (N39)? mem[1954] :
                        (N41)? mem[2088] : 1'b0;
  assign r_data_o[77] = (N26)? mem[77] :
                        (N28)? mem[211] :
                        (N30)? mem[345] :
                        (N32)? mem[479] :
                        (N34)? mem[613] :
                        (N36)? mem[747] :
                        (N38)? mem[881] :
                        (N40)? mem[1015] :
                        (N27)? mem[1149] :
                        (N29)? mem[1283] :
                        (N31)? mem[1417] :
                        (N33)? mem[1551] :
                        (N35)? mem[1685] :
                        (N37)? mem[1819] :
                        (N39)? mem[1953] :
                        (N41)? mem[2087] : 1'b0;
  assign r_data_o[76] = (N26)? mem[76] :
                        (N28)? mem[210] :
                        (N30)? mem[344] :
                        (N32)? mem[478] :
                        (N34)? mem[612] :
                        (N36)? mem[746] :
                        (N38)? mem[880] :
                        (N40)? mem[1014] :
                        (N27)? mem[1148] :
                        (N29)? mem[1282] :
                        (N31)? mem[1416] :
                        (N33)? mem[1550] :
                        (N35)? mem[1684] :
                        (N37)? mem[1818] :
                        (N39)? mem[1952] :
                        (N41)? mem[2086] : 1'b0;
  assign r_data_o[75] = (N26)? mem[75] :
                        (N28)? mem[209] :
                        (N30)? mem[343] :
                        (N32)? mem[477] :
                        (N34)? mem[611] :
                        (N36)? mem[745] :
                        (N38)? mem[879] :
                        (N40)? mem[1013] :
                        (N27)? mem[1147] :
                        (N29)? mem[1281] :
                        (N31)? mem[1415] :
                        (N33)? mem[1549] :
                        (N35)? mem[1683] :
                        (N37)? mem[1817] :
                        (N39)? mem[1951] :
                        (N41)? mem[2085] : 1'b0;
  assign r_data_o[74] = (N26)? mem[74] :
                        (N28)? mem[208] :
                        (N30)? mem[342] :
                        (N32)? mem[476] :
                        (N34)? mem[610] :
                        (N36)? mem[744] :
                        (N38)? mem[878] :
                        (N40)? mem[1012] :
                        (N27)? mem[1146] :
                        (N29)? mem[1280] :
                        (N31)? mem[1414] :
                        (N33)? mem[1548] :
                        (N35)? mem[1682] :
                        (N37)? mem[1816] :
                        (N39)? mem[1950] :
                        (N41)? mem[2084] : 1'b0;
  assign r_data_o[73] = (N26)? mem[73] :
                        (N28)? mem[207] :
                        (N30)? mem[341] :
                        (N32)? mem[475] :
                        (N34)? mem[609] :
                        (N36)? mem[743] :
                        (N38)? mem[877] :
                        (N40)? mem[1011] :
                        (N27)? mem[1145] :
                        (N29)? mem[1279] :
                        (N31)? mem[1413] :
                        (N33)? mem[1547] :
                        (N35)? mem[1681] :
                        (N37)? mem[1815] :
                        (N39)? mem[1949] :
                        (N41)? mem[2083] : 1'b0;
  assign r_data_o[72] = (N26)? mem[72] :
                        (N28)? mem[206] :
                        (N30)? mem[340] :
                        (N32)? mem[474] :
                        (N34)? mem[608] :
                        (N36)? mem[742] :
                        (N38)? mem[876] :
                        (N40)? mem[1010] :
                        (N27)? mem[1144] :
                        (N29)? mem[1278] :
                        (N31)? mem[1412] :
                        (N33)? mem[1546] :
                        (N35)? mem[1680] :
                        (N37)? mem[1814] :
                        (N39)? mem[1948] :
                        (N41)? mem[2082] : 1'b0;
  assign r_data_o[71] = (N26)? mem[71] :
                        (N28)? mem[205] :
                        (N30)? mem[339] :
                        (N32)? mem[473] :
                        (N34)? mem[607] :
                        (N36)? mem[741] :
                        (N38)? mem[875] :
                        (N40)? mem[1009] :
                        (N27)? mem[1143] :
                        (N29)? mem[1277] :
                        (N31)? mem[1411] :
                        (N33)? mem[1545] :
                        (N35)? mem[1679] :
                        (N37)? mem[1813] :
                        (N39)? mem[1947] :
                        (N41)? mem[2081] : 1'b0;
  assign r_data_o[70] = (N26)? mem[70] :
                        (N28)? mem[204] :
                        (N30)? mem[338] :
                        (N32)? mem[472] :
                        (N34)? mem[606] :
                        (N36)? mem[740] :
                        (N38)? mem[874] :
                        (N40)? mem[1008] :
                        (N27)? mem[1142] :
                        (N29)? mem[1276] :
                        (N31)? mem[1410] :
                        (N33)? mem[1544] :
                        (N35)? mem[1678] :
                        (N37)? mem[1812] :
                        (N39)? mem[1946] :
                        (N41)? mem[2080] : 1'b0;
  assign r_data_o[69] = (N26)? mem[69] :
                        (N28)? mem[203] :
                        (N30)? mem[337] :
                        (N32)? mem[471] :
                        (N34)? mem[605] :
                        (N36)? mem[739] :
                        (N38)? mem[873] :
                        (N40)? mem[1007] :
                        (N27)? mem[1141] :
                        (N29)? mem[1275] :
                        (N31)? mem[1409] :
                        (N33)? mem[1543] :
                        (N35)? mem[1677] :
                        (N37)? mem[1811] :
                        (N39)? mem[1945] :
                        (N41)? mem[2079] : 1'b0;
  assign r_data_o[68] = (N26)? mem[68] :
                        (N28)? mem[202] :
                        (N30)? mem[336] :
                        (N32)? mem[470] :
                        (N34)? mem[604] :
                        (N36)? mem[738] :
                        (N38)? mem[872] :
                        (N40)? mem[1006] :
                        (N27)? mem[1140] :
                        (N29)? mem[1274] :
                        (N31)? mem[1408] :
                        (N33)? mem[1542] :
                        (N35)? mem[1676] :
                        (N37)? mem[1810] :
                        (N39)? mem[1944] :
                        (N41)? mem[2078] : 1'b0;
  assign r_data_o[67] = (N26)? mem[67] :
                        (N28)? mem[201] :
                        (N30)? mem[335] :
                        (N32)? mem[469] :
                        (N34)? mem[603] :
                        (N36)? mem[737] :
                        (N38)? mem[871] :
                        (N40)? mem[1005] :
                        (N27)? mem[1139] :
                        (N29)? mem[1273] :
                        (N31)? mem[1407] :
                        (N33)? mem[1541] :
                        (N35)? mem[1675] :
                        (N37)? mem[1809] :
                        (N39)? mem[1943] :
                        (N41)? mem[2077] : 1'b0;
  assign r_data_o[66] = (N26)? mem[66] :
                        (N28)? mem[200] :
                        (N30)? mem[334] :
                        (N32)? mem[468] :
                        (N34)? mem[602] :
                        (N36)? mem[736] :
                        (N38)? mem[870] :
                        (N40)? mem[1004] :
                        (N27)? mem[1138] :
                        (N29)? mem[1272] :
                        (N31)? mem[1406] :
                        (N33)? mem[1540] :
                        (N35)? mem[1674] :
                        (N37)? mem[1808] :
                        (N39)? mem[1942] :
                        (N41)? mem[2076] : 1'b0;
  assign r_data_o[65] = (N26)? mem[65] :
                        (N28)? mem[199] :
                        (N30)? mem[333] :
                        (N32)? mem[467] :
                        (N34)? mem[601] :
                        (N36)? mem[735] :
                        (N38)? mem[869] :
                        (N40)? mem[1003] :
                        (N27)? mem[1137] :
                        (N29)? mem[1271] :
                        (N31)? mem[1405] :
                        (N33)? mem[1539] :
                        (N35)? mem[1673] :
                        (N37)? mem[1807] :
                        (N39)? mem[1941] :
                        (N41)? mem[2075] : 1'b0;
  assign r_data_o[64] = (N26)? mem[64] :
                        (N28)? mem[198] :
                        (N30)? mem[332] :
                        (N32)? mem[466] :
                        (N34)? mem[600] :
                        (N36)? mem[734] :
                        (N38)? mem[868] :
                        (N40)? mem[1002] :
                        (N27)? mem[1136] :
                        (N29)? mem[1270] :
                        (N31)? mem[1404] :
                        (N33)? mem[1538] :
                        (N35)? mem[1672] :
                        (N37)? mem[1806] :
                        (N39)? mem[1940] :
                        (N41)? mem[2074] : 1'b0;
  assign r_data_o[63] = (N26)? mem[63] :
                        (N28)? mem[197] :
                        (N30)? mem[331] :
                        (N32)? mem[465] :
                        (N34)? mem[599] :
                        (N36)? mem[733] :
                        (N38)? mem[867] :
                        (N40)? mem[1001] :
                        (N27)? mem[1135] :
                        (N29)? mem[1269] :
                        (N31)? mem[1403] :
                        (N33)? mem[1537] :
                        (N35)? mem[1671] :
                        (N37)? mem[1805] :
                        (N39)? mem[1939] :
                        (N41)? mem[2073] : 1'b0;
  assign r_data_o[62] = (N26)? mem[62] :
                        (N28)? mem[196] :
                        (N30)? mem[330] :
                        (N32)? mem[464] :
                        (N34)? mem[598] :
                        (N36)? mem[732] :
                        (N38)? mem[866] :
                        (N40)? mem[1000] :
                        (N27)? mem[1134] :
                        (N29)? mem[1268] :
                        (N31)? mem[1402] :
                        (N33)? mem[1536] :
                        (N35)? mem[1670] :
                        (N37)? mem[1804] :
                        (N39)? mem[1938] :
                        (N41)? mem[2072] : 1'b0;
  assign r_data_o[61] = (N26)? mem[61] :
                        (N28)? mem[195] :
                        (N30)? mem[329] :
                        (N32)? mem[463] :
                        (N34)? mem[597] :
                        (N36)? mem[731] :
                        (N38)? mem[865] :
                        (N40)? mem[999] :
                        (N27)? mem[1133] :
                        (N29)? mem[1267] :
                        (N31)? mem[1401] :
                        (N33)? mem[1535] :
                        (N35)? mem[1669] :
                        (N37)? mem[1803] :
                        (N39)? mem[1937] :
                        (N41)? mem[2071] : 1'b0;
  assign r_data_o[60] = (N26)? mem[60] :
                        (N28)? mem[194] :
                        (N30)? mem[328] :
                        (N32)? mem[462] :
                        (N34)? mem[596] :
                        (N36)? mem[730] :
                        (N38)? mem[864] :
                        (N40)? mem[998] :
                        (N27)? mem[1132] :
                        (N29)? mem[1266] :
                        (N31)? mem[1400] :
                        (N33)? mem[1534] :
                        (N35)? mem[1668] :
                        (N37)? mem[1802] :
                        (N39)? mem[1936] :
                        (N41)? mem[2070] : 1'b0;
  assign r_data_o[59] = (N26)? mem[59] :
                        (N28)? mem[193] :
                        (N30)? mem[327] :
                        (N32)? mem[461] :
                        (N34)? mem[595] :
                        (N36)? mem[729] :
                        (N38)? mem[863] :
                        (N40)? mem[997] :
                        (N27)? mem[1131] :
                        (N29)? mem[1265] :
                        (N31)? mem[1399] :
                        (N33)? mem[1533] :
                        (N35)? mem[1667] :
                        (N37)? mem[1801] :
                        (N39)? mem[1935] :
                        (N41)? mem[2069] : 1'b0;
  assign r_data_o[58] = (N26)? mem[58] :
                        (N28)? mem[192] :
                        (N30)? mem[326] :
                        (N32)? mem[460] :
                        (N34)? mem[594] :
                        (N36)? mem[728] :
                        (N38)? mem[862] :
                        (N40)? mem[996] :
                        (N27)? mem[1130] :
                        (N29)? mem[1264] :
                        (N31)? mem[1398] :
                        (N33)? mem[1532] :
                        (N35)? mem[1666] :
                        (N37)? mem[1800] :
                        (N39)? mem[1934] :
                        (N41)? mem[2068] : 1'b0;
  assign r_data_o[57] = (N26)? mem[57] :
                        (N28)? mem[191] :
                        (N30)? mem[325] :
                        (N32)? mem[459] :
                        (N34)? mem[593] :
                        (N36)? mem[727] :
                        (N38)? mem[861] :
                        (N40)? mem[995] :
                        (N27)? mem[1129] :
                        (N29)? mem[1263] :
                        (N31)? mem[1397] :
                        (N33)? mem[1531] :
                        (N35)? mem[1665] :
                        (N37)? mem[1799] :
                        (N39)? mem[1933] :
                        (N41)? mem[2067] : 1'b0;
  assign r_data_o[56] = (N26)? mem[56] :
                        (N28)? mem[190] :
                        (N30)? mem[324] :
                        (N32)? mem[458] :
                        (N34)? mem[592] :
                        (N36)? mem[726] :
                        (N38)? mem[860] :
                        (N40)? mem[994] :
                        (N27)? mem[1128] :
                        (N29)? mem[1262] :
                        (N31)? mem[1396] :
                        (N33)? mem[1530] :
                        (N35)? mem[1664] :
                        (N37)? mem[1798] :
                        (N39)? mem[1932] :
                        (N41)? mem[2066] : 1'b0;
  assign r_data_o[55] = (N26)? mem[55] :
                        (N28)? mem[189] :
                        (N30)? mem[323] :
                        (N32)? mem[457] :
                        (N34)? mem[591] :
                        (N36)? mem[725] :
                        (N38)? mem[859] :
                        (N40)? mem[993] :
                        (N27)? mem[1127] :
                        (N29)? mem[1261] :
                        (N31)? mem[1395] :
                        (N33)? mem[1529] :
                        (N35)? mem[1663] :
                        (N37)? mem[1797] :
                        (N39)? mem[1931] :
                        (N41)? mem[2065] : 1'b0;
  assign r_data_o[54] = (N26)? mem[54] :
                        (N28)? mem[188] :
                        (N30)? mem[322] :
                        (N32)? mem[456] :
                        (N34)? mem[590] :
                        (N36)? mem[724] :
                        (N38)? mem[858] :
                        (N40)? mem[992] :
                        (N27)? mem[1126] :
                        (N29)? mem[1260] :
                        (N31)? mem[1394] :
                        (N33)? mem[1528] :
                        (N35)? mem[1662] :
                        (N37)? mem[1796] :
                        (N39)? mem[1930] :
                        (N41)? mem[2064] : 1'b0;
  assign r_data_o[53] = (N26)? mem[53] :
                        (N28)? mem[187] :
                        (N30)? mem[321] :
                        (N32)? mem[455] :
                        (N34)? mem[589] :
                        (N36)? mem[723] :
                        (N38)? mem[857] :
                        (N40)? mem[991] :
                        (N27)? mem[1125] :
                        (N29)? mem[1259] :
                        (N31)? mem[1393] :
                        (N33)? mem[1527] :
                        (N35)? mem[1661] :
                        (N37)? mem[1795] :
                        (N39)? mem[1929] :
                        (N41)? mem[2063] : 1'b0;
  assign r_data_o[52] = (N26)? mem[52] :
                        (N28)? mem[186] :
                        (N30)? mem[320] :
                        (N32)? mem[454] :
                        (N34)? mem[588] :
                        (N36)? mem[722] :
                        (N38)? mem[856] :
                        (N40)? mem[990] :
                        (N27)? mem[1124] :
                        (N29)? mem[1258] :
                        (N31)? mem[1392] :
                        (N33)? mem[1526] :
                        (N35)? mem[1660] :
                        (N37)? mem[1794] :
                        (N39)? mem[1928] :
                        (N41)? mem[2062] : 1'b0;
  assign r_data_o[51] = (N26)? mem[51] :
                        (N28)? mem[185] :
                        (N30)? mem[319] :
                        (N32)? mem[453] :
                        (N34)? mem[587] :
                        (N36)? mem[721] :
                        (N38)? mem[855] :
                        (N40)? mem[989] :
                        (N27)? mem[1123] :
                        (N29)? mem[1257] :
                        (N31)? mem[1391] :
                        (N33)? mem[1525] :
                        (N35)? mem[1659] :
                        (N37)? mem[1793] :
                        (N39)? mem[1927] :
                        (N41)? mem[2061] : 1'b0;
  assign r_data_o[50] = (N26)? mem[50] :
                        (N28)? mem[184] :
                        (N30)? mem[318] :
                        (N32)? mem[452] :
                        (N34)? mem[586] :
                        (N36)? mem[720] :
                        (N38)? mem[854] :
                        (N40)? mem[988] :
                        (N27)? mem[1122] :
                        (N29)? mem[1256] :
                        (N31)? mem[1390] :
                        (N33)? mem[1524] :
                        (N35)? mem[1658] :
                        (N37)? mem[1792] :
                        (N39)? mem[1926] :
                        (N41)? mem[2060] : 1'b0;
  assign r_data_o[49] = (N26)? mem[49] :
                        (N28)? mem[183] :
                        (N30)? mem[317] :
                        (N32)? mem[451] :
                        (N34)? mem[585] :
                        (N36)? mem[719] :
                        (N38)? mem[853] :
                        (N40)? mem[987] :
                        (N27)? mem[1121] :
                        (N29)? mem[1255] :
                        (N31)? mem[1389] :
                        (N33)? mem[1523] :
                        (N35)? mem[1657] :
                        (N37)? mem[1791] :
                        (N39)? mem[1925] :
                        (N41)? mem[2059] : 1'b0;
  assign r_data_o[48] = (N26)? mem[48] :
                        (N28)? mem[182] :
                        (N30)? mem[316] :
                        (N32)? mem[450] :
                        (N34)? mem[584] :
                        (N36)? mem[718] :
                        (N38)? mem[852] :
                        (N40)? mem[986] :
                        (N27)? mem[1120] :
                        (N29)? mem[1254] :
                        (N31)? mem[1388] :
                        (N33)? mem[1522] :
                        (N35)? mem[1656] :
                        (N37)? mem[1790] :
                        (N39)? mem[1924] :
                        (N41)? mem[2058] : 1'b0;
  assign r_data_o[47] = (N26)? mem[47] :
                        (N28)? mem[181] :
                        (N30)? mem[315] :
                        (N32)? mem[449] :
                        (N34)? mem[583] :
                        (N36)? mem[717] :
                        (N38)? mem[851] :
                        (N40)? mem[985] :
                        (N27)? mem[1119] :
                        (N29)? mem[1253] :
                        (N31)? mem[1387] :
                        (N33)? mem[1521] :
                        (N35)? mem[1655] :
                        (N37)? mem[1789] :
                        (N39)? mem[1923] :
                        (N41)? mem[2057] : 1'b0;
  assign r_data_o[46] = (N26)? mem[46] :
                        (N28)? mem[180] :
                        (N30)? mem[314] :
                        (N32)? mem[448] :
                        (N34)? mem[582] :
                        (N36)? mem[716] :
                        (N38)? mem[850] :
                        (N40)? mem[984] :
                        (N27)? mem[1118] :
                        (N29)? mem[1252] :
                        (N31)? mem[1386] :
                        (N33)? mem[1520] :
                        (N35)? mem[1654] :
                        (N37)? mem[1788] :
                        (N39)? mem[1922] :
                        (N41)? mem[2056] : 1'b0;
  assign r_data_o[45] = (N26)? mem[45] :
                        (N28)? mem[179] :
                        (N30)? mem[313] :
                        (N32)? mem[447] :
                        (N34)? mem[581] :
                        (N36)? mem[715] :
                        (N38)? mem[849] :
                        (N40)? mem[983] :
                        (N27)? mem[1117] :
                        (N29)? mem[1251] :
                        (N31)? mem[1385] :
                        (N33)? mem[1519] :
                        (N35)? mem[1653] :
                        (N37)? mem[1787] :
                        (N39)? mem[1921] :
                        (N41)? mem[2055] : 1'b0;
  assign r_data_o[44] = (N26)? mem[44] :
                        (N28)? mem[178] :
                        (N30)? mem[312] :
                        (N32)? mem[446] :
                        (N34)? mem[580] :
                        (N36)? mem[714] :
                        (N38)? mem[848] :
                        (N40)? mem[982] :
                        (N27)? mem[1116] :
                        (N29)? mem[1250] :
                        (N31)? mem[1384] :
                        (N33)? mem[1518] :
                        (N35)? mem[1652] :
                        (N37)? mem[1786] :
                        (N39)? mem[1920] :
                        (N41)? mem[2054] : 1'b0;
  assign r_data_o[43] = (N26)? mem[43] :
                        (N28)? mem[177] :
                        (N30)? mem[311] :
                        (N32)? mem[445] :
                        (N34)? mem[579] :
                        (N36)? mem[713] :
                        (N38)? mem[847] :
                        (N40)? mem[981] :
                        (N27)? mem[1115] :
                        (N29)? mem[1249] :
                        (N31)? mem[1383] :
                        (N33)? mem[1517] :
                        (N35)? mem[1651] :
                        (N37)? mem[1785] :
                        (N39)? mem[1919] :
                        (N41)? mem[2053] : 1'b0;
  assign r_data_o[42] = (N26)? mem[42] :
                        (N28)? mem[176] :
                        (N30)? mem[310] :
                        (N32)? mem[444] :
                        (N34)? mem[578] :
                        (N36)? mem[712] :
                        (N38)? mem[846] :
                        (N40)? mem[980] :
                        (N27)? mem[1114] :
                        (N29)? mem[1248] :
                        (N31)? mem[1382] :
                        (N33)? mem[1516] :
                        (N35)? mem[1650] :
                        (N37)? mem[1784] :
                        (N39)? mem[1918] :
                        (N41)? mem[2052] : 1'b0;
  assign r_data_o[41] = (N26)? mem[41] :
                        (N28)? mem[175] :
                        (N30)? mem[309] :
                        (N32)? mem[443] :
                        (N34)? mem[577] :
                        (N36)? mem[711] :
                        (N38)? mem[845] :
                        (N40)? mem[979] :
                        (N27)? mem[1113] :
                        (N29)? mem[1247] :
                        (N31)? mem[1381] :
                        (N33)? mem[1515] :
                        (N35)? mem[1649] :
                        (N37)? mem[1783] :
                        (N39)? mem[1917] :
                        (N41)? mem[2051] : 1'b0;
  assign r_data_o[40] = (N26)? mem[40] :
                        (N28)? mem[174] :
                        (N30)? mem[308] :
                        (N32)? mem[442] :
                        (N34)? mem[576] :
                        (N36)? mem[710] :
                        (N38)? mem[844] :
                        (N40)? mem[978] :
                        (N27)? mem[1112] :
                        (N29)? mem[1246] :
                        (N31)? mem[1380] :
                        (N33)? mem[1514] :
                        (N35)? mem[1648] :
                        (N37)? mem[1782] :
                        (N39)? mem[1916] :
                        (N41)? mem[2050] : 1'b0;
  assign r_data_o[39] = (N26)? mem[39] :
                        (N28)? mem[173] :
                        (N30)? mem[307] :
                        (N32)? mem[441] :
                        (N34)? mem[575] :
                        (N36)? mem[709] :
                        (N38)? mem[843] :
                        (N40)? mem[977] :
                        (N27)? mem[1111] :
                        (N29)? mem[1245] :
                        (N31)? mem[1379] :
                        (N33)? mem[1513] :
                        (N35)? mem[1647] :
                        (N37)? mem[1781] :
                        (N39)? mem[1915] :
                        (N41)? mem[2049] : 1'b0;
  assign r_data_o[38] = (N26)? mem[38] :
                        (N28)? mem[172] :
                        (N30)? mem[306] :
                        (N32)? mem[440] :
                        (N34)? mem[574] :
                        (N36)? mem[708] :
                        (N38)? mem[842] :
                        (N40)? mem[976] :
                        (N27)? mem[1110] :
                        (N29)? mem[1244] :
                        (N31)? mem[1378] :
                        (N33)? mem[1512] :
                        (N35)? mem[1646] :
                        (N37)? mem[1780] :
                        (N39)? mem[1914] :
                        (N41)? mem[2048] : 1'b0;
  assign r_data_o[37] = (N26)? mem[37] :
                        (N28)? mem[171] :
                        (N30)? mem[305] :
                        (N32)? mem[439] :
                        (N34)? mem[573] :
                        (N36)? mem[707] :
                        (N38)? mem[841] :
                        (N40)? mem[975] :
                        (N27)? mem[1109] :
                        (N29)? mem[1243] :
                        (N31)? mem[1377] :
                        (N33)? mem[1511] :
                        (N35)? mem[1645] :
                        (N37)? mem[1779] :
                        (N39)? mem[1913] :
                        (N41)? mem[2047] : 1'b0;
  assign r_data_o[36] = (N26)? mem[36] :
                        (N28)? mem[170] :
                        (N30)? mem[304] :
                        (N32)? mem[438] :
                        (N34)? mem[572] :
                        (N36)? mem[706] :
                        (N38)? mem[840] :
                        (N40)? mem[974] :
                        (N27)? mem[1108] :
                        (N29)? mem[1242] :
                        (N31)? mem[1376] :
                        (N33)? mem[1510] :
                        (N35)? mem[1644] :
                        (N37)? mem[1778] :
                        (N39)? mem[1912] :
                        (N41)? mem[2046] : 1'b0;
  assign r_data_o[35] = (N26)? mem[35] :
                        (N28)? mem[169] :
                        (N30)? mem[303] :
                        (N32)? mem[437] :
                        (N34)? mem[571] :
                        (N36)? mem[705] :
                        (N38)? mem[839] :
                        (N40)? mem[973] :
                        (N27)? mem[1107] :
                        (N29)? mem[1241] :
                        (N31)? mem[1375] :
                        (N33)? mem[1509] :
                        (N35)? mem[1643] :
                        (N37)? mem[1777] :
                        (N39)? mem[1911] :
                        (N41)? mem[2045] : 1'b0;
  assign r_data_o[34] = (N26)? mem[34] :
                        (N28)? mem[168] :
                        (N30)? mem[302] :
                        (N32)? mem[436] :
                        (N34)? mem[570] :
                        (N36)? mem[704] :
                        (N38)? mem[838] :
                        (N40)? mem[972] :
                        (N27)? mem[1106] :
                        (N29)? mem[1240] :
                        (N31)? mem[1374] :
                        (N33)? mem[1508] :
                        (N35)? mem[1642] :
                        (N37)? mem[1776] :
                        (N39)? mem[1910] :
                        (N41)? mem[2044] : 1'b0;
  assign r_data_o[33] = (N26)? mem[33] :
                        (N28)? mem[167] :
                        (N30)? mem[301] :
                        (N32)? mem[435] :
                        (N34)? mem[569] :
                        (N36)? mem[703] :
                        (N38)? mem[837] :
                        (N40)? mem[971] :
                        (N27)? mem[1105] :
                        (N29)? mem[1239] :
                        (N31)? mem[1373] :
                        (N33)? mem[1507] :
                        (N35)? mem[1641] :
                        (N37)? mem[1775] :
                        (N39)? mem[1909] :
                        (N41)? mem[2043] : 1'b0;
  assign r_data_o[32] = (N26)? mem[32] :
                        (N28)? mem[166] :
                        (N30)? mem[300] :
                        (N32)? mem[434] :
                        (N34)? mem[568] :
                        (N36)? mem[702] :
                        (N38)? mem[836] :
                        (N40)? mem[970] :
                        (N27)? mem[1104] :
                        (N29)? mem[1238] :
                        (N31)? mem[1372] :
                        (N33)? mem[1506] :
                        (N35)? mem[1640] :
                        (N37)? mem[1774] :
                        (N39)? mem[1908] :
                        (N41)? mem[2042] : 1'b0;
  assign r_data_o[31] = (N26)? mem[31] :
                        (N28)? mem[165] :
                        (N30)? mem[299] :
                        (N32)? mem[433] :
                        (N34)? mem[567] :
                        (N36)? mem[701] :
                        (N38)? mem[835] :
                        (N40)? mem[969] :
                        (N27)? mem[1103] :
                        (N29)? mem[1237] :
                        (N31)? mem[1371] :
                        (N33)? mem[1505] :
                        (N35)? mem[1639] :
                        (N37)? mem[1773] :
                        (N39)? mem[1907] :
                        (N41)? mem[2041] : 1'b0;
  assign r_data_o[30] = (N26)? mem[30] :
                        (N28)? mem[164] :
                        (N30)? mem[298] :
                        (N32)? mem[432] :
                        (N34)? mem[566] :
                        (N36)? mem[700] :
                        (N38)? mem[834] :
                        (N40)? mem[968] :
                        (N27)? mem[1102] :
                        (N29)? mem[1236] :
                        (N31)? mem[1370] :
                        (N33)? mem[1504] :
                        (N35)? mem[1638] :
                        (N37)? mem[1772] :
                        (N39)? mem[1906] :
                        (N41)? mem[2040] : 1'b0;
  assign r_data_o[29] = (N26)? mem[29] :
                        (N28)? mem[163] :
                        (N30)? mem[297] :
                        (N32)? mem[431] :
                        (N34)? mem[565] :
                        (N36)? mem[699] :
                        (N38)? mem[833] :
                        (N40)? mem[967] :
                        (N27)? mem[1101] :
                        (N29)? mem[1235] :
                        (N31)? mem[1369] :
                        (N33)? mem[1503] :
                        (N35)? mem[1637] :
                        (N37)? mem[1771] :
                        (N39)? mem[1905] :
                        (N41)? mem[2039] : 1'b0;
  assign r_data_o[28] = (N26)? mem[28] :
                        (N28)? mem[162] :
                        (N30)? mem[296] :
                        (N32)? mem[430] :
                        (N34)? mem[564] :
                        (N36)? mem[698] :
                        (N38)? mem[832] :
                        (N40)? mem[966] :
                        (N27)? mem[1100] :
                        (N29)? mem[1234] :
                        (N31)? mem[1368] :
                        (N33)? mem[1502] :
                        (N35)? mem[1636] :
                        (N37)? mem[1770] :
                        (N39)? mem[1904] :
                        (N41)? mem[2038] : 1'b0;
  assign r_data_o[27] = (N26)? mem[27] :
                        (N28)? mem[161] :
                        (N30)? mem[295] :
                        (N32)? mem[429] :
                        (N34)? mem[563] :
                        (N36)? mem[697] :
                        (N38)? mem[831] :
                        (N40)? mem[965] :
                        (N27)? mem[1099] :
                        (N29)? mem[1233] :
                        (N31)? mem[1367] :
                        (N33)? mem[1501] :
                        (N35)? mem[1635] :
                        (N37)? mem[1769] :
                        (N39)? mem[1903] :
                        (N41)? mem[2037] : 1'b0;
  assign r_data_o[26] = (N26)? mem[26] :
                        (N28)? mem[160] :
                        (N30)? mem[294] :
                        (N32)? mem[428] :
                        (N34)? mem[562] :
                        (N36)? mem[696] :
                        (N38)? mem[830] :
                        (N40)? mem[964] :
                        (N27)? mem[1098] :
                        (N29)? mem[1232] :
                        (N31)? mem[1366] :
                        (N33)? mem[1500] :
                        (N35)? mem[1634] :
                        (N37)? mem[1768] :
                        (N39)? mem[1902] :
                        (N41)? mem[2036] : 1'b0;
  assign r_data_o[25] = (N26)? mem[25] :
                        (N28)? mem[159] :
                        (N30)? mem[293] :
                        (N32)? mem[427] :
                        (N34)? mem[561] :
                        (N36)? mem[695] :
                        (N38)? mem[829] :
                        (N40)? mem[963] :
                        (N27)? mem[1097] :
                        (N29)? mem[1231] :
                        (N31)? mem[1365] :
                        (N33)? mem[1499] :
                        (N35)? mem[1633] :
                        (N37)? mem[1767] :
                        (N39)? mem[1901] :
                        (N41)? mem[2035] : 1'b0;
  assign r_data_o[24] = (N26)? mem[24] :
                        (N28)? mem[158] :
                        (N30)? mem[292] :
                        (N32)? mem[426] :
                        (N34)? mem[560] :
                        (N36)? mem[694] :
                        (N38)? mem[828] :
                        (N40)? mem[962] :
                        (N27)? mem[1096] :
                        (N29)? mem[1230] :
                        (N31)? mem[1364] :
                        (N33)? mem[1498] :
                        (N35)? mem[1632] :
                        (N37)? mem[1766] :
                        (N39)? mem[1900] :
                        (N41)? mem[2034] : 1'b0;
  assign r_data_o[23] = (N26)? mem[23] :
                        (N28)? mem[157] :
                        (N30)? mem[291] :
                        (N32)? mem[425] :
                        (N34)? mem[559] :
                        (N36)? mem[693] :
                        (N38)? mem[827] :
                        (N40)? mem[961] :
                        (N27)? mem[1095] :
                        (N29)? mem[1229] :
                        (N31)? mem[1363] :
                        (N33)? mem[1497] :
                        (N35)? mem[1631] :
                        (N37)? mem[1765] :
                        (N39)? mem[1899] :
                        (N41)? mem[2033] : 1'b0;
  assign r_data_o[22] = (N26)? mem[22] :
                        (N28)? mem[156] :
                        (N30)? mem[290] :
                        (N32)? mem[424] :
                        (N34)? mem[558] :
                        (N36)? mem[692] :
                        (N38)? mem[826] :
                        (N40)? mem[960] :
                        (N27)? mem[1094] :
                        (N29)? mem[1228] :
                        (N31)? mem[1362] :
                        (N33)? mem[1496] :
                        (N35)? mem[1630] :
                        (N37)? mem[1764] :
                        (N39)? mem[1898] :
                        (N41)? mem[2032] : 1'b0;
  assign r_data_o[21] = (N26)? mem[21] :
                        (N28)? mem[155] :
                        (N30)? mem[289] :
                        (N32)? mem[423] :
                        (N34)? mem[557] :
                        (N36)? mem[691] :
                        (N38)? mem[825] :
                        (N40)? mem[959] :
                        (N27)? mem[1093] :
                        (N29)? mem[1227] :
                        (N31)? mem[1361] :
                        (N33)? mem[1495] :
                        (N35)? mem[1629] :
                        (N37)? mem[1763] :
                        (N39)? mem[1897] :
                        (N41)? mem[2031] : 1'b0;
  assign r_data_o[20] = (N26)? mem[20] :
                        (N28)? mem[154] :
                        (N30)? mem[288] :
                        (N32)? mem[422] :
                        (N34)? mem[556] :
                        (N36)? mem[690] :
                        (N38)? mem[824] :
                        (N40)? mem[958] :
                        (N27)? mem[1092] :
                        (N29)? mem[1226] :
                        (N31)? mem[1360] :
                        (N33)? mem[1494] :
                        (N35)? mem[1628] :
                        (N37)? mem[1762] :
                        (N39)? mem[1896] :
                        (N41)? mem[2030] : 1'b0;
  assign r_data_o[19] = (N26)? mem[19] :
                        (N28)? mem[153] :
                        (N30)? mem[287] :
                        (N32)? mem[421] :
                        (N34)? mem[555] :
                        (N36)? mem[689] :
                        (N38)? mem[823] :
                        (N40)? mem[957] :
                        (N27)? mem[1091] :
                        (N29)? mem[1225] :
                        (N31)? mem[1359] :
                        (N33)? mem[1493] :
                        (N35)? mem[1627] :
                        (N37)? mem[1761] :
                        (N39)? mem[1895] :
                        (N41)? mem[2029] : 1'b0;
  assign r_data_o[18] = (N26)? mem[18] :
                        (N28)? mem[152] :
                        (N30)? mem[286] :
                        (N32)? mem[420] :
                        (N34)? mem[554] :
                        (N36)? mem[688] :
                        (N38)? mem[822] :
                        (N40)? mem[956] :
                        (N27)? mem[1090] :
                        (N29)? mem[1224] :
                        (N31)? mem[1358] :
                        (N33)? mem[1492] :
                        (N35)? mem[1626] :
                        (N37)? mem[1760] :
                        (N39)? mem[1894] :
                        (N41)? mem[2028] : 1'b0;
  assign r_data_o[17] = (N26)? mem[17] :
                        (N28)? mem[151] :
                        (N30)? mem[285] :
                        (N32)? mem[419] :
                        (N34)? mem[553] :
                        (N36)? mem[687] :
                        (N38)? mem[821] :
                        (N40)? mem[955] :
                        (N27)? mem[1089] :
                        (N29)? mem[1223] :
                        (N31)? mem[1357] :
                        (N33)? mem[1491] :
                        (N35)? mem[1625] :
                        (N37)? mem[1759] :
                        (N39)? mem[1893] :
                        (N41)? mem[2027] : 1'b0;
  assign r_data_o[16] = (N26)? mem[16] :
                        (N28)? mem[150] :
                        (N30)? mem[284] :
                        (N32)? mem[418] :
                        (N34)? mem[552] :
                        (N36)? mem[686] :
                        (N38)? mem[820] :
                        (N40)? mem[954] :
                        (N27)? mem[1088] :
                        (N29)? mem[1222] :
                        (N31)? mem[1356] :
                        (N33)? mem[1490] :
                        (N35)? mem[1624] :
                        (N37)? mem[1758] :
                        (N39)? mem[1892] :
                        (N41)? mem[2026] : 1'b0;
  assign r_data_o[15] = (N26)? mem[15] :
                        (N28)? mem[149] :
                        (N30)? mem[283] :
                        (N32)? mem[417] :
                        (N34)? mem[551] :
                        (N36)? mem[685] :
                        (N38)? mem[819] :
                        (N40)? mem[953] :
                        (N27)? mem[1087] :
                        (N29)? mem[1221] :
                        (N31)? mem[1355] :
                        (N33)? mem[1489] :
                        (N35)? mem[1623] :
                        (N37)? mem[1757] :
                        (N39)? mem[1891] :
                        (N41)? mem[2025] : 1'b0;
  assign r_data_o[14] = (N26)? mem[14] :
                        (N28)? mem[148] :
                        (N30)? mem[282] :
                        (N32)? mem[416] :
                        (N34)? mem[550] :
                        (N36)? mem[684] :
                        (N38)? mem[818] :
                        (N40)? mem[952] :
                        (N27)? mem[1086] :
                        (N29)? mem[1220] :
                        (N31)? mem[1354] :
                        (N33)? mem[1488] :
                        (N35)? mem[1622] :
                        (N37)? mem[1756] :
                        (N39)? mem[1890] :
                        (N41)? mem[2024] : 1'b0;
  assign r_data_o[13] = (N26)? mem[13] :
                        (N28)? mem[147] :
                        (N30)? mem[281] :
                        (N32)? mem[415] :
                        (N34)? mem[549] :
                        (N36)? mem[683] :
                        (N38)? mem[817] :
                        (N40)? mem[951] :
                        (N27)? mem[1085] :
                        (N29)? mem[1219] :
                        (N31)? mem[1353] :
                        (N33)? mem[1487] :
                        (N35)? mem[1621] :
                        (N37)? mem[1755] :
                        (N39)? mem[1889] :
                        (N41)? mem[2023] : 1'b0;
  assign r_data_o[12] = (N26)? mem[12] :
                        (N28)? mem[146] :
                        (N30)? mem[280] :
                        (N32)? mem[414] :
                        (N34)? mem[548] :
                        (N36)? mem[682] :
                        (N38)? mem[816] :
                        (N40)? mem[950] :
                        (N27)? mem[1084] :
                        (N29)? mem[1218] :
                        (N31)? mem[1352] :
                        (N33)? mem[1486] :
                        (N35)? mem[1620] :
                        (N37)? mem[1754] :
                        (N39)? mem[1888] :
                        (N41)? mem[2022] : 1'b0;
  assign r_data_o[11] = (N26)? mem[11] :
                        (N28)? mem[145] :
                        (N30)? mem[279] :
                        (N32)? mem[413] :
                        (N34)? mem[547] :
                        (N36)? mem[681] :
                        (N38)? mem[815] :
                        (N40)? mem[949] :
                        (N27)? mem[1083] :
                        (N29)? mem[1217] :
                        (N31)? mem[1351] :
                        (N33)? mem[1485] :
                        (N35)? mem[1619] :
                        (N37)? mem[1753] :
                        (N39)? mem[1887] :
                        (N41)? mem[2021] : 1'b0;
  assign r_data_o[10] = (N26)? mem[10] :
                        (N28)? mem[144] :
                        (N30)? mem[278] :
                        (N32)? mem[412] :
                        (N34)? mem[546] :
                        (N36)? mem[680] :
                        (N38)? mem[814] :
                        (N40)? mem[948] :
                        (N27)? mem[1082] :
                        (N29)? mem[1216] :
                        (N31)? mem[1350] :
                        (N33)? mem[1484] :
                        (N35)? mem[1618] :
                        (N37)? mem[1752] :
                        (N39)? mem[1886] :
                        (N41)? mem[2020] : 1'b0;
  assign r_data_o[9] = (N26)? mem[9] :
                       (N28)? mem[143] :
                       (N30)? mem[277] :
                       (N32)? mem[411] :
                       (N34)? mem[545] :
                       (N36)? mem[679] :
                       (N38)? mem[813] :
                       (N40)? mem[947] :
                       (N27)? mem[1081] :
                       (N29)? mem[1215] :
                       (N31)? mem[1349] :
                       (N33)? mem[1483] :
                       (N35)? mem[1617] :
                       (N37)? mem[1751] :
                       (N39)? mem[1885] :
                       (N41)? mem[2019] : 1'b0;
  assign r_data_o[8] = (N26)? mem[8] :
                       (N28)? mem[142] :
                       (N30)? mem[276] :
                       (N32)? mem[410] :
                       (N34)? mem[544] :
                       (N36)? mem[678] :
                       (N38)? mem[812] :
                       (N40)? mem[946] :
                       (N27)? mem[1080] :
                       (N29)? mem[1214] :
                       (N31)? mem[1348] :
                       (N33)? mem[1482] :
                       (N35)? mem[1616] :
                       (N37)? mem[1750] :
                       (N39)? mem[1884] :
                       (N41)? mem[2018] : 1'b0;
  assign r_data_o[7] = (N26)? mem[7] :
                       (N28)? mem[141] :
                       (N30)? mem[275] :
                       (N32)? mem[409] :
                       (N34)? mem[543] :
                       (N36)? mem[677] :
                       (N38)? mem[811] :
                       (N40)? mem[945] :
                       (N27)? mem[1079] :
                       (N29)? mem[1213] :
                       (N31)? mem[1347] :
                       (N33)? mem[1481] :
                       (N35)? mem[1615] :
                       (N37)? mem[1749] :
                       (N39)? mem[1883] :
                       (N41)? mem[2017] : 1'b0;
  assign r_data_o[6] = (N26)? mem[6] :
                       (N28)? mem[140] :
                       (N30)? mem[274] :
                       (N32)? mem[408] :
                       (N34)? mem[542] :
                       (N36)? mem[676] :
                       (N38)? mem[810] :
                       (N40)? mem[944] :
                       (N27)? mem[1078] :
                       (N29)? mem[1212] :
                       (N31)? mem[1346] :
                       (N33)? mem[1480] :
                       (N35)? mem[1614] :
                       (N37)? mem[1748] :
                       (N39)? mem[1882] :
                       (N41)? mem[2016] : 1'b0;
  assign r_data_o[5] = (N26)? mem[5] :
                       (N28)? mem[139] :
                       (N30)? mem[273] :
                       (N32)? mem[407] :
                       (N34)? mem[541] :
                       (N36)? mem[675] :
                       (N38)? mem[809] :
                       (N40)? mem[943] :
                       (N27)? mem[1077] :
                       (N29)? mem[1211] :
                       (N31)? mem[1345] :
                       (N33)? mem[1479] :
                       (N35)? mem[1613] :
                       (N37)? mem[1747] :
                       (N39)? mem[1881] :
                       (N41)? mem[2015] : 1'b0;
  assign r_data_o[4] = (N26)? mem[4] :
                       (N28)? mem[138] :
                       (N30)? mem[272] :
                       (N32)? mem[406] :
                       (N34)? mem[540] :
                       (N36)? mem[674] :
                       (N38)? mem[808] :
                       (N40)? mem[942] :
                       (N27)? mem[1076] :
                       (N29)? mem[1210] :
                       (N31)? mem[1344] :
                       (N33)? mem[1478] :
                       (N35)? mem[1612] :
                       (N37)? mem[1746] :
                       (N39)? mem[1880] :
                       (N41)? mem[2014] : 1'b0;
  assign r_data_o[3] = (N26)? mem[3] :
                       (N28)? mem[137] :
                       (N30)? mem[271] :
                       (N32)? mem[405] :
                       (N34)? mem[539] :
                       (N36)? mem[673] :
                       (N38)? mem[807] :
                       (N40)? mem[941] :
                       (N27)? mem[1075] :
                       (N29)? mem[1209] :
                       (N31)? mem[1343] :
                       (N33)? mem[1477] :
                       (N35)? mem[1611] :
                       (N37)? mem[1745] :
                       (N39)? mem[1879] :
                       (N41)? mem[2013] : 1'b0;
  assign r_data_o[2] = (N26)? mem[2] :
                       (N28)? mem[136] :
                       (N30)? mem[270] :
                       (N32)? mem[404] :
                       (N34)? mem[538] :
                       (N36)? mem[672] :
                       (N38)? mem[806] :
                       (N40)? mem[940] :
                       (N27)? mem[1074] :
                       (N29)? mem[1208] :
                       (N31)? mem[1342] :
                       (N33)? mem[1476] :
                       (N35)? mem[1610] :
                       (N37)? mem[1744] :
                       (N39)? mem[1878] :
                       (N41)? mem[2012] : 1'b0;
  assign r_data_o[1] = (N26)? mem[1] :
                       (N28)? mem[135] :
                       (N30)? mem[269] :
                       (N32)? mem[403] :
                       (N34)? mem[537] :
                       (N36)? mem[671] :
                       (N38)? mem[805] :
                       (N40)? mem[939] :
                       (N27)? mem[1073] :
                       (N29)? mem[1207] :
                       (N31)? mem[1341] :
                       (N33)? mem[1475] :
                       (N35)? mem[1609] :
                       (N37)? mem[1743] :
                       (N39)? mem[1877] :
                       (N41)? mem[2011] : 1'b0;
  assign r_data_o[0] = (N26)? mem[0] :
                       (N28)? mem[134] :
                       (N30)? mem[268] :
                       (N32)? mem[402] :
                       (N34)? mem[536] :
                       (N36)? mem[670] :
                       (N38)? mem[804] :
                       (N40)? mem[938] :
                       (N27)? mem[1072] :
                       (N29)? mem[1206] :
                       (N31)? mem[1340] :
                       (N33)? mem[1474] :
                       (N35)? mem[1608] :
                       (N37)? mem[1742] :
                       (N39)? mem[1876] :
                       (N41)? mem[2010] : 1'b0;
  assign N91 = w_addr_i[2] & w_addr_i[3];
  assign N92 = N0 & w_addr_i[3];
  assign N0 = ~w_addr_i[2];
  assign N93 = w_addr_i[2] & N1;
  assign N1 = ~w_addr_i[3];
  assign N94 = N2 & N3;
  assign N2 = ~w_addr_i[2];
  assign N3 = ~w_addr_i[3];
  assign N95 = w_addr_i[0] & w_addr_i[1];
  assign N96 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N97 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N98 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N58 = N91 & N95;
  assign N57 = N91 & N96;
  assign N56 = N91 & N97;
  assign N55 = N91 & N98;
  assign N54 = N92 & N95;
  assign N53 = N92 & N96;
  assign N52 = N92 & N97;
  assign N51 = N92 & N98;
  assign N50 = N93 & N95;
  assign N49 = N93 & N96;
  assign N48 = N93 & N97;
  assign N47 = N93 & N98;
  assign N46 = N94 & N95;
  assign N45 = N94 & N96;
  assign N44 = N94 & N97;
  assign N43 = N94 & N98;
  assign { N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59 } = (N8)? { N58, N58, N57, N57, N56, N56, N55, N55, N54, N54, N53, N53, N52, N52, N51, N51, N50, N50, N49, N49, N48, N48, N47, N47, N46, N46, N45, N45, N44, N44, N43, N43 } :
                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N42;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~r_addr_i[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_i[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_i[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_i[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_i[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N89) begin
      { mem[2143:2045], mem[2010:2010] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N90) begin
      { mem[2044:2011] } <= { w_data_i[34:1] };
    end
    if(N87) begin
      { mem[2009:1911], mem[1876:1876] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N88) begin
      { mem[1910:1877] } <= { w_data_i[34:1] };
    end
    if(N85) begin
      { mem[1875:1777], mem[1742:1742] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N86) begin
      { mem[1776:1743] } <= { w_data_i[34:1] };
    end
    if(N83) begin
      { mem[1741:1643], mem[1608:1608] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N84) begin
      { mem[1642:1609] } <= { w_data_i[34:1] };
    end
    if(N81) begin
      { mem[1607:1509], mem[1474:1474] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N82) begin
      { mem[1508:1475] } <= { w_data_i[34:1] };
    end
    if(N79) begin
      { mem[1473:1375], mem[1340:1340] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N80) begin
      { mem[1374:1341] } <= { w_data_i[34:1] };
    end
    if(N77) begin
      { mem[1339:1241], mem[1206:1206] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N78) begin
      { mem[1240:1207] } <= { w_data_i[34:1] };
    end
    if(N75) begin
      { mem[1205:1107], mem[1072:1072] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N76) begin
      { mem[1106:1073] } <= { w_data_i[34:1] };
    end
    if(N73) begin
      { mem[1071:973], mem[938:938] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N74) begin
      { mem[972:939] } <= { w_data_i[34:1] };
    end
    if(N71) begin
      { mem[937:839], mem[804:804] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N72) begin
      { mem[838:805] } <= { w_data_i[34:1] };
    end
    if(N69) begin
      { mem[803:705], mem[670:670] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N70) begin
      { mem[704:671] } <= { w_data_i[34:1] };
    end
    if(N67) begin
      { mem[669:571], mem[536:536] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N68) begin
      { mem[570:537] } <= { w_data_i[34:1] };
    end
    if(N65) begin
      { mem[535:437], mem[402:402] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N66) begin
      { mem[436:403] } <= { w_data_i[34:1] };
    end
    if(N63) begin
      { mem[401:303], mem[268:268] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N64) begin
      { mem[302:269] } <= { w_data_i[34:1] };
    end
    if(N61) begin
      { mem[267:169], mem[134:134] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N62) begin
      { mem[168:135] } <= { w_data_i[34:1] };
    end
    if(N59) begin
      { mem[133:35], mem[0:0] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N60) begin
      { mem[34:1] } <= { w_data_i[34:1] };
    end
  end


endmodule