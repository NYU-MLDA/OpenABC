module bsg_mem_1rw_sync_mask_write_bit_synth_width_p15_els_p128
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [14:0] data_i;
  input [6:0] addr_i;
  input [14:0] w_mask_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [14:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,
  N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,
  N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,
  N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,
  N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,
  N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,
  N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,
  N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,
  N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,
  N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,
  N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
  N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
  N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,
  N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,
  N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,
  N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,
  N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,
  N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,
  N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,
  N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,
  N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,
  N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,
  N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,
  N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,
  N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,
  N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,
  N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,
  N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,
  N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,
  N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,
  N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,
  N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,
  N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,
  N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,
  N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,
  N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,
  N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,
  N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,
  N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,
  N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,
  N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,
  N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,
  N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,
  N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,
  N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,
  N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,
  N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,
  N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,
  N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,
  N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,
  N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,
  N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,
  N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,
  N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,
  N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,
  N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,
  N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,
  N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,
  N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,
  N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,
  N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,
  N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,
  N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,
  N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,
  N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,
  N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,
  N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,
  N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,
  N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104,
  N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,
  N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,N4130,
  N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,N4143,N4144,
  N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,
  N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,N4170,
  N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,N4183,N4184,
  N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
  N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,N4210,
  N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,N4223,N4224,
  N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,
  N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,N4250,
  N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,N4263,N4264,
  N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,
  N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,N4290,
  N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,N4303,N4304,
  N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,
  N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,N4330,
  N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,N4343,N4344,
  N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,
  N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,N4370,
  N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,N4383,N4384,
  N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,
  N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,N4410,
  N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,N4423,N4424,
  N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,
  N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,N4450,
  N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,N4463,N4464,
  N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
  N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,
  N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,
  N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
  N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,
  N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,
  N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,
  N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,N4570,
  N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,N4583,N4584,
  N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,
  N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4610,
  N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,
  N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,
  N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,
  N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,N4663,N4664,
  N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,
  N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,N4690,
  N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4703,N4704,
  N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,
  N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,N4730,
  N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,N4743,N4744,
  N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,
  N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4770,
  N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
  N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,
  N4798,N4799,N4800,N4801,N4802,N4803,N4804;
  wire [6:0] addr_r;
  wire [1919:0] mem;
  reg addr_r_6_sv2v_reg,addr_r_5_sv2v_reg,addr_r_4_sv2v_reg,addr_r_3_sv2v_reg,
  addr_r_2_sv2v_reg,addr_r_1_sv2v_reg,addr_r_0_sv2v_reg,mem_1919_sv2v_reg,
  mem_1918_sv2v_reg,mem_1917_sv2v_reg,mem_1916_sv2v_reg,mem_1915_sv2v_reg,mem_1914_sv2v_reg,
  mem_1913_sv2v_reg,mem_1912_sv2v_reg,mem_1911_sv2v_reg,mem_1910_sv2v_reg,
  mem_1909_sv2v_reg,mem_1908_sv2v_reg,mem_1907_sv2v_reg,mem_1906_sv2v_reg,mem_1905_sv2v_reg,
  mem_1904_sv2v_reg,mem_1903_sv2v_reg,mem_1902_sv2v_reg,mem_1901_sv2v_reg,
  mem_1900_sv2v_reg,mem_1899_sv2v_reg,mem_1898_sv2v_reg,mem_1897_sv2v_reg,mem_1896_sv2v_reg,
  mem_1895_sv2v_reg,mem_1894_sv2v_reg,mem_1893_sv2v_reg,mem_1892_sv2v_reg,
  mem_1891_sv2v_reg,mem_1890_sv2v_reg,mem_1889_sv2v_reg,mem_1888_sv2v_reg,mem_1887_sv2v_reg,
  mem_1886_sv2v_reg,mem_1885_sv2v_reg,mem_1884_sv2v_reg,mem_1883_sv2v_reg,
  mem_1882_sv2v_reg,mem_1881_sv2v_reg,mem_1880_sv2v_reg,mem_1879_sv2v_reg,
  mem_1878_sv2v_reg,mem_1877_sv2v_reg,mem_1876_sv2v_reg,mem_1875_sv2v_reg,mem_1874_sv2v_reg,
  mem_1873_sv2v_reg,mem_1872_sv2v_reg,mem_1871_sv2v_reg,mem_1870_sv2v_reg,
  mem_1869_sv2v_reg,mem_1868_sv2v_reg,mem_1867_sv2v_reg,mem_1866_sv2v_reg,mem_1865_sv2v_reg,
  mem_1864_sv2v_reg,mem_1863_sv2v_reg,mem_1862_sv2v_reg,mem_1861_sv2v_reg,
  mem_1860_sv2v_reg,mem_1859_sv2v_reg,mem_1858_sv2v_reg,mem_1857_sv2v_reg,mem_1856_sv2v_reg,
  mem_1855_sv2v_reg,mem_1854_sv2v_reg,mem_1853_sv2v_reg,mem_1852_sv2v_reg,
  mem_1851_sv2v_reg,mem_1850_sv2v_reg,mem_1849_sv2v_reg,mem_1848_sv2v_reg,mem_1847_sv2v_reg,
  mem_1846_sv2v_reg,mem_1845_sv2v_reg,mem_1844_sv2v_reg,mem_1843_sv2v_reg,
  mem_1842_sv2v_reg,mem_1841_sv2v_reg,mem_1840_sv2v_reg,mem_1839_sv2v_reg,
  mem_1838_sv2v_reg,mem_1837_sv2v_reg,mem_1836_sv2v_reg,mem_1835_sv2v_reg,mem_1834_sv2v_reg,
  mem_1833_sv2v_reg,mem_1832_sv2v_reg,mem_1831_sv2v_reg,mem_1830_sv2v_reg,
  mem_1829_sv2v_reg,mem_1828_sv2v_reg,mem_1827_sv2v_reg,mem_1826_sv2v_reg,mem_1825_sv2v_reg,
  mem_1824_sv2v_reg,mem_1823_sv2v_reg,mem_1822_sv2v_reg,mem_1821_sv2v_reg,
  mem_1820_sv2v_reg,mem_1819_sv2v_reg,mem_1818_sv2v_reg,mem_1817_sv2v_reg,mem_1816_sv2v_reg,
  mem_1815_sv2v_reg,mem_1814_sv2v_reg,mem_1813_sv2v_reg,mem_1812_sv2v_reg,
  mem_1811_sv2v_reg,mem_1810_sv2v_reg,mem_1809_sv2v_reg,mem_1808_sv2v_reg,mem_1807_sv2v_reg,
  mem_1806_sv2v_reg,mem_1805_sv2v_reg,mem_1804_sv2v_reg,mem_1803_sv2v_reg,
  mem_1802_sv2v_reg,mem_1801_sv2v_reg,mem_1800_sv2v_reg,mem_1799_sv2v_reg,
  mem_1798_sv2v_reg,mem_1797_sv2v_reg,mem_1796_sv2v_reg,mem_1795_sv2v_reg,mem_1794_sv2v_reg,
  mem_1793_sv2v_reg,mem_1792_sv2v_reg,mem_1791_sv2v_reg,mem_1790_sv2v_reg,
  mem_1789_sv2v_reg,mem_1788_sv2v_reg,mem_1787_sv2v_reg,mem_1786_sv2v_reg,mem_1785_sv2v_reg,
  mem_1784_sv2v_reg,mem_1783_sv2v_reg,mem_1782_sv2v_reg,mem_1781_sv2v_reg,
  mem_1780_sv2v_reg,mem_1779_sv2v_reg,mem_1778_sv2v_reg,mem_1777_sv2v_reg,mem_1776_sv2v_reg,
  mem_1775_sv2v_reg,mem_1774_sv2v_reg,mem_1773_sv2v_reg,mem_1772_sv2v_reg,
  mem_1771_sv2v_reg,mem_1770_sv2v_reg,mem_1769_sv2v_reg,mem_1768_sv2v_reg,mem_1767_sv2v_reg,
  mem_1766_sv2v_reg,mem_1765_sv2v_reg,mem_1764_sv2v_reg,mem_1763_sv2v_reg,
  mem_1762_sv2v_reg,mem_1761_sv2v_reg,mem_1760_sv2v_reg,mem_1759_sv2v_reg,
  mem_1758_sv2v_reg,mem_1757_sv2v_reg,mem_1756_sv2v_reg,mem_1755_sv2v_reg,mem_1754_sv2v_reg,
  mem_1753_sv2v_reg,mem_1752_sv2v_reg,mem_1751_sv2v_reg,mem_1750_sv2v_reg,
  mem_1749_sv2v_reg,mem_1748_sv2v_reg,mem_1747_sv2v_reg,mem_1746_sv2v_reg,mem_1745_sv2v_reg,
  mem_1744_sv2v_reg,mem_1743_sv2v_reg,mem_1742_sv2v_reg,mem_1741_sv2v_reg,
  mem_1740_sv2v_reg,mem_1739_sv2v_reg,mem_1738_sv2v_reg,mem_1737_sv2v_reg,mem_1736_sv2v_reg,
  mem_1735_sv2v_reg,mem_1734_sv2v_reg,mem_1733_sv2v_reg,mem_1732_sv2v_reg,
  mem_1731_sv2v_reg,mem_1730_sv2v_reg,mem_1729_sv2v_reg,mem_1728_sv2v_reg,mem_1727_sv2v_reg,
  mem_1726_sv2v_reg,mem_1725_sv2v_reg,mem_1724_sv2v_reg,mem_1723_sv2v_reg,
  mem_1722_sv2v_reg,mem_1721_sv2v_reg,mem_1720_sv2v_reg,mem_1719_sv2v_reg,
  mem_1718_sv2v_reg,mem_1717_sv2v_reg,mem_1716_sv2v_reg,mem_1715_sv2v_reg,mem_1714_sv2v_reg,
  mem_1713_sv2v_reg,mem_1712_sv2v_reg,mem_1711_sv2v_reg,mem_1710_sv2v_reg,
  mem_1709_sv2v_reg,mem_1708_sv2v_reg,mem_1707_sv2v_reg,mem_1706_sv2v_reg,mem_1705_sv2v_reg,
  mem_1704_sv2v_reg,mem_1703_sv2v_reg,mem_1702_sv2v_reg,mem_1701_sv2v_reg,
  mem_1700_sv2v_reg,mem_1699_sv2v_reg,mem_1698_sv2v_reg,mem_1697_sv2v_reg,mem_1696_sv2v_reg,
  mem_1695_sv2v_reg,mem_1694_sv2v_reg,mem_1693_sv2v_reg,mem_1692_sv2v_reg,
  mem_1691_sv2v_reg,mem_1690_sv2v_reg,mem_1689_sv2v_reg,mem_1688_sv2v_reg,mem_1687_sv2v_reg,
  mem_1686_sv2v_reg,mem_1685_sv2v_reg,mem_1684_sv2v_reg,mem_1683_sv2v_reg,
  mem_1682_sv2v_reg,mem_1681_sv2v_reg,mem_1680_sv2v_reg,mem_1679_sv2v_reg,
  mem_1678_sv2v_reg,mem_1677_sv2v_reg,mem_1676_sv2v_reg,mem_1675_sv2v_reg,mem_1674_sv2v_reg,
  mem_1673_sv2v_reg,mem_1672_sv2v_reg,mem_1671_sv2v_reg,mem_1670_sv2v_reg,
  mem_1669_sv2v_reg,mem_1668_sv2v_reg,mem_1667_sv2v_reg,mem_1666_sv2v_reg,mem_1665_sv2v_reg,
  mem_1664_sv2v_reg,mem_1663_sv2v_reg,mem_1662_sv2v_reg,mem_1661_sv2v_reg,
  mem_1660_sv2v_reg,mem_1659_sv2v_reg,mem_1658_sv2v_reg,mem_1657_sv2v_reg,mem_1656_sv2v_reg,
  mem_1655_sv2v_reg,mem_1654_sv2v_reg,mem_1653_sv2v_reg,mem_1652_sv2v_reg,
  mem_1651_sv2v_reg,mem_1650_sv2v_reg,mem_1649_sv2v_reg,mem_1648_sv2v_reg,mem_1647_sv2v_reg,
  mem_1646_sv2v_reg,mem_1645_sv2v_reg,mem_1644_sv2v_reg,mem_1643_sv2v_reg,
  mem_1642_sv2v_reg,mem_1641_sv2v_reg,mem_1640_sv2v_reg,mem_1639_sv2v_reg,
  mem_1638_sv2v_reg,mem_1637_sv2v_reg,mem_1636_sv2v_reg,mem_1635_sv2v_reg,mem_1634_sv2v_reg,
  mem_1633_sv2v_reg,mem_1632_sv2v_reg,mem_1631_sv2v_reg,mem_1630_sv2v_reg,
  mem_1629_sv2v_reg,mem_1628_sv2v_reg,mem_1627_sv2v_reg,mem_1626_sv2v_reg,mem_1625_sv2v_reg,
  mem_1624_sv2v_reg,mem_1623_sv2v_reg,mem_1622_sv2v_reg,mem_1621_sv2v_reg,
  mem_1620_sv2v_reg,mem_1619_sv2v_reg,mem_1618_sv2v_reg,mem_1617_sv2v_reg,mem_1616_sv2v_reg,
  mem_1615_sv2v_reg,mem_1614_sv2v_reg,mem_1613_sv2v_reg,mem_1612_sv2v_reg,
  mem_1611_sv2v_reg,mem_1610_sv2v_reg,mem_1609_sv2v_reg,mem_1608_sv2v_reg,mem_1607_sv2v_reg,
  mem_1606_sv2v_reg,mem_1605_sv2v_reg,mem_1604_sv2v_reg,mem_1603_sv2v_reg,
  mem_1602_sv2v_reg,mem_1601_sv2v_reg,mem_1600_sv2v_reg,mem_1599_sv2v_reg,
  mem_1598_sv2v_reg,mem_1597_sv2v_reg,mem_1596_sv2v_reg,mem_1595_sv2v_reg,mem_1594_sv2v_reg,
  mem_1593_sv2v_reg,mem_1592_sv2v_reg,mem_1591_sv2v_reg,mem_1590_sv2v_reg,
  mem_1589_sv2v_reg,mem_1588_sv2v_reg,mem_1587_sv2v_reg,mem_1586_sv2v_reg,mem_1585_sv2v_reg,
  mem_1584_sv2v_reg,mem_1583_sv2v_reg,mem_1582_sv2v_reg,mem_1581_sv2v_reg,
  mem_1580_sv2v_reg,mem_1579_sv2v_reg,mem_1578_sv2v_reg,mem_1577_sv2v_reg,mem_1576_sv2v_reg,
  mem_1575_sv2v_reg,mem_1574_sv2v_reg,mem_1573_sv2v_reg,mem_1572_sv2v_reg,
  mem_1571_sv2v_reg,mem_1570_sv2v_reg,mem_1569_sv2v_reg,mem_1568_sv2v_reg,mem_1567_sv2v_reg,
  mem_1566_sv2v_reg,mem_1565_sv2v_reg,mem_1564_sv2v_reg,mem_1563_sv2v_reg,
  mem_1562_sv2v_reg,mem_1561_sv2v_reg,mem_1560_sv2v_reg,mem_1559_sv2v_reg,
  mem_1558_sv2v_reg,mem_1557_sv2v_reg,mem_1556_sv2v_reg,mem_1555_sv2v_reg,mem_1554_sv2v_reg,
  mem_1553_sv2v_reg,mem_1552_sv2v_reg,mem_1551_sv2v_reg,mem_1550_sv2v_reg,
  mem_1549_sv2v_reg,mem_1548_sv2v_reg,mem_1547_sv2v_reg,mem_1546_sv2v_reg,mem_1545_sv2v_reg,
  mem_1544_sv2v_reg,mem_1543_sv2v_reg,mem_1542_sv2v_reg,mem_1541_sv2v_reg,
  mem_1540_sv2v_reg,mem_1539_sv2v_reg,mem_1538_sv2v_reg,mem_1537_sv2v_reg,mem_1536_sv2v_reg,
  mem_1535_sv2v_reg,mem_1534_sv2v_reg,mem_1533_sv2v_reg,mem_1532_sv2v_reg,
  mem_1531_sv2v_reg,mem_1530_sv2v_reg,mem_1529_sv2v_reg,mem_1528_sv2v_reg,mem_1527_sv2v_reg,
  mem_1526_sv2v_reg,mem_1525_sv2v_reg,mem_1524_sv2v_reg,mem_1523_sv2v_reg,
  mem_1522_sv2v_reg,mem_1521_sv2v_reg,mem_1520_sv2v_reg,mem_1519_sv2v_reg,
  mem_1518_sv2v_reg,mem_1517_sv2v_reg,mem_1516_sv2v_reg,mem_1515_sv2v_reg,mem_1514_sv2v_reg,
  mem_1513_sv2v_reg,mem_1512_sv2v_reg,mem_1511_sv2v_reg,mem_1510_sv2v_reg,
  mem_1509_sv2v_reg,mem_1508_sv2v_reg,mem_1507_sv2v_reg,mem_1506_sv2v_reg,mem_1505_sv2v_reg,
  mem_1504_sv2v_reg,mem_1503_sv2v_reg,mem_1502_sv2v_reg,mem_1501_sv2v_reg,
  mem_1500_sv2v_reg,mem_1499_sv2v_reg,mem_1498_sv2v_reg,mem_1497_sv2v_reg,mem_1496_sv2v_reg,
  mem_1495_sv2v_reg,mem_1494_sv2v_reg,mem_1493_sv2v_reg,mem_1492_sv2v_reg,
  mem_1491_sv2v_reg,mem_1490_sv2v_reg,mem_1489_sv2v_reg,mem_1488_sv2v_reg,mem_1487_sv2v_reg,
  mem_1486_sv2v_reg,mem_1485_sv2v_reg,mem_1484_sv2v_reg,mem_1483_sv2v_reg,
  mem_1482_sv2v_reg,mem_1481_sv2v_reg,mem_1480_sv2v_reg,mem_1479_sv2v_reg,
  mem_1478_sv2v_reg,mem_1477_sv2v_reg,mem_1476_sv2v_reg,mem_1475_sv2v_reg,mem_1474_sv2v_reg,
  mem_1473_sv2v_reg,mem_1472_sv2v_reg,mem_1471_sv2v_reg,mem_1470_sv2v_reg,
  mem_1469_sv2v_reg,mem_1468_sv2v_reg,mem_1467_sv2v_reg,mem_1466_sv2v_reg,mem_1465_sv2v_reg,
  mem_1464_sv2v_reg,mem_1463_sv2v_reg,mem_1462_sv2v_reg,mem_1461_sv2v_reg,
  mem_1460_sv2v_reg,mem_1459_sv2v_reg,mem_1458_sv2v_reg,mem_1457_sv2v_reg,mem_1456_sv2v_reg,
  mem_1455_sv2v_reg,mem_1454_sv2v_reg,mem_1453_sv2v_reg,mem_1452_sv2v_reg,
  mem_1451_sv2v_reg,mem_1450_sv2v_reg,mem_1449_sv2v_reg,mem_1448_sv2v_reg,mem_1447_sv2v_reg,
  mem_1446_sv2v_reg,mem_1445_sv2v_reg,mem_1444_sv2v_reg,mem_1443_sv2v_reg,
  mem_1442_sv2v_reg,mem_1441_sv2v_reg,mem_1440_sv2v_reg,mem_1439_sv2v_reg,
  mem_1438_sv2v_reg,mem_1437_sv2v_reg,mem_1436_sv2v_reg,mem_1435_sv2v_reg,mem_1434_sv2v_reg,
  mem_1433_sv2v_reg,mem_1432_sv2v_reg,mem_1431_sv2v_reg,mem_1430_sv2v_reg,
  mem_1429_sv2v_reg,mem_1428_sv2v_reg,mem_1427_sv2v_reg,mem_1426_sv2v_reg,mem_1425_sv2v_reg,
  mem_1424_sv2v_reg,mem_1423_sv2v_reg,mem_1422_sv2v_reg,mem_1421_sv2v_reg,
  mem_1420_sv2v_reg,mem_1419_sv2v_reg,mem_1418_sv2v_reg,mem_1417_sv2v_reg,mem_1416_sv2v_reg,
  mem_1415_sv2v_reg,mem_1414_sv2v_reg,mem_1413_sv2v_reg,mem_1412_sv2v_reg,
  mem_1411_sv2v_reg,mem_1410_sv2v_reg,mem_1409_sv2v_reg,mem_1408_sv2v_reg,mem_1407_sv2v_reg,
  mem_1406_sv2v_reg,mem_1405_sv2v_reg,mem_1404_sv2v_reg,mem_1403_sv2v_reg,
  mem_1402_sv2v_reg,mem_1401_sv2v_reg,mem_1400_sv2v_reg,mem_1399_sv2v_reg,
  mem_1398_sv2v_reg,mem_1397_sv2v_reg,mem_1396_sv2v_reg,mem_1395_sv2v_reg,mem_1394_sv2v_reg,
  mem_1393_sv2v_reg,mem_1392_sv2v_reg,mem_1391_sv2v_reg,mem_1390_sv2v_reg,
  mem_1389_sv2v_reg,mem_1388_sv2v_reg,mem_1387_sv2v_reg,mem_1386_sv2v_reg,mem_1385_sv2v_reg,
  mem_1384_sv2v_reg,mem_1383_sv2v_reg,mem_1382_sv2v_reg,mem_1381_sv2v_reg,
  mem_1380_sv2v_reg,mem_1379_sv2v_reg,mem_1378_sv2v_reg,mem_1377_sv2v_reg,mem_1376_sv2v_reg,
  mem_1375_sv2v_reg,mem_1374_sv2v_reg,mem_1373_sv2v_reg,mem_1372_sv2v_reg,
  mem_1371_sv2v_reg,mem_1370_sv2v_reg,mem_1369_sv2v_reg,mem_1368_sv2v_reg,mem_1367_sv2v_reg,
  mem_1366_sv2v_reg,mem_1365_sv2v_reg,mem_1364_sv2v_reg,mem_1363_sv2v_reg,
  mem_1362_sv2v_reg,mem_1361_sv2v_reg,mem_1360_sv2v_reg,mem_1359_sv2v_reg,
  mem_1358_sv2v_reg,mem_1357_sv2v_reg,mem_1356_sv2v_reg,mem_1355_sv2v_reg,mem_1354_sv2v_reg,
  mem_1353_sv2v_reg,mem_1352_sv2v_reg,mem_1351_sv2v_reg,mem_1350_sv2v_reg,
  mem_1349_sv2v_reg,mem_1348_sv2v_reg,mem_1347_sv2v_reg,mem_1346_sv2v_reg,mem_1345_sv2v_reg,
  mem_1344_sv2v_reg,mem_1343_sv2v_reg,mem_1342_sv2v_reg,mem_1341_sv2v_reg,
  mem_1340_sv2v_reg,mem_1339_sv2v_reg,mem_1338_sv2v_reg,mem_1337_sv2v_reg,mem_1336_sv2v_reg,
  mem_1335_sv2v_reg,mem_1334_sv2v_reg,mem_1333_sv2v_reg,mem_1332_sv2v_reg,
  mem_1331_sv2v_reg,mem_1330_sv2v_reg,mem_1329_sv2v_reg,mem_1328_sv2v_reg,mem_1327_sv2v_reg,
  mem_1326_sv2v_reg,mem_1325_sv2v_reg,mem_1324_sv2v_reg,mem_1323_sv2v_reg,
  mem_1322_sv2v_reg,mem_1321_sv2v_reg,mem_1320_sv2v_reg,mem_1319_sv2v_reg,
  mem_1318_sv2v_reg,mem_1317_sv2v_reg,mem_1316_sv2v_reg,mem_1315_sv2v_reg,mem_1314_sv2v_reg,
  mem_1313_sv2v_reg,mem_1312_sv2v_reg,mem_1311_sv2v_reg,mem_1310_sv2v_reg,
  mem_1309_sv2v_reg,mem_1308_sv2v_reg,mem_1307_sv2v_reg,mem_1306_sv2v_reg,mem_1305_sv2v_reg,
  mem_1304_sv2v_reg,mem_1303_sv2v_reg,mem_1302_sv2v_reg,mem_1301_sv2v_reg,
  mem_1300_sv2v_reg,mem_1299_sv2v_reg,mem_1298_sv2v_reg,mem_1297_sv2v_reg,mem_1296_sv2v_reg,
  mem_1295_sv2v_reg,mem_1294_sv2v_reg,mem_1293_sv2v_reg,mem_1292_sv2v_reg,
  mem_1291_sv2v_reg,mem_1290_sv2v_reg,mem_1289_sv2v_reg,mem_1288_sv2v_reg,mem_1287_sv2v_reg,
  mem_1286_sv2v_reg,mem_1285_sv2v_reg,mem_1284_sv2v_reg,mem_1283_sv2v_reg,
  mem_1282_sv2v_reg,mem_1281_sv2v_reg,mem_1280_sv2v_reg,mem_1279_sv2v_reg,
  mem_1278_sv2v_reg,mem_1277_sv2v_reg,mem_1276_sv2v_reg,mem_1275_sv2v_reg,mem_1274_sv2v_reg,
  mem_1273_sv2v_reg,mem_1272_sv2v_reg,mem_1271_sv2v_reg,mem_1270_sv2v_reg,
  mem_1269_sv2v_reg,mem_1268_sv2v_reg,mem_1267_sv2v_reg,mem_1266_sv2v_reg,mem_1265_sv2v_reg,
  mem_1264_sv2v_reg,mem_1263_sv2v_reg,mem_1262_sv2v_reg,mem_1261_sv2v_reg,
  mem_1260_sv2v_reg,mem_1259_sv2v_reg,mem_1258_sv2v_reg,mem_1257_sv2v_reg,mem_1256_sv2v_reg,
  mem_1255_sv2v_reg,mem_1254_sv2v_reg,mem_1253_sv2v_reg,mem_1252_sv2v_reg,
  mem_1251_sv2v_reg,mem_1250_sv2v_reg,mem_1249_sv2v_reg,mem_1248_sv2v_reg,mem_1247_sv2v_reg,
  mem_1246_sv2v_reg,mem_1245_sv2v_reg,mem_1244_sv2v_reg,mem_1243_sv2v_reg,
  mem_1242_sv2v_reg,mem_1241_sv2v_reg,mem_1240_sv2v_reg,mem_1239_sv2v_reg,
  mem_1238_sv2v_reg,mem_1237_sv2v_reg,mem_1236_sv2v_reg,mem_1235_sv2v_reg,mem_1234_sv2v_reg,
  mem_1233_sv2v_reg,mem_1232_sv2v_reg,mem_1231_sv2v_reg,mem_1230_sv2v_reg,
  mem_1229_sv2v_reg,mem_1228_sv2v_reg,mem_1227_sv2v_reg,mem_1226_sv2v_reg,mem_1225_sv2v_reg,
  mem_1224_sv2v_reg,mem_1223_sv2v_reg,mem_1222_sv2v_reg,mem_1221_sv2v_reg,
  mem_1220_sv2v_reg,mem_1219_sv2v_reg,mem_1218_sv2v_reg,mem_1217_sv2v_reg,mem_1216_sv2v_reg,
  mem_1215_sv2v_reg,mem_1214_sv2v_reg,mem_1213_sv2v_reg,mem_1212_sv2v_reg,
  mem_1211_sv2v_reg,mem_1210_sv2v_reg,mem_1209_sv2v_reg,mem_1208_sv2v_reg,mem_1207_sv2v_reg,
  mem_1206_sv2v_reg,mem_1205_sv2v_reg,mem_1204_sv2v_reg,mem_1203_sv2v_reg,
  mem_1202_sv2v_reg,mem_1201_sv2v_reg,mem_1200_sv2v_reg,mem_1199_sv2v_reg,
  mem_1198_sv2v_reg,mem_1197_sv2v_reg,mem_1196_sv2v_reg,mem_1195_sv2v_reg,mem_1194_sv2v_reg,
  mem_1193_sv2v_reg,mem_1192_sv2v_reg,mem_1191_sv2v_reg,mem_1190_sv2v_reg,
  mem_1189_sv2v_reg,mem_1188_sv2v_reg,mem_1187_sv2v_reg,mem_1186_sv2v_reg,mem_1185_sv2v_reg,
  mem_1184_sv2v_reg,mem_1183_sv2v_reg,mem_1182_sv2v_reg,mem_1181_sv2v_reg,
  mem_1180_sv2v_reg,mem_1179_sv2v_reg,mem_1178_sv2v_reg,mem_1177_sv2v_reg,mem_1176_sv2v_reg,
  mem_1175_sv2v_reg,mem_1174_sv2v_reg,mem_1173_sv2v_reg,mem_1172_sv2v_reg,
  mem_1171_sv2v_reg,mem_1170_sv2v_reg,mem_1169_sv2v_reg,mem_1168_sv2v_reg,mem_1167_sv2v_reg,
  mem_1166_sv2v_reg,mem_1165_sv2v_reg,mem_1164_sv2v_reg,mem_1163_sv2v_reg,
  mem_1162_sv2v_reg,mem_1161_sv2v_reg,mem_1160_sv2v_reg,mem_1159_sv2v_reg,
  mem_1158_sv2v_reg,mem_1157_sv2v_reg,mem_1156_sv2v_reg,mem_1155_sv2v_reg,mem_1154_sv2v_reg,
  mem_1153_sv2v_reg,mem_1152_sv2v_reg,mem_1151_sv2v_reg,mem_1150_sv2v_reg,
  mem_1149_sv2v_reg,mem_1148_sv2v_reg,mem_1147_sv2v_reg,mem_1146_sv2v_reg,mem_1145_sv2v_reg,
  mem_1144_sv2v_reg,mem_1143_sv2v_reg,mem_1142_sv2v_reg,mem_1141_sv2v_reg,
  mem_1140_sv2v_reg,mem_1139_sv2v_reg,mem_1138_sv2v_reg,mem_1137_sv2v_reg,mem_1136_sv2v_reg,
  mem_1135_sv2v_reg,mem_1134_sv2v_reg,mem_1133_sv2v_reg,mem_1132_sv2v_reg,
  mem_1131_sv2v_reg,mem_1130_sv2v_reg,mem_1129_sv2v_reg,mem_1128_sv2v_reg,mem_1127_sv2v_reg,
  mem_1126_sv2v_reg,mem_1125_sv2v_reg,mem_1124_sv2v_reg,mem_1123_sv2v_reg,
  mem_1122_sv2v_reg,mem_1121_sv2v_reg,mem_1120_sv2v_reg,mem_1119_sv2v_reg,
  mem_1118_sv2v_reg,mem_1117_sv2v_reg,mem_1116_sv2v_reg,mem_1115_sv2v_reg,mem_1114_sv2v_reg,
  mem_1113_sv2v_reg,mem_1112_sv2v_reg,mem_1111_sv2v_reg,mem_1110_sv2v_reg,
  mem_1109_sv2v_reg,mem_1108_sv2v_reg,mem_1107_sv2v_reg,mem_1106_sv2v_reg,mem_1105_sv2v_reg,
  mem_1104_sv2v_reg,mem_1103_sv2v_reg,mem_1102_sv2v_reg,mem_1101_sv2v_reg,
  mem_1100_sv2v_reg,mem_1099_sv2v_reg,mem_1098_sv2v_reg,mem_1097_sv2v_reg,mem_1096_sv2v_reg,
  mem_1095_sv2v_reg,mem_1094_sv2v_reg,mem_1093_sv2v_reg,mem_1092_sv2v_reg,
  mem_1091_sv2v_reg,mem_1090_sv2v_reg,mem_1089_sv2v_reg,mem_1088_sv2v_reg,mem_1087_sv2v_reg,
  mem_1086_sv2v_reg,mem_1085_sv2v_reg,mem_1084_sv2v_reg,mem_1083_sv2v_reg,
  mem_1082_sv2v_reg,mem_1081_sv2v_reg,mem_1080_sv2v_reg,mem_1079_sv2v_reg,
  mem_1078_sv2v_reg,mem_1077_sv2v_reg,mem_1076_sv2v_reg,mem_1075_sv2v_reg,mem_1074_sv2v_reg,
  mem_1073_sv2v_reg,mem_1072_sv2v_reg,mem_1071_sv2v_reg,mem_1070_sv2v_reg,
  mem_1069_sv2v_reg,mem_1068_sv2v_reg,mem_1067_sv2v_reg,mem_1066_sv2v_reg,mem_1065_sv2v_reg,
  mem_1064_sv2v_reg,mem_1063_sv2v_reg,mem_1062_sv2v_reg,mem_1061_sv2v_reg,
  mem_1060_sv2v_reg,mem_1059_sv2v_reg,mem_1058_sv2v_reg,mem_1057_sv2v_reg,mem_1056_sv2v_reg,
  mem_1055_sv2v_reg,mem_1054_sv2v_reg,mem_1053_sv2v_reg,mem_1052_sv2v_reg,
  mem_1051_sv2v_reg,mem_1050_sv2v_reg,mem_1049_sv2v_reg,mem_1048_sv2v_reg,mem_1047_sv2v_reg,
  mem_1046_sv2v_reg,mem_1045_sv2v_reg,mem_1044_sv2v_reg,mem_1043_sv2v_reg,
  mem_1042_sv2v_reg,mem_1041_sv2v_reg,mem_1040_sv2v_reg,mem_1039_sv2v_reg,
  mem_1038_sv2v_reg,mem_1037_sv2v_reg,mem_1036_sv2v_reg,mem_1035_sv2v_reg,mem_1034_sv2v_reg,
  mem_1033_sv2v_reg,mem_1032_sv2v_reg,mem_1031_sv2v_reg,mem_1030_sv2v_reg,
  mem_1029_sv2v_reg,mem_1028_sv2v_reg,mem_1027_sv2v_reg,mem_1026_sv2v_reg,mem_1025_sv2v_reg,
  mem_1024_sv2v_reg,mem_1023_sv2v_reg,mem_1022_sv2v_reg,mem_1021_sv2v_reg,
  mem_1020_sv2v_reg,mem_1019_sv2v_reg,mem_1018_sv2v_reg,mem_1017_sv2v_reg,mem_1016_sv2v_reg,
  mem_1015_sv2v_reg,mem_1014_sv2v_reg,mem_1013_sv2v_reg,mem_1012_sv2v_reg,
  mem_1011_sv2v_reg,mem_1010_sv2v_reg,mem_1009_sv2v_reg,mem_1008_sv2v_reg,mem_1007_sv2v_reg,
  mem_1006_sv2v_reg,mem_1005_sv2v_reg,mem_1004_sv2v_reg,mem_1003_sv2v_reg,
  mem_1002_sv2v_reg,mem_1001_sv2v_reg,mem_1000_sv2v_reg,mem_999_sv2v_reg,mem_998_sv2v_reg,
  mem_997_sv2v_reg,mem_996_sv2v_reg,mem_995_sv2v_reg,mem_994_sv2v_reg,
  mem_993_sv2v_reg,mem_992_sv2v_reg,mem_991_sv2v_reg,mem_990_sv2v_reg,mem_989_sv2v_reg,
  mem_988_sv2v_reg,mem_987_sv2v_reg,mem_986_sv2v_reg,mem_985_sv2v_reg,mem_984_sv2v_reg,
  mem_983_sv2v_reg,mem_982_sv2v_reg,mem_981_sv2v_reg,mem_980_sv2v_reg,
  mem_979_sv2v_reg,mem_978_sv2v_reg,mem_977_sv2v_reg,mem_976_sv2v_reg,mem_975_sv2v_reg,
  mem_974_sv2v_reg,mem_973_sv2v_reg,mem_972_sv2v_reg,mem_971_sv2v_reg,mem_970_sv2v_reg,
  mem_969_sv2v_reg,mem_968_sv2v_reg,mem_967_sv2v_reg,mem_966_sv2v_reg,
  mem_965_sv2v_reg,mem_964_sv2v_reg,mem_963_sv2v_reg,mem_962_sv2v_reg,mem_961_sv2v_reg,
  mem_960_sv2v_reg,mem_959_sv2v_reg,mem_958_sv2v_reg,mem_957_sv2v_reg,mem_956_sv2v_reg,
  mem_955_sv2v_reg,mem_954_sv2v_reg,mem_953_sv2v_reg,mem_952_sv2v_reg,mem_951_sv2v_reg,
  mem_950_sv2v_reg,mem_949_sv2v_reg,mem_948_sv2v_reg,mem_947_sv2v_reg,
  mem_946_sv2v_reg,mem_945_sv2v_reg,mem_944_sv2v_reg,mem_943_sv2v_reg,mem_942_sv2v_reg,
  mem_941_sv2v_reg,mem_940_sv2v_reg,mem_939_sv2v_reg,mem_938_sv2v_reg,mem_937_sv2v_reg,
  mem_936_sv2v_reg,mem_935_sv2v_reg,mem_934_sv2v_reg,mem_933_sv2v_reg,
  mem_932_sv2v_reg,mem_931_sv2v_reg,mem_930_sv2v_reg,mem_929_sv2v_reg,mem_928_sv2v_reg,
  mem_927_sv2v_reg,mem_926_sv2v_reg,mem_925_sv2v_reg,mem_924_sv2v_reg,mem_923_sv2v_reg,
  mem_922_sv2v_reg,mem_921_sv2v_reg,mem_920_sv2v_reg,mem_919_sv2v_reg,mem_918_sv2v_reg,
  mem_917_sv2v_reg,mem_916_sv2v_reg,mem_915_sv2v_reg,mem_914_sv2v_reg,
  mem_913_sv2v_reg,mem_912_sv2v_reg,mem_911_sv2v_reg,mem_910_sv2v_reg,mem_909_sv2v_reg,
  mem_908_sv2v_reg,mem_907_sv2v_reg,mem_906_sv2v_reg,mem_905_sv2v_reg,mem_904_sv2v_reg,
  mem_903_sv2v_reg,mem_902_sv2v_reg,mem_901_sv2v_reg,mem_900_sv2v_reg,
  mem_899_sv2v_reg,mem_898_sv2v_reg,mem_897_sv2v_reg,mem_896_sv2v_reg,mem_895_sv2v_reg,
  mem_894_sv2v_reg,mem_893_sv2v_reg,mem_892_sv2v_reg,mem_891_sv2v_reg,mem_890_sv2v_reg,
  mem_889_sv2v_reg,mem_888_sv2v_reg,mem_887_sv2v_reg,mem_886_sv2v_reg,
  mem_885_sv2v_reg,mem_884_sv2v_reg,mem_883_sv2v_reg,mem_882_sv2v_reg,mem_881_sv2v_reg,
  mem_880_sv2v_reg,mem_879_sv2v_reg,mem_878_sv2v_reg,mem_877_sv2v_reg,mem_876_sv2v_reg,
  mem_875_sv2v_reg,mem_874_sv2v_reg,mem_873_sv2v_reg,mem_872_sv2v_reg,mem_871_sv2v_reg,
  mem_870_sv2v_reg,mem_869_sv2v_reg,mem_868_sv2v_reg,mem_867_sv2v_reg,
  mem_866_sv2v_reg,mem_865_sv2v_reg,mem_864_sv2v_reg,mem_863_sv2v_reg,mem_862_sv2v_reg,
  mem_861_sv2v_reg,mem_860_sv2v_reg,mem_859_sv2v_reg,mem_858_sv2v_reg,mem_857_sv2v_reg,
  mem_856_sv2v_reg,mem_855_sv2v_reg,mem_854_sv2v_reg,mem_853_sv2v_reg,
  mem_852_sv2v_reg,mem_851_sv2v_reg,mem_850_sv2v_reg,mem_849_sv2v_reg,mem_848_sv2v_reg,
  mem_847_sv2v_reg,mem_846_sv2v_reg,mem_845_sv2v_reg,mem_844_sv2v_reg,mem_843_sv2v_reg,
  mem_842_sv2v_reg,mem_841_sv2v_reg,mem_840_sv2v_reg,mem_839_sv2v_reg,mem_838_sv2v_reg,
  mem_837_sv2v_reg,mem_836_sv2v_reg,mem_835_sv2v_reg,mem_834_sv2v_reg,
  mem_833_sv2v_reg,mem_832_sv2v_reg,mem_831_sv2v_reg,mem_830_sv2v_reg,mem_829_sv2v_reg,
  mem_828_sv2v_reg,mem_827_sv2v_reg,mem_826_sv2v_reg,mem_825_sv2v_reg,mem_824_sv2v_reg,
  mem_823_sv2v_reg,mem_822_sv2v_reg,mem_821_sv2v_reg,mem_820_sv2v_reg,
  mem_819_sv2v_reg,mem_818_sv2v_reg,mem_817_sv2v_reg,mem_816_sv2v_reg,mem_815_sv2v_reg,
  mem_814_sv2v_reg,mem_813_sv2v_reg,mem_812_sv2v_reg,mem_811_sv2v_reg,mem_810_sv2v_reg,
  mem_809_sv2v_reg,mem_808_sv2v_reg,mem_807_sv2v_reg,mem_806_sv2v_reg,
  mem_805_sv2v_reg,mem_804_sv2v_reg,mem_803_sv2v_reg,mem_802_sv2v_reg,mem_801_sv2v_reg,
  mem_800_sv2v_reg,mem_799_sv2v_reg,mem_798_sv2v_reg,mem_797_sv2v_reg,mem_796_sv2v_reg,
  mem_795_sv2v_reg,mem_794_sv2v_reg,mem_793_sv2v_reg,mem_792_sv2v_reg,mem_791_sv2v_reg,
  mem_790_sv2v_reg,mem_789_sv2v_reg,mem_788_sv2v_reg,mem_787_sv2v_reg,
  mem_786_sv2v_reg,mem_785_sv2v_reg,mem_784_sv2v_reg,mem_783_sv2v_reg,mem_782_sv2v_reg,
  mem_781_sv2v_reg,mem_780_sv2v_reg,mem_779_sv2v_reg,mem_778_sv2v_reg,mem_777_sv2v_reg,
  mem_776_sv2v_reg,mem_775_sv2v_reg,mem_774_sv2v_reg,mem_773_sv2v_reg,
  mem_772_sv2v_reg,mem_771_sv2v_reg,mem_770_sv2v_reg,mem_769_sv2v_reg,mem_768_sv2v_reg,
  mem_767_sv2v_reg,mem_766_sv2v_reg,mem_765_sv2v_reg,mem_764_sv2v_reg,mem_763_sv2v_reg,
  mem_762_sv2v_reg,mem_761_sv2v_reg,mem_760_sv2v_reg,mem_759_sv2v_reg,mem_758_sv2v_reg,
  mem_757_sv2v_reg,mem_756_sv2v_reg,mem_755_sv2v_reg,mem_754_sv2v_reg,
  mem_753_sv2v_reg,mem_752_sv2v_reg,mem_751_sv2v_reg,mem_750_sv2v_reg,mem_749_sv2v_reg,
  mem_748_sv2v_reg,mem_747_sv2v_reg,mem_746_sv2v_reg,mem_745_sv2v_reg,mem_744_sv2v_reg,
  mem_743_sv2v_reg,mem_742_sv2v_reg,mem_741_sv2v_reg,mem_740_sv2v_reg,
  mem_739_sv2v_reg,mem_738_sv2v_reg,mem_737_sv2v_reg,mem_736_sv2v_reg,mem_735_sv2v_reg,
  mem_734_sv2v_reg,mem_733_sv2v_reg,mem_732_sv2v_reg,mem_731_sv2v_reg,mem_730_sv2v_reg,
  mem_729_sv2v_reg,mem_728_sv2v_reg,mem_727_sv2v_reg,mem_726_sv2v_reg,
  mem_725_sv2v_reg,mem_724_sv2v_reg,mem_723_sv2v_reg,mem_722_sv2v_reg,mem_721_sv2v_reg,
  mem_720_sv2v_reg,mem_719_sv2v_reg,mem_718_sv2v_reg,mem_717_sv2v_reg,mem_716_sv2v_reg,
  mem_715_sv2v_reg,mem_714_sv2v_reg,mem_713_sv2v_reg,mem_712_sv2v_reg,mem_711_sv2v_reg,
  mem_710_sv2v_reg,mem_709_sv2v_reg,mem_708_sv2v_reg,mem_707_sv2v_reg,
  mem_706_sv2v_reg,mem_705_sv2v_reg,mem_704_sv2v_reg,mem_703_sv2v_reg,mem_702_sv2v_reg,
  mem_701_sv2v_reg,mem_700_sv2v_reg,mem_699_sv2v_reg,mem_698_sv2v_reg,mem_697_sv2v_reg,
  mem_696_sv2v_reg,mem_695_sv2v_reg,mem_694_sv2v_reg,mem_693_sv2v_reg,
  mem_692_sv2v_reg,mem_691_sv2v_reg,mem_690_sv2v_reg,mem_689_sv2v_reg,mem_688_sv2v_reg,
  mem_687_sv2v_reg,mem_686_sv2v_reg,mem_685_sv2v_reg,mem_684_sv2v_reg,mem_683_sv2v_reg,
  mem_682_sv2v_reg,mem_681_sv2v_reg,mem_680_sv2v_reg,mem_679_sv2v_reg,mem_678_sv2v_reg,
  mem_677_sv2v_reg,mem_676_sv2v_reg,mem_675_sv2v_reg,mem_674_sv2v_reg,
  mem_673_sv2v_reg,mem_672_sv2v_reg,mem_671_sv2v_reg,mem_670_sv2v_reg,mem_669_sv2v_reg,
  mem_668_sv2v_reg,mem_667_sv2v_reg,mem_666_sv2v_reg,mem_665_sv2v_reg,mem_664_sv2v_reg,
  mem_663_sv2v_reg,mem_662_sv2v_reg,mem_661_sv2v_reg,mem_660_sv2v_reg,
  mem_659_sv2v_reg,mem_658_sv2v_reg,mem_657_sv2v_reg,mem_656_sv2v_reg,mem_655_sv2v_reg,
  mem_654_sv2v_reg,mem_653_sv2v_reg,mem_652_sv2v_reg,mem_651_sv2v_reg,mem_650_sv2v_reg,
  mem_649_sv2v_reg,mem_648_sv2v_reg,mem_647_sv2v_reg,mem_646_sv2v_reg,
  mem_645_sv2v_reg,mem_644_sv2v_reg,mem_643_sv2v_reg,mem_642_sv2v_reg,mem_641_sv2v_reg,
  mem_640_sv2v_reg,mem_639_sv2v_reg,mem_638_sv2v_reg,mem_637_sv2v_reg,mem_636_sv2v_reg,
  mem_635_sv2v_reg,mem_634_sv2v_reg,mem_633_sv2v_reg,mem_632_sv2v_reg,mem_631_sv2v_reg,
  mem_630_sv2v_reg,mem_629_sv2v_reg,mem_628_sv2v_reg,mem_627_sv2v_reg,
  mem_626_sv2v_reg,mem_625_sv2v_reg,mem_624_sv2v_reg,mem_623_sv2v_reg,mem_622_sv2v_reg,
  mem_621_sv2v_reg,mem_620_sv2v_reg,mem_619_sv2v_reg,mem_618_sv2v_reg,mem_617_sv2v_reg,
  mem_616_sv2v_reg,mem_615_sv2v_reg,mem_614_sv2v_reg,mem_613_sv2v_reg,
  mem_612_sv2v_reg,mem_611_sv2v_reg,mem_610_sv2v_reg,mem_609_sv2v_reg,mem_608_sv2v_reg,
  mem_607_sv2v_reg,mem_606_sv2v_reg,mem_605_sv2v_reg,mem_604_sv2v_reg,mem_603_sv2v_reg,
  mem_602_sv2v_reg,mem_601_sv2v_reg,mem_600_sv2v_reg,mem_599_sv2v_reg,mem_598_sv2v_reg,
  mem_597_sv2v_reg,mem_596_sv2v_reg,mem_595_sv2v_reg,mem_594_sv2v_reg,
  mem_593_sv2v_reg,mem_592_sv2v_reg,mem_591_sv2v_reg,mem_590_sv2v_reg,mem_589_sv2v_reg,
  mem_588_sv2v_reg,mem_587_sv2v_reg,mem_586_sv2v_reg,mem_585_sv2v_reg,mem_584_sv2v_reg,
  mem_583_sv2v_reg,mem_582_sv2v_reg,mem_581_sv2v_reg,mem_580_sv2v_reg,
  mem_579_sv2v_reg,mem_578_sv2v_reg,mem_577_sv2v_reg,mem_576_sv2v_reg,mem_575_sv2v_reg,
  mem_574_sv2v_reg,mem_573_sv2v_reg,mem_572_sv2v_reg,mem_571_sv2v_reg,mem_570_sv2v_reg,
  mem_569_sv2v_reg,mem_568_sv2v_reg,mem_567_sv2v_reg,mem_566_sv2v_reg,
  mem_565_sv2v_reg,mem_564_sv2v_reg,mem_563_sv2v_reg,mem_562_sv2v_reg,mem_561_sv2v_reg,
  mem_560_sv2v_reg,mem_559_sv2v_reg,mem_558_sv2v_reg,mem_557_sv2v_reg,mem_556_sv2v_reg,
  mem_555_sv2v_reg,mem_554_sv2v_reg,mem_553_sv2v_reg,mem_552_sv2v_reg,mem_551_sv2v_reg,
  mem_550_sv2v_reg,mem_549_sv2v_reg,mem_548_sv2v_reg,mem_547_sv2v_reg,
  mem_546_sv2v_reg,mem_545_sv2v_reg,mem_544_sv2v_reg,mem_543_sv2v_reg,mem_542_sv2v_reg,
  mem_541_sv2v_reg,mem_540_sv2v_reg,mem_539_sv2v_reg,mem_538_sv2v_reg,mem_537_sv2v_reg,
  mem_536_sv2v_reg,mem_535_sv2v_reg,mem_534_sv2v_reg,mem_533_sv2v_reg,
  mem_532_sv2v_reg,mem_531_sv2v_reg,mem_530_sv2v_reg,mem_529_sv2v_reg,mem_528_sv2v_reg,
  mem_527_sv2v_reg,mem_526_sv2v_reg,mem_525_sv2v_reg,mem_524_sv2v_reg,mem_523_sv2v_reg,
  mem_522_sv2v_reg,mem_521_sv2v_reg,mem_520_sv2v_reg,mem_519_sv2v_reg,mem_518_sv2v_reg,
  mem_517_sv2v_reg,mem_516_sv2v_reg,mem_515_sv2v_reg,mem_514_sv2v_reg,
  mem_513_sv2v_reg,mem_512_sv2v_reg,mem_511_sv2v_reg,mem_510_sv2v_reg,mem_509_sv2v_reg,
  mem_508_sv2v_reg,mem_507_sv2v_reg,mem_506_sv2v_reg,mem_505_sv2v_reg,mem_504_sv2v_reg,
  mem_503_sv2v_reg,mem_502_sv2v_reg,mem_501_sv2v_reg,mem_500_sv2v_reg,
  mem_499_sv2v_reg,mem_498_sv2v_reg,mem_497_sv2v_reg,mem_496_sv2v_reg,mem_495_sv2v_reg,
  mem_494_sv2v_reg,mem_493_sv2v_reg,mem_492_sv2v_reg,mem_491_sv2v_reg,mem_490_sv2v_reg,
  mem_489_sv2v_reg,mem_488_sv2v_reg,mem_487_sv2v_reg,mem_486_sv2v_reg,
  mem_485_sv2v_reg,mem_484_sv2v_reg,mem_483_sv2v_reg,mem_482_sv2v_reg,mem_481_sv2v_reg,
  mem_480_sv2v_reg,mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,mem_476_sv2v_reg,
  mem_475_sv2v_reg,mem_474_sv2v_reg,mem_473_sv2v_reg,mem_472_sv2v_reg,mem_471_sv2v_reg,
  mem_470_sv2v_reg,mem_469_sv2v_reg,mem_468_sv2v_reg,mem_467_sv2v_reg,
  mem_466_sv2v_reg,mem_465_sv2v_reg,mem_464_sv2v_reg,mem_463_sv2v_reg,mem_462_sv2v_reg,
  mem_461_sv2v_reg,mem_460_sv2v_reg,mem_459_sv2v_reg,mem_458_sv2v_reg,mem_457_sv2v_reg,
  mem_456_sv2v_reg,mem_455_sv2v_reg,mem_454_sv2v_reg,mem_453_sv2v_reg,
  mem_452_sv2v_reg,mem_451_sv2v_reg,mem_450_sv2v_reg,mem_449_sv2v_reg,mem_448_sv2v_reg,
  mem_447_sv2v_reg,mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,mem_443_sv2v_reg,
  mem_442_sv2v_reg,mem_441_sv2v_reg,mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,
  mem_437_sv2v_reg,mem_436_sv2v_reg,mem_435_sv2v_reg,mem_434_sv2v_reg,
  mem_433_sv2v_reg,mem_432_sv2v_reg,mem_431_sv2v_reg,mem_430_sv2v_reg,mem_429_sv2v_reg,
  mem_428_sv2v_reg,mem_427_sv2v_reg,mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,
  mem_423_sv2v_reg,mem_422_sv2v_reg,mem_421_sv2v_reg,mem_420_sv2v_reg,
  mem_419_sv2v_reg,mem_418_sv2v_reg,mem_417_sv2v_reg,mem_416_sv2v_reg,mem_415_sv2v_reg,
  mem_414_sv2v_reg,mem_413_sv2v_reg,mem_412_sv2v_reg,mem_411_sv2v_reg,mem_410_sv2v_reg,
  mem_409_sv2v_reg,mem_408_sv2v_reg,mem_407_sv2v_reg,mem_406_sv2v_reg,
  mem_405_sv2v_reg,mem_404_sv2v_reg,mem_403_sv2v_reg,mem_402_sv2v_reg,mem_401_sv2v_reg,
  mem_400_sv2v_reg,mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,mem_396_sv2v_reg,
  mem_395_sv2v_reg,mem_394_sv2v_reg,mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,
  mem_390_sv2v_reg,mem_389_sv2v_reg,mem_388_sv2v_reg,mem_387_sv2v_reg,
  mem_386_sv2v_reg,mem_385_sv2v_reg,mem_384_sv2v_reg,mem_383_sv2v_reg,mem_382_sv2v_reg,
  mem_381_sv2v_reg,mem_380_sv2v_reg,mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,
  mem_376_sv2v_reg,mem_375_sv2v_reg,mem_374_sv2v_reg,mem_373_sv2v_reg,
  mem_372_sv2v_reg,mem_371_sv2v_reg,mem_370_sv2v_reg,mem_369_sv2v_reg,mem_368_sv2v_reg,
  mem_367_sv2v_reg,mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,mem_363_sv2v_reg,
  mem_362_sv2v_reg,mem_361_sv2v_reg,mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,
  mem_357_sv2v_reg,mem_356_sv2v_reg,mem_355_sv2v_reg,mem_354_sv2v_reg,
  mem_353_sv2v_reg,mem_352_sv2v_reg,mem_351_sv2v_reg,mem_350_sv2v_reg,mem_349_sv2v_reg,
  mem_348_sv2v_reg,mem_347_sv2v_reg,mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,
  mem_343_sv2v_reg,mem_342_sv2v_reg,mem_341_sv2v_reg,mem_340_sv2v_reg,
  mem_339_sv2v_reg,mem_338_sv2v_reg,mem_337_sv2v_reg,mem_336_sv2v_reg,mem_335_sv2v_reg,
  mem_334_sv2v_reg,mem_333_sv2v_reg,mem_332_sv2v_reg,mem_331_sv2v_reg,mem_330_sv2v_reg,
  mem_329_sv2v_reg,mem_328_sv2v_reg,mem_327_sv2v_reg,mem_326_sv2v_reg,
  mem_325_sv2v_reg,mem_324_sv2v_reg,mem_323_sv2v_reg,mem_322_sv2v_reg,mem_321_sv2v_reg,
  mem_320_sv2v_reg,mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,mem_316_sv2v_reg,
  mem_315_sv2v_reg,mem_314_sv2v_reg,mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,
  mem_310_sv2v_reg,mem_309_sv2v_reg,mem_308_sv2v_reg,mem_307_sv2v_reg,
  mem_306_sv2v_reg,mem_305_sv2v_reg,mem_304_sv2v_reg,mem_303_sv2v_reg,mem_302_sv2v_reg,
  mem_301_sv2v_reg,mem_300_sv2v_reg,mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,
  mem_296_sv2v_reg,mem_295_sv2v_reg,mem_294_sv2v_reg,mem_293_sv2v_reg,
  mem_292_sv2v_reg,mem_291_sv2v_reg,mem_290_sv2v_reg,mem_289_sv2v_reg,mem_288_sv2v_reg,
  mem_287_sv2v_reg,mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,mem_283_sv2v_reg,
  mem_282_sv2v_reg,mem_281_sv2v_reg,mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,
  mem_277_sv2v_reg,mem_276_sv2v_reg,mem_275_sv2v_reg,mem_274_sv2v_reg,
  mem_273_sv2v_reg,mem_272_sv2v_reg,mem_271_sv2v_reg,mem_270_sv2v_reg,mem_269_sv2v_reg,
  mem_268_sv2v_reg,mem_267_sv2v_reg,mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,
  mem_263_sv2v_reg,mem_262_sv2v_reg,mem_261_sv2v_reg,mem_260_sv2v_reg,
  mem_259_sv2v_reg,mem_258_sv2v_reg,mem_257_sv2v_reg,mem_256_sv2v_reg,mem_255_sv2v_reg,
  mem_254_sv2v_reg,mem_253_sv2v_reg,mem_252_sv2v_reg,mem_251_sv2v_reg,mem_250_sv2v_reg,
  mem_249_sv2v_reg,mem_248_sv2v_reg,mem_247_sv2v_reg,mem_246_sv2v_reg,
  mem_245_sv2v_reg,mem_244_sv2v_reg,mem_243_sv2v_reg,mem_242_sv2v_reg,mem_241_sv2v_reg,
  mem_240_sv2v_reg,mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,mem_236_sv2v_reg,
  mem_235_sv2v_reg,mem_234_sv2v_reg,mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,
  mem_230_sv2v_reg,mem_229_sv2v_reg,mem_228_sv2v_reg,mem_227_sv2v_reg,
  mem_226_sv2v_reg,mem_225_sv2v_reg,mem_224_sv2v_reg,mem_223_sv2v_reg,mem_222_sv2v_reg,
  mem_221_sv2v_reg,mem_220_sv2v_reg,mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,
  mem_216_sv2v_reg,mem_215_sv2v_reg,mem_214_sv2v_reg,mem_213_sv2v_reg,
  mem_212_sv2v_reg,mem_211_sv2v_reg,mem_210_sv2v_reg,mem_209_sv2v_reg,mem_208_sv2v_reg,
  mem_207_sv2v_reg,mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,mem_203_sv2v_reg,
  mem_202_sv2v_reg,mem_201_sv2v_reg,mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,
  mem_197_sv2v_reg,mem_196_sv2v_reg,mem_195_sv2v_reg,mem_194_sv2v_reg,
  mem_193_sv2v_reg,mem_192_sv2v_reg,mem_191_sv2v_reg,mem_190_sv2v_reg,mem_189_sv2v_reg,
  mem_188_sv2v_reg,mem_187_sv2v_reg,mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,
  mem_183_sv2v_reg,mem_182_sv2v_reg,mem_181_sv2v_reg,mem_180_sv2v_reg,
  mem_179_sv2v_reg,mem_178_sv2v_reg,mem_177_sv2v_reg,mem_176_sv2v_reg,mem_175_sv2v_reg,
  mem_174_sv2v_reg,mem_173_sv2v_reg,mem_172_sv2v_reg,mem_171_sv2v_reg,mem_170_sv2v_reg,
  mem_169_sv2v_reg,mem_168_sv2v_reg,mem_167_sv2v_reg,mem_166_sv2v_reg,
  mem_165_sv2v_reg,mem_164_sv2v_reg,mem_163_sv2v_reg,mem_162_sv2v_reg,mem_161_sv2v_reg,
  mem_160_sv2v_reg,mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,mem_156_sv2v_reg,
  mem_155_sv2v_reg,mem_154_sv2v_reg,mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,
  mem_150_sv2v_reg,mem_149_sv2v_reg,mem_148_sv2v_reg,mem_147_sv2v_reg,
  mem_146_sv2v_reg,mem_145_sv2v_reg,mem_144_sv2v_reg,mem_143_sv2v_reg,mem_142_sv2v_reg,
  mem_141_sv2v_reg,mem_140_sv2v_reg,mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,
  mem_136_sv2v_reg,mem_135_sv2v_reg,mem_134_sv2v_reg,mem_133_sv2v_reg,
  mem_132_sv2v_reg,mem_131_sv2v_reg,mem_130_sv2v_reg,mem_129_sv2v_reg,mem_128_sv2v_reg,
  mem_127_sv2v_reg,mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,mem_123_sv2v_reg,
  mem_122_sv2v_reg,mem_121_sv2v_reg,mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,
  mem_117_sv2v_reg,mem_116_sv2v_reg,mem_115_sv2v_reg,mem_114_sv2v_reg,
  mem_113_sv2v_reg,mem_112_sv2v_reg,mem_111_sv2v_reg,mem_110_sv2v_reg,mem_109_sv2v_reg,
  mem_108_sv2v_reg,mem_107_sv2v_reg,mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,
  mem_103_sv2v_reg,mem_102_sv2v_reg,mem_101_sv2v_reg,mem_100_sv2v_reg,
  mem_99_sv2v_reg,mem_98_sv2v_reg,mem_97_sv2v_reg,mem_96_sv2v_reg,mem_95_sv2v_reg,
  mem_94_sv2v_reg,mem_93_sv2v_reg,mem_92_sv2v_reg,mem_91_sv2v_reg,mem_90_sv2v_reg,
  mem_89_sv2v_reg,mem_88_sv2v_reg,mem_87_sv2v_reg,mem_86_sv2v_reg,mem_85_sv2v_reg,
  mem_84_sv2v_reg,mem_83_sv2v_reg,mem_82_sv2v_reg,mem_81_sv2v_reg,mem_80_sv2v_reg,
  mem_79_sv2v_reg,mem_78_sv2v_reg,mem_77_sv2v_reg,mem_76_sv2v_reg,mem_75_sv2v_reg,
  mem_74_sv2v_reg,mem_73_sv2v_reg,mem_72_sv2v_reg,mem_71_sv2v_reg,mem_70_sv2v_reg,
  mem_69_sv2v_reg,mem_68_sv2v_reg,mem_67_sv2v_reg,mem_66_sv2v_reg,mem_65_sv2v_reg,
  mem_64_sv2v_reg,mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,
  mem_59_sv2v_reg,mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,
  mem_54_sv2v_reg,mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,
  mem_49_sv2v_reg,mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,
  mem_44_sv2v_reg,mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,
  mem_39_sv2v_reg,mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,
  mem_34_sv2v_reg,mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,
  mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,
  mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,
  mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,
  mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,
  mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,
  mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign addr_r[6] = addr_r_6_sv2v_reg;
  assign addr_r[5] = addr_r_5_sv2v_reg;
  assign addr_r[4] = addr_r_4_sv2v_reg;
  assign addr_r[3] = addr_r_3_sv2v_reg;
  assign addr_r[2] = addr_r_2_sv2v_reg;
  assign addr_r[1] = addr_r_1_sv2v_reg;
  assign addr_r[0] = addr_r_0_sv2v_reg;
  assign mem[1919] = mem_1919_sv2v_reg;
  assign mem[1918] = mem_1918_sv2v_reg;
  assign mem[1917] = mem_1917_sv2v_reg;
  assign mem[1916] = mem_1916_sv2v_reg;
  assign mem[1915] = mem_1915_sv2v_reg;
  assign mem[1914] = mem_1914_sv2v_reg;
  assign mem[1913] = mem_1913_sv2v_reg;
  assign mem[1912] = mem_1912_sv2v_reg;
  assign mem[1911] = mem_1911_sv2v_reg;
  assign mem[1910] = mem_1910_sv2v_reg;
  assign mem[1909] = mem_1909_sv2v_reg;
  assign mem[1908] = mem_1908_sv2v_reg;
  assign mem[1907] = mem_1907_sv2v_reg;
  assign mem[1906] = mem_1906_sv2v_reg;
  assign mem[1905] = mem_1905_sv2v_reg;
  assign mem[1904] = mem_1904_sv2v_reg;
  assign mem[1903] = mem_1903_sv2v_reg;
  assign mem[1902] = mem_1902_sv2v_reg;
  assign mem[1901] = mem_1901_sv2v_reg;
  assign mem[1900] = mem_1900_sv2v_reg;
  assign mem[1899] = mem_1899_sv2v_reg;
  assign mem[1898] = mem_1898_sv2v_reg;
  assign mem[1897] = mem_1897_sv2v_reg;
  assign mem[1896] = mem_1896_sv2v_reg;
  assign mem[1895] = mem_1895_sv2v_reg;
  assign mem[1894] = mem_1894_sv2v_reg;
  assign mem[1893] = mem_1893_sv2v_reg;
  assign mem[1892] = mem_1892_sv2v_reg;
  assign mem[1891] = mem_1891_sv2v_reg;
  assign mem[1890] = mem_1890_sv2v_reg;
  assign mem[1889] = mem_1889_sv2v_reg;
  assign mem[1888] = mem_1888_sv2v_reg;
  assign mem[1887] = mem_1887_sv2v_reg;
  assign mem[1886] = mem_1886_sv2v_reg;
  assign mem[1885] = mem_1885_sv2v_reg;
  assign mem[1884] = mem_1884_sv2v_reg;
  assign mem[1883] = mem_1883_sv2v_reg;
  assign mem[1882] = mem_1882_sv2v_reg;
  assign mem[1881] = mem_1881_sv2v_reg;
  assign mem[1880] = mem_1880_sv2v_reg;
  assign mem[1879] = mem_1879_sv2v_reg;
  assign mem[1878] = mem_1878_sv2v_reg;
  assign mem[1877] = mem_1877_sv2v_reg;
  assign mem[1876] = mem_1876_sv2v_reg;
  assign mem[1875] = mem_1875_sv2v_reg;
  assign mem[1874] = mem_1874_sv2v_reg;
  assign mem[1873] = mem_1873_sv2v_reg;
  assign mem[1872] = mem_1872_sv2v_reg;
  assign mem[1871] = mem_1871_sv2v_reg;
  assign mem[1870] = mem_1870_sv2v_reg;
  assign mem[1869] = mem_1869_sv2v_reg;
  assign mem[1868] = mem_1868_sv2v_reg;
  assign mem[1867] = mem_1867_sv2v_reg;
  assign mem[1866] = mem_1866_sv2v_reg;
  assign mem[1865] = mem_1865_sv2v_reg;
  assign mem[1864] = mem_1864_sv2v_reg;
  assign mem[1863] = mem_1863_sv2v_reg;
  assign mem[1862] = mem_1862_sv2v_reg;
  assign mem[1861] = mem_1861_sv2v_reg;
  assign mem[1860] = mem_1860_sv2v_reg;
  assign mem[1859] = mem_1859_sv2v_reg;
  assign mem[1858] = mem_1858_sv2v_reg;
  assign mem[1857] = mem_1857_sv2v_reg;
  assign mem[1856] = mem_1856_sv2v_reg;
  assign mem[1855] = mem_1855_sv2v_reg;
  assign mem[1854] = mem_1854_sv2v_reg;
  assign mem[1853] = mem_1853_sv2v_reg;
  assign mem[1852] = mem_1852_sv2v_reg;
  assign mem[1851] = mem_1851_sv2v_reg;
  assign mem[1850] = mem_1850_sv2v_reg;
  assign mem[1849] = mem_1849_sv2v_reg;
  assign mem[1848] = mem_1848_sv2v_reg;
  assign mem[1847] = mem_1847_sv2v_reg;
  assign mem[1846] = mem_1846_sv2v_reg;
  assign mem[1845] = mem_1845_sv2v_reg;
  assign mem[1844] = mem_1844_sv2v_reg;
  assign mem[1843] = mem_1843_sv2v_reg;
  assign mem[1842] = mem_1842_sv2v_reg;
  assign mem[1841] = mem_1841_sv2v_reg;
  assign mem[1840] = mem_1840_sv2v_reg;
  assign mem[1839] = mem_1839_sv2v_reg;
  assign mem[1838] = mem_1838_sv2v_reg;
  assign mem[1837] = mem_1837_sv2v_reg;
  assign mem[1836] = mem_1836_sv2v_reg;
  assign mem[1835] = mem_1835_sv2v_reg;
  assign mem[1834] = mem_1834_sv2v_reg;
  assign mem[1833] = mem_1833_sv2v_reg;
  assign mem[1832] = mem_1832_sv2v_reg;
  assign mem[1831] = mem_1831_sv2v_reg;
  assign mem[1830] = mem_1830_sv2v_reg;
  assign mem[1829] = mem_1829_sv2v_reg;
  assign mem[1828] = mem_1828_sv2v_reg;
  assign mem[1827] = mem_1827_sv2v_reg;
  assign mem[1826] = mem_1826_sv2v_reg;
  assign mem[1825] = mem_1825_sv2v_reg;
  assign mem[1824] = mem_1824_sv2v_reg;
  assign mem[1823] = mem_1823_sv2v_reg;
  assign mem[1822] = mem_1822_sv2v_reg;
  assign mem[1821] = mem_1821_sv2v_reg;
  assign mem[1820] = mem_1820_sv2v_reg;
  assign mem[1819] = mem_1819_sv2v_reg;
  assign mem[1818] = mem_1818_sv2v_reg;
  assign mem[1817] = mem_1817_sv2v_reg;
  assign mem[1816] = mem_1816_sv2v_reg;
  assign mem[1815] = mem_1815_sv2v_reg;
  assign mem[1814] = mem_1814_sv2v_reg;
  assign mem[1813] = mem_1813_sv2v_reg;
  assign mem[1812] = mem_1812_sv2v_reg;
  assign mem[1811] = mem_1811_sv2v_reg;
  assign mem[1810] = mem_1810_sv2v_reg;
  assign mem[1809] = mem_1809_sv2v_reg;
  assign mem[1808] = mem_1808_sv2v_reg;
  assign mem[1807] = mem_1807_sv2v_reg;
  assign mem[1806] = mem_1806_sv2v_reg;
  assign mem[1805] = mem_1805_sv2v_reg;
  assign mem[1804] = mem_1804_sv2v_reg;
  assign mem[1803] = mem_1803_sv2v_reg;
  assign mem[1802] = mem_1802_sv2v_reg;
  assign mem[1801] = mem_1801_sv2v_reg;
  assign mem[1800] = mem_1800_sv2v_reg;
  assign mem[1799] = mem_1799_sv2v_reg;
  assign mem[1798] = mem_1798_sv2v_reg;
  assign mem[1797] = mem_1797_sv2v_reg;
  assign mem[1796] = mem_1796_sv2v_reg;
  assign mem[1795] = mem_1795_sv2v_reg;
  assign mem[1794] = mem_1794_sv2v_reg;
  assign mem[1793] = mem_1793_sv2v_reg;
  assign mem[1792] = mem_1792_sv2v_reg;
  assign mem[1791] = mem_1791_sv2v_reg;
  assign mem[1790] = mem_1790_sv2v_reg;
  assign mem[1789] = mem_1789_sv2v_reg;
  assign mem[1788] = mem_1788_sv2v_reg;
  assign mem[1787] = mem_1787_sv2v_reg;
  assign mem[1786] = mem_1786_sv2v_reg;
  assign mem[1785] = mem_1785_sv2v_reg;
  assign mem[1784] = mem_1784_sv2v_reg;
  assign mem[1783] = mem_1783_sv2v_reg;
  assign mem[1782] = mem_1782_sv2v_reg;
  assign mem[1781] = mem_1781_sv2v_reg;
  assign mem[1780] = mem_1780_sv2v_reg;
  assign mem[1779] = mem_1779_sv2v_reg;
  assign mem[1778] = mem_1778_sv2v_reg;
  assign mem[1777] = mem_1777_sv2v_reg;
  assign mem[1776] = mem_1776_sv2v_reg;
  assign mem[1775] = mem_1775_sv2v_reg;
  assign mem[1774] = mem_1774_sv2v_reg;
  assign mem[1773] = mem_1773_sv2v_reg;
  assign mem[1772] = mem_1772_sv2v_reg;
  assign mem[1771] = mem_1771_sv2v_reg;
  assign mem[1770] = mem_1770_sv2v_reg;
  assign mem[1769] = mem_1769_sv2v_reg;
  assign mem[1768] = mem_1768_sv2v_reg;
  assign mem[1767] = mem_1767_sv2v_reg;
  assign mem[1766] = mem_1766_sv2v_reg;
  assign mem[1765] = mem_1765_sv2v_reg;
  assign mem[1764] = mem_1764_sv2v_reg;
  assign mem[1763] = mem_1763_sv2v_reg;
  assign mem[1762] = mem_1762_sv2v_reg;
  assign mem[1761] = mem_1761_sv2v_reg;
  assign mem[1760] = mem_1760_sv2v_reg;
  assign mem[1759] = mem_1759_sv2v_reg;
  assign mem[1758] = mem_1758_sv2v_reg;
  assign mem[1757] = mem_1757_sv2v_reg;
  assign mem[1756] = mem_1756_sv2v_reg;
  assign mem[1755] = mem_1755_sv2v_reg;
  assign mem[1754] = mem_1754_sv2v_reg;
  assign mem[1753] = mem_1753_sv2v_reg;
  assign mem[1752] = mem_1752_sv2v_reg;
  assign mem[1751] = mem_1751_sv2v_reg;
  assign mem[1750] = mem_1750_sv2v_reg;
  assign mem[1749] = mem_1749_sv2v_reg;
  assign mem[1748] = mem_1748_sv2v_reg;
  assign mem[1747] = mem_1747_sv2v_reg;
  assign mem[1746] = mem_1746_sv2v_reg;
  assign mem[1745] = mem_1745_sv2v_reg;
  assign mem[1744] = mem_1744_sv2v_reg;
  assign mem[1743] = mem_1743_sv2v_reg;
  assign mem[1742] = mem_1742_sv2v_reg;
  assign mem[1741] = mem_1741_sv2v_reg;
  assign mem[1740] = mem_1740_sv2v_reg;
  assign mem[1739] = mem_1739_sv2v_reg;
  assign mem[1738] = mem_1738_sv2v_reg;
  assign mem[1737] = mem_1737_sv2v_reg;
  assign mem[1736] = mem_1736_sv2v_reg;
  assign mem[1735] = mem_1735_sv2v_reg;
  assign mem[1734] = mem_1734_sv2v_reg;
  assign mem[1733] = mem_1733_sv2v_reg;
  assign mem[1732] = mem_1732_sv2v_reg;
  assign mem[1731] = mem_1731_sv2v_reg;
  assign mem[1730] = mem_1730_sv2v_reg;
  assign mem[1729] = mem_1729_sv2v_reg;
  assign mem[1728] = mem_1728_sv2v_reg;
  assign mem[1727] = mem_1727_sv2v_reg;
  assign mem[1726] = mem_1726_sv2v_reg;
  assign mem[1725] = mem_1725_sv2v_reg;
  assign mem[1724] = mem_1724_sv2v_reg;
  assign mem[1723] = mem_1723_sv2v_reg;
  assign mem[1722] = mem_1722_sv2v_reg;
  assign mem[1721] = mem_1721_sv2v_reg;
  assign mem[1720] = mem_1720_sv2v_reg;
  assign mem[1719] = mem_1719_sv2v_reg;
  assign mem[1718] = mem_1718_sv2v_reg;
  assign mem[1717] = mem_1717_sv2v_reg;
  assign mem[1716] = mem_1716_sv2v_reg;
  assign mem[1715] = mem_1715_sv2v_reg;
  assign mem[1714] = mem_1714_sv2v_reg;
  assign mem[1713] = mem_1713_sv2v_reg;
  assign mem[1712] = mem_1712_sv2v_reg;
  assign mem[1711] = mem_1711_sv2v_reg;
  assign mem[1710] = mem_1710_sv2v_reg;
  assign mem[1709] = mem_1709_sv2v_reg;
  assign mem[1708] = mem_1708_sv2v_reg;
  assign mem[1707] = mem_1707_sv2v_reg;
  assign mem[1706] = mem_1706_sv2v_reg;
  assign mem[1705] = mem_1705_sv2v_reg;
  assign mem[1704] = mem_1704_sv2v_reg;
  assign mem[1703] = mem_1703_sv2v_reg;
  assign mem[1702] = mem_1702_sv2v_reg;
  assign mem[1701] = mem_1701_sv2v_reg;
  assign mem[1700] = mem_1700_sv2v_reg;
  assign mem[1699] = mem_1699_sv2v_reg;
  assign mem[1698] = mem_1698_sv2v_reg;
  assign mem[1697] = mem_1697_sv2v_reg;
  assign mem[1696] = mem_1696_sv2v_reg;
  assign mem[1695] = mem_1695_sv2v_reg;
  assign mem[1694] = mem_1694_sv2v_reg;
  assign mem[1693] = mem_1693_sv2v_reg;
  assign mem[1692] = mem_1692_sv2v_reg;
  assign mem[1691] = mem_1691_sv2v_reg;
  assign mem[1690] = mem_1690_sv2v_reg;
  assign mem[1689] = mem_1689_sv2v_reg;
  assign mem[1688] = mem_1688_sv2v_reg;
  assign mem[1687] = mem_1687_sv2v_reg;
  assign mem[1686] = mem_1686_sv2v_reg;
  assign mem[1685] = mem_1685_sv2v_reg;
  assign mem[1684] = mem_1684_sv2v_reg;
  assign mem[1683] = mem_1683_sv2v_reg;
  assign mem[1682] = mem_1682_sv2v_reg;
  assign mem[1681] = mem_1681_sv2v_reg;
  assign mem[1680] = mem_1680_sv2v_reg;
  assign mem[1679] = mem_1679_sv2v_reg;
  assign mem[1678] = mem_1678_sv2v_reg;
  assign mem[1677] = mem_1677_sv2v_reg;
  assign mem[1676] = mem_1676_sv2v_reg;
  assign mem[1675] = mem_1675_sv2v_reg;
  assign mem[1674] = mem_1674_sv2v_reg;
  assign mem[1673] = mem_1673_sv2v_reg;
  assign mem[1672] = mem_1672_sv2v_reg;
  assign mem[1671] = mem_1671_sv2v_reg;
  assign mem[1670] = mem_1670_sv2v_reg;
  assign mem[1669] = mem_1669_sv2v_reg;
  assign mem[1668] = mem_1668_sv2v_reg;
  assign mem[1667] = mem_1667_sv2v_reg;
  assign mem[1666] = mem_1666_sv2v_reg;
  assign mem[1665] = mem_1665_sv2v_reg;
  assign mem[1664] = mem_1664_sv2v_reg;
  assign mem[1663] = mem_1663_sv2v_reg;
  assign mem[1662] = mem_1662_sv2v_reg;
  assign mem[1661] = mem_1661_sv2v_reg;
  assign mem[1660] = mem_1660_sv2v_reg;
  assign mem[1659] = mem_1659_sv2v_reg;
  assign mem[1658] = mem_1658_sv2v_reg;
  assign mem[1657] = mem_1657_sv2v_reg;
  assign mem[1656] = mem_1656_sv2v_reg;
  assign mem[1655] = mem_1655_sv2v_reg;
  assign mem[1654] = mem_1654_sv2v_reg;
  assign mem[1653] = mem_1653_sv2v_reg;
  assign mem[1652] = mem_1652_sv2v_reg;
  assign mem[1651] = mem_1651_sv2v_reg;
  assign mem[1650] = mem_1650_sv2v_reg;
  assign mem[1649] = mem_1649_sv2v_reg;
  assign mem[1648] = mem_1648_sv2v_reg;
  assign mem[1647] = mem_1647_sv2v_reg;
  assign mem[1646] = mem_1646_sv2v_reg;
  assign mem[1645] = mem_1645_sv2v_reg;
  assign mem[1644] = mem_1644_sv2v_reg;
  assign mem[1643] = mem_1643_sv2v_reg;
  assign mem[1642] = mem_1642_sv2v_reg;
  assign mem[1641] = mem_1641_sv2v_reg;
  assign mem[1640] = mem_1640_sv2v_reg;
  assign mem[1639] = mem_1639_sv2v_reg;
  assign mem[1638] = mem_1638_sv2v_reg;
  assign mem[1637] = mem_1637_sv2v_reg;
  assign mem[1636] = mem_1636_sv2v_reg;
  assign mem[1635] = mem_1635_sv2v_reg;
  assign mem[1634] = mem_1634_sv2v_reg;
  assign mem[1633] = mem_1633_sv2v_reg;
  assign mem[1632] = mem_1632_sv2v_reg;
  assign mem[1631] = mem_1631_sv2v_reg;
  assign mem[1630] = mem_1630_sv2v_reg;
  assign mem[1629] = mem_1629_sv2v_reg;
  assign mem[1628] = mem_1628_sv2v_reg;
  assign mem[1627] = mem_1627_sv2v_reg;
  assign mem[1626] = mem_1626_sv2v_reg;
  assign mem[1625] = mem_1625_sv2v_reg;
  assign mem[1624] = mem_1624_sv2v_reg;
  assign mem[1623] = mem_1623_sv2v_reg;
  assign mem[1622] = mem_1622_sv2v_reg;
  assign mem[1621] = mem_1621_sv2v_reg;
  assign mem[1620] = mem_1620_sv2v_reg;
  assign mem[1619] = mem_1619_sv2v_reg;
  assign mem[1618] = mem_1618_sv2v_reg;
  assign mem[1617] = mem_1617_sv2v_reg;
  assign mem[1616] = mem_1616_sv2v_reg;
  assign mem[1615] = mem_1615_sv2v_reg;
  assign mem[1614] = mem_1614_sv2v_reg;
  assign mem[1613] = mem_1613_sv2v_reg;
  assign mem[1612] = mem_1612_sv2v_reg;
  assign mem[1611] = mem_1611_sv2v_reg;
  assign mem[1610] = mem_1610_sv2v_reg;
  assign mem[1609] = mem_1609_sv2v_reg;
  assign mem[1608] = mem_1608_sv2v_reg;
  assign mem[1607] = mem_1607_sv2v_reg;
  assign mem[1606] = mem_1606_sv2v_reg;
  assign mem[1605] = mem_1605_sv2v_reg;
  assign mem[1604] = mem_1604_sv2v_reg;
  assign mem[1603] = mem_1603_sv2v_reg;
  assign mem[1602] = mem_1602_sv2v_reg;
  assign mem[1601] = mem_1601_sv2v_reg;
  assign mem[1600] = mem_1600_sv2v_reg;
  assign mem[1599] = mem_1599_sv2v_reg;
  assign mem[1598] = mem_1598_sv2v_reg;
  assign mem[1597] = mem_1597_sv2v_reg;
  assign mem[1596] = mem_1596_sv2v_reg;
  assign mem[1595] = mem_1595_sv2v_reg;
  assign mem[1594] = mem_1594_sv2v_reg;
  assign mem[1593] = mem_1593_sv2v_reg;
  assign mem[1592] = mem_1592_sv2v_reg;
  assign mem[1591] = mem_1591_sv2v_reg;
  assign mem[1590] = mem_1590_sv2v_reg;
  assign mem[1589] = mem_1589_sv2v_reg;
  assign mem[1588] = mem_1588_sv2v_reg;
  assign mem[1587] = mem_1587_sv2v_reg;
  assign mem[1586] = mem_1586_sv2v_reg;
  assign mem[1585] = mem_1585_sv2v_reg;
  assign mem[1584] = mem_1584_sv2v_reg;
  assign mem[1583] = mem_1583_sv2v_reg;
  assign mem[1582] = mem_1582_sv2v_reg;
  assign mem[1581] = mem_1581_sv2v_reg;
  assign mem[1580] = mem_1580_sv2v_reg;
  assign mem[1579] = mem_1579_sv2v_reg;
  assign mem[1578] = mem_1578_sv2v_reg;
  assign mem[1577] = mem_1577_sv2v_reg;
  assign mem[1576] = mem_1576_sv2v_reg;
  assign mem[1575] = mem_1575_sv2v_reg;
  assign mem[1574] = mem_1574_sv2v_reg;
  assign mem[1573] = mem_1573_sv2v_reg;
  assign mem[1572] = mem_1572_sv2v_reg;
  assign mem[1571] = mem_1571_sv2v_reg;
  assign mem[1570] = mem_1570_sv2v_reg;
  assign mem[1569] = mem_1569_sv2v_reg;
  assign mem[1568] = mem_1568_sv2v_reg;
  assign mem[1567] = mem_1567_sv2v_reg;
  assign mem[1566] = mem_1566_sv2v_reg;
  assign mem[1565] = mem_1565_sv2v_reg;
  assign mem[1564] = mem_1564_sv2v_reg;
  assign mem[1563] = mem_1563_sv2v_reg;
  assign mem[1562] = mem_1562_sv2v_reg;
  assign mem[1561] = mem_1561_sv2v_reg;
  assign mem[1560] = mem_1560_sv2v_reg;
  assign mem[1559] = mem_1559_sv2v_reg;
  assign mem[1558] = mem_1558_sv2v_reg;
  assign mem[1557] = mem_1557_sv2v_reg;
  assign mem[1556] = mem_1556_sv2v_reg;
  assign mem[1555] = mem_1555_sv2v_reg;
  assign mem[1554] = mem_1554_sv2v_reg;
  assign mem[1553] = mem_1553_sv2v_reg;
  assign mem[1552] = mem_1552_sv2v_reg;
  assign mem[1551] = mem_1551_sv2v_reg;
  assign mem[1550] = mem_1550_sv2v_reg;
  assign mem[1549] = mem_1549_sv2v_reg;
  assign mem[1548] = mem_1548_sv2v_reg;
  assign mem[1547] = mem_1547_sv2v_reg;
  assign mem[1546] = mem_1546_sv2v_reg;
  assign mem[1545] = mem_1545_sv2v_reg;
  assign mem[1544] = mem_1544_sv2v_reg;
  assign mem[1543] = mem_1543_sv2v_reg;
  assign mem[1542] = mem_1542_sv2v_reg;
  assign mem[1541] = mem_1541_sv2v_reg;
  assign mem[1540] = mem_1540_sv2v_reg;
  assign mem[1539] = mem_1539_sv2v_reg;
  assign mem[1538] = mem_1538_sv2v_reg;
  assign mem[1537] = mem_1537_sv2v_reg;
  assign mem[1536] = mem_1536_sv2v_reg;
  assign mem[1535] = mem_1535_sv2v_reg;
  assign mem[1534] = mem_1534_sv2v_reg;
  assign mem[1533] = mem_1533_sv2v_reg;
  assign mem[1532] = mem_1532_sv2v_reg;
  assign mem[1531] = mem_1531_sv2v_reg;
  assign mem[1530] = mem_1530_sv2v_reg;
  assign mem[1529] = mem_1529_sv2v_reg;
  assign mem[1528] = mem_1528_sv2v_reg;
  assign mem[1527] = mem_1527_sv2v_reg;
  assign mem[1526] = mem_1526_sv2v_reg;
  assign mem[1525] = mem_1525_sv2v_reg;
  assign mem[1524] = mem_1524_sv2v_reg;
  assign mem[1523] = mem_1523_sv2v_reg;
  assign mem[1522] = mem_1522_sv2v_reg;
  assign mem[1521] = mem_1521_sv2v_reg;
  assign mem[1520] = mem_1520_sv2v_reg;
  assign mem[1519] = mem_1519_sv2v_reg;
  assign mem[1518] = mem_1518_sv2v_reg;
  assign mem[1517] = mem_1517_sv2v_reg;
  assign mem[1516] = mem_1516_sv2v_reg;
  assign mem[1515] = mem_1515_sv2v_reg;
  assign mem[1514] = mem_1514_sv2v_reg;
  assign mem[1513] = mem_1513_sv2v_reg;
  assign mem[1512] = mem_1512_sv2v_reg;
  assign mem[1511] = mem_1511_sv2v_reg;
  assign mem[1510] = mem_1510_sv2v_reg;
  assign mem[1509] = mem_1509_sv2v_reg;
  assign mem[1508] = mem_1508_sv2v_reg;
  assign mem[1507] = mem_1507_sv2v_reg;
  assign mem[1506] = mem_1506_sv2v_reg;
  assign mem[1505] = mem_1505_sv2v_reg;
  assign mem[1504] = mem_1504_sv2v_reg;
  assign mem[1503] = mem_1503_sv2v_reg;
  assign mem[1502] = mem_1502_sv2v_reg;
  assign mem[1501] = mem_1501_sv2v_reg;
  assign mem[1500] = mem_1500_sv2v_reg;
  assign mem[1499] = mem_1499_sv2v_reg;
  assign mem[1498] = mem_1498_sv2v_reg;
  assign mem[1497] = mem_1497_sv2v_reg;
  assign mem[1496] = mem_1496_sv2v_reg;
  assign mem[1495] = mem_1495_sv2v_reg;
  assign mem[1494] = mem_1494_sv2v_reg;
  assign mem[1493] = mem_1493_sv2v_reg;
  assign mem[1492] = mem_1492_sv2v_reg;
  assign mem[1491] = mem_1491_sv2v_reg;
  assign mem[1490] = mem_1490_sv2v_reg;
  assign mem[1489] = mem_1489_sv2v_reg;
  assign mem[1488] = mem_1488_sv2v_reg;
  assign mem[1487] = mem_1487_sv2v_reg;
  assign mem[1486] = mem_1486_sv2v_reg;
  assign mem[1485] = mem_1485_sv2v_reg;
  assign mem[1484] = mem_1484_sv2v_reg;
  assign mem[1483] = mem_1483_sv2v_reg;
  assign mem[1482] = mem_1482_sv2v_reg;
  assign mem[1481] = mem_1481_sv2v_reg;
  assign mem[1480] = mem_1480_sv2v_reg;
  assign mem[1479] = mem_1479_sv2v_reg;
  assign mem[1478] = mem_1478_sv2v_reg;
  assign mem[1477] = mem_1477_sv2v_reg;
  assign mem[1476] = mem_1476_sv2v_reg;
  assign mem[1475] = mem_1475_sv2v_reg;
  assign mem[1474] = mem_1474_sv2v_reg;
  assign mem[1473] = mem_1473_sv2v_reg;
  assign mem[1472] = mem_1472_sv2v_reg;
  assign mem[1471] = mem_1471_sv2v_reg;
  assign mem[1470] = mem_1470_sv2v_reg;
  assign mem[1469] = mem_1469_sv2v_reg;
  assign mem[1468] = mem_1468_sv2v_reg;
  assign mem[1467] = mem_1467_sv2v_reg;
  assign mem[1466] = mem_1466_sv2v_reg;
  assign mem[1465] = mem_1465_sv2v_reg;
  assign mem[1464] = mem_1464_sv2v_reg;
  assign mem[1463] = mem_1463_sv2v_reg;
  assign mem[1462] = mem_1462_sv2v_reg;
  assign mem[1461] = mem_1461_sv2v_reg;
  assign mem[1460] = mem_1460_sv2v_reg;
  assign mem[1459] = mem_1459_sv2v_reg;
  assign mem[1458] = mem_1458_sv2v_reg;
  assign mem[1457] = mem_1457_sv2v_reg;
  assign mem[1456] = mem_1456_sv2v_reg;
  assign mem[1455] = mem_1455_sv2v_reg;
  assign mem[1454] = mem_1454_sv2v_reg;
  assign mem[1453] = mem_1453_sv2v_reg;
  assign mem[1452] = mem_1452_sv2v_reg;
  assign mem[1451] = mem_1451_sv2v_reg;
  assign mem[1450] = mem_1450_sv2v_reg;
  assign mem[1449] = mem_1449_sv2v_reg;
  assign mem[1448] = mem_1448_sv2v_reg;
  assign mem[1447] = mem_1447_sv2v_reg;
  assign mem[1446] = mem_1446_sv2v_reg;
  assign mem[1445] = mem_1445_sv2v_reg;
  assign mem[1444] = mem_1444_sv2v_reg;
  assign mem[1443] = mem_1443_sv2v_reg;
  assign mem[1442] = mem_1442_sv2v_reg;
  assign mem[1441] = mem_1441_sv2v_reg;
  assign mem[1440] = mem_1440_sv2v_reg;
  assign mem[1439] = mem_1439_sv2v_reg;
  assign mem[1438] = mem_1438_sv2v_reg;
  assign mem[1437] = mem_1437_sv2v_reg;
  assign mem[1436] = mem_1436_sv2v_reg;
  assign mem[1435] = mem_1435_sv2v_reg;
  assign mem[1434] = mem_1434_sv2v_reg;
  assign mem[1433] = mem_1433_sv2v_reg;
  assign mem[1432] = mem_1432_sv2v_reg;
  assign mem[1431] = mem_1431_sv2v_reg;
  assign mem[1430] = mem_1430_sv2v_reg;
  assign mem[1429] = mem_1429_sv2v_reg;
  assign mem[1428] = mem_1428_sv2v_reg;
  assign mem[1427] = mem_1427_sv2v_reg;
  assign mem[1426] = mem_1426_sv2v_reg;
  assign mem[1425] = mem_1425_sv2v_reg;
  assign mem[1424] = mem_1424_sv2v_reg;
  assign mem[1423] = mem_1423_sv2v_reg;
  assign mem[1422] = mem_1422_sv2v_reg;
  assign mem[1421] = mem_1421_sv2v_reg;
  assign mem[1420] = mem_1420_sv2v_reg;
  assign mem[1419] = mem_1419_sv2v_reg;
  assign mem[1418] = mem_1418_sv2v_reg;
  assign mem[1417] = mem_1417_sv2v_reg;
  assign mem[1416] = mem_1416_sv2v_reg;
  assign mem[1415] = mem_1415_sv2v_reg;
  assign mem[1414] = mem_1414_sv2v_reg;
  assign mem[1413] = mem_1413_sv2v_reg;
  assign mem[1412] = mem_1412_sv2v_reg;
  assign mem[1411] = mem_1411_sv2v_reg;
  assign mem[1410] = mem_1410_sv2v_reg;
  assign mem[1409] = mem_1409_sv2v_reg;
  assign mem[1408] = mem_1408_sv2v_reg;
  assign mem[1407] = mem_1407_sv2v_reg;
  assign mem[1406] = mem_1406_sv2v_reg;
  assign mem[1405] = mem_1405_sv2v_reg;
  assign mem[1404] = mem_1404_sv2v_reg;
  assign mem[1403] = mem_1403_sv2v_reg;
  assign mem[1402] = mem_1402_sv2v_reg;
  assign mem[1401] = mem_1401_sv2v_reg;
  assign mem[1400] = mem_1400_sv2v_reg;
  assign mem[1399] = mem_1399_sv2v_reg;
  assign mem[1398] = mem_1398_sv2v_reg;
  assign mem[1397] = mem_1397_sv2v_reg;
  assign mem[1396] = mem_1396_sv2v_reg;
  assign mem[1395] = mem_1395_sv2v_reg;
  assign mem[1394] = mem_1394_sv2v_reg;
  assign mem[1393] = mem_1393_sv2v_reg;
  assign mem[1392] = mem_1392_sv2v_reg;
  assign mem[1391] = mem_1391_sv2v_reg;
  assign mem[1390] = mem_1390_sv2v_reg;
  assign mem[1389] = mem_1389_sv2v_reg;
  assign mem[1388] = mem_1388_sv2v_reg;
  assign mem[1387] = mem_1387_sv2v_reg;
  assign mem[1386] = mem_1386_sv2v_reg;
  assign mem[1385] = mem_1385_sv2v_reg;
  assign mem[1384] = mem_1384_sv2v_reg;
  assign mem[1383] = mem_1383_sv2v_reg;
  assign mem[1382] = mem_1382_sv2v_reg;
  assign mem[1381] = mem_1381_sv2v_reg;
  assign mem[1380] = mem_1380_sv2v_reg;
  assign mem[1379] = mem_1379_sv2v_reg;
  assign mem[1378] = mem_1378_sv2v_reg;
  assign mem[1377] = mem_1377_sv2v_reg;
  assign mem[1376] = mem_1376_sv2v_reg;
  assign mem[1375] = mem_1375_sv2v_reg;
  assign mem[1374] = mem_1374_sv2v_reg;
  assign mem[1373] = mem_1373_sv2v_reg;
  assign mem[1372] = mem_1372_sv2v_reg;
  assign mem[1371] = mem_1371_sv2v_reg;
  assign mem[1370] = mem_1370_sv2v_reg;
  assign mem[1369] = mem_1369_sv2v_reg;
  assign mem[1368] = mem_1368_sv2v_reg;
  assign mem[1367] = mem_1367_sv2v_reg;
  assign mem[1366] = mem_1366_sv2v_reg;
  assign mem[1365] = mem_1365_sv2v_reg;
  assign mem[1364] = mem_1364_sv2v_reg;
  assign mem[1363] = mem_1363_sv2v_reg;
  assign mem[1362] = mem_1362_sv2v_reg;
  assign mem[1361] = mem_1361_sv2v_reg;
  assign mem[1360] = mem_1360_sv2v_reg;
  assign mem[1359] = mem_1359_sv2v_reg;
  assign mem[1358] = mem_1358_sv2v_reg;
  assign mem[1357] = mem_1357_sv2v_reg;
  assign mem[1356] = mem_1356_sv2v_reg;
  assign mem[1355] = mem_1355_sv2v_reg;
  assign mem[1354] = mem_1354_sv2v_reg;
  assign mem[1353] = mem_1353_sv2v_reg;
  assign mem[1352] = mem_1352_sv2v_reg;
  assign mem[1351] = mem_1351_sv2v_reg;
  assign mem[1350] = mem_1350_sv2v_reg;
  assign mem[1349] = mem_1349_sv2v_reg;
  assign mem[1348] = mem_1348_sv2v_reg;
  assign mem[1347] = mem_1347_sv2v_reg;
  assign mem[1346] = mem_1346_sv2v_reg;
  assign mem[1345] = mem_1345_sv2v_reg;
  assign mem[1344] = mem_1344_sv2v_reg;
  assign mem[1343] = mem_1343_sv2v_reg;
  assign mem[1342] = mem_1342_sv2v_reg;
  assign mem[1341] = mem_1341_sv2v_reg;
  assign mem[1340] = mem_1340_sv2v_reg;
  assign mem[1339] = mem_1339_sv2v_reg;
  assign mem[1338] = mem_1338_sv2v_reg;
  assign mem[1337] = mem_1337_sv2v_reg;
  assign mem[1336] = mem_1336_sv2v_reg;
  assign mem[1335] = mem_1335_sv2v_reg;
  assign mem[1334] = mem_1334_sv2v_reg;
  assign mem[1333] = mem_1333_sv2v_reg;
  assign mem[1332] = mem_1332_sv2v_reg;
  assign mem[1331] = mem_1331_sv2v_reg;
  assign mem[1330] = mem_1330_sv2v_reg;
  assign mem[1329] = mem_1329_sv2v_reg;
  assign mem[1328] = mem_1328_sv2v_reg;
  assign mem[1327] = mem_1327_sv2v_reg;
  assign mem[1326] = mem_1326_sv2v_reg;
  assign mem[1325] = mem_1325_sv2v_reg;
  assign mem[1324] = mem_1324_sv2v_reg;
  assign mem[1323] = mem_1323_sv2v_reg;
  assign mem[1322] = mem_1322_sv2v_reg;
  assign mem[1321] = mem_1321_sv2v_reg;
  assign mem[1320] = mem_1320_sv2v_reg;
  assign mem[1319] = mem_1319_sv2v_reg;
  assign mem[1318] = mem_1318_sv2v_reg;
  assign mem[1317] = mem_1317_sv2v_reg;
  assign mem[1316] = mem_1316_sv2v_reg;
  assign mem[1315] = mem_1315_sv2v_reg;
  assign mem[1314] = mem_1314_sv2v_reg;
  assign mem[1313] = mem_1313_sv2v_reg;
  assign mem[1312] = mem_1312_sv2v_reg;
  assign mem[1311] = mem_1311_sv2v_reg;
  assign mem[1310] = mem_1310_sv2v_reg;
  assign mem[1309] = mem_1309_sv2v_reg;
  assign mem[1308] = mem_1308_sv2v_reg;
  assign mem[1307] = mem_1307_sv2v_reg;
  assign mem[1306] = mem_1306_sv2v_reg;
  assign mem[1305] = mem_1305_sv2v_reg;
  assign mem[1304] = mem_1304_sv2v_reg;
  assign mem[1303] = mem_1303_sv2v_reg;
  assign mem[1302] = mem_1302_sv2v_reg;
  assign mem[1301] = mem_1301_sv2v_reg;
  assign mem[1300] = mem_1300_sv2v_reg;
  assign mem[1299] = mem_1299_sv2v_reg;
  assign mem[1298] = mem_1298_sv2v_reg;
  assign mem[1297] = mem_1297_sv2v_reg;
  assign mem[1296] = mem_1296_sv2v_reg;
  assign mem[1295] = mem_1295_sv2v_reg;
  assign mem[1294] = mem_1294_sv2v_reg;
  assign mem[1293] = mem_1293_sv2v_reg;
  assign mem[1292] = mem_1292_sv2v_reg;
  assign mem[1291] = mem_1291_sv2v_reg;
  assign mem[1290] = mem_1290_sv2v_reg;
  assign mem[1289] = mem_1289_sv2v_reg;
  assign mem[1288] = mem_1288_sv2v_reg;
  assign mem[1287] = mem_1287_sv2v_reg;
  assign mem[1286] = mem_1286_sv2v_reg;
  assign mem[1285] = mem_1285_sv2v_reg;
  assign mem[1284] = mem_1284_sv2v_reg;
  assign mem[1283] = mem_1283_sv2v_reg;
  assign mem[1282] = mem_1282_sv2v_reg;
  assign mem[1281] = mem_1281_sv2v_reg;
  assign mem[1280] = mem_1280_sv2v_reg;
  assign mem[1279] = mem_1279_sv2v_reg;
  assign mem[1278] = mem_1278_sv2v_reg;
  assign mem[1277] = mem_1277_sv2v_reg;
  assign mem[1276] = mem_1276_sv2v_reg;
  assign mem[1275] = mem_1275_sv2v_reg;
  assign mem[1274] = mem_1274_sv2v_reg;
  assign mem[1273] = mem_1273_sv2v_reg;
  assign mem[1272] = mem_1272_sv2v_reg;
  assign mem[1271] = mem_1271_sv2v_reg;
  assign mem[1270] = mem_1270_sv2v_reg;
  assign mem[1269] = mem_1269_sv2v_reg;
  assign mem[1268] = mem_1268_sv2v_reg;
  assign mem[1267] = mem_1267_sv2v_reg;
  assign mem[1266] = mem_1266_sv2v_reg;
  assign mem[1265] = mem_1265_sv2v_reg;
  assign mem[1264] = mem_1264_sv2v_reg;
  assign mem[1263] = mem_1263_sv2v_reg;
  assign mem[1262] = mem_1262_sv2v_reg;
  assign mem[1261] = mem_1261_sv2v_reg;
  assign mem[1260] = mem_1260_sv2v_reg;
  assign mem[1259] = mem_1259_sv2v_reg;
  assign mem[1258] = mem_1258_sv2v_reg;
  assign mem[1257] = mem_1257_sv2v_reg;
  assign mem[1256] = mem_1256_sv2v_reg;
  assign mem[1255] = mem_1255_sv2v_reg;
  assign mem[1254] = mem_1254_sv2v_reg;
  assign mem[1253] = mem_1253_sv2v_reg;
  assign mem[1252] = mem_1252_sv2v_reg;
  assign mem[1251] = mem_1251_sv2v_reg;
  assign mem[1250] = mem_1250_sv2v_reg;
  assign mem[1249] = mem_1249_sv2v_reg;
  assign mem[1248] = mem_1248_sv2v_reg;
  assign mem[1247] = mem_1247_sv2v_reg;
  assign mem[1246] = mem_1246_sv2v_reg;
  assign mem[1245] = mem_1245_sv2v_reg;
  assign mem[1244] = mem_1244_sv2v_reg;
  assign mem[1243] = mem_1243_sv2v_reg;
  assign mem[1242] = mem_1242_sv2v_reg;
  assign mem[1241] = mem_1241_sv2v_reg;
  assign mem[1240] = mem_1240_sv2v_reg;
  assign mem[1239] = mem_1239_sv2v_reg;
  assign mem[1238] = mem_1238_sv2v_reg;
  assign mem[1237] = mem_1237_sv2v_reg;
  assign mem[1236] = mem_1236_sv2v_reg;
  assign mem[1235] = mem_1235_sv2v_reg;
  assign mem[1234] = mem_1234_sv2v_reg;
  assign mem[1233] = mem_1233_sv2v_reg;
  assign mem[1232] = mem_1232_sv2v_reg;
  assign mem[1231] = mem_1231_sv2v_reg;
  assign mem[1230] = mem_1230_sv2v_reg;
  assign mem[1229] = mem_1229_sv2v_reg;
  assign mem[1228] = mem_1228_sv2v_reg;
  assign mem[1227] = mem_1227_sv2v_reg;
  assign mem[1226] = mem_1226_sv2v_reg;
  assign mem[1225] = mem_1225_sv2v_reg;
  assign mem[1224] = mem_1224_sv2v_reg;
  assign mem[1223] = mem_1223_sv2v_reg;
  assign mem[1222] = mem_1222_sv2v_reg;
  assign mem[1221] = mem_1221_sv2v_reg;
  assign mem[1220] = mem_1220_sv2v_reg;
  assign mem[1219] = mem_1219_sv2v_reg;
  assign mem[1218] = mem_1218_sv2v_reg;
  assign mem[1217] = mem_1217_sv2v_reg;
  assign mem[1216] = mem_1216_sv2v_reg;
  assign mem[1215] = mem_1215_sv2v_reg;
  assign mem[1214] = mem_1214_sv2v_reg;
  assign mem[1213] = mem_1213_sv2v_reg;
  assign mem[1212] = mem_1212_sv2v_reg;
  assign mem[1211] = mem_1211_sv2v_reg;
  assign mem[1210] = mem_1210_sv2v_reg;
  assign mem[1209] = mem_1209_sv2v_reg;
  assign mem[1208] = mem_1208_sv2v_reg;
  assign mem[1207] = mem_1207_sv2v_reg;
  assign mem[1206] = mem_1206_sv2v_reg;
  assign mem[1205] = mem_1205_sv2v_reg;
  assign mem[1204] = mem_1204_sv2v_reg;
  assign mem[1203] = mem_1203_sv2v_reg;
  assign mem[1202] = mem_1202_sv2v_reg;
  assign mem[1201] = mem_1201_sv2v_reg;
  assign mem[1200] = mem_1200_sv2v_reg;
  assign mem[1199] = mem_1199_sv2v_reg;
  assign mem[1198] = mem_1198_sv2v_reg;
  assign mem[1197] = mem_1197_sv2v_reg;
  assign mem[1196] = mem_1196_sv2v_reg;
  assign mem[1195] = mem_1195_sv2v_reg;
  assign mem[1194] = mem_1194_sv2v_reg;
  assign mem[1193] = mem_1193_sv2v_reg;
  assign mem[1192] = mem_1192_sv2v_reg;
  assign mem[1191] = mem_1191_sv2v_reg;
  assign mem[1190] = mem_1190_sv2v_reg;
  assign mem[1189] = mem_1189_sv2v_reg;
  assign mem[1188] = mem_1188_sv2v_reg;
  assign mem[1187] = mem_1187_sv2v_reg;
  assign mem[1186] = mem_1186_sv2v_reg;
  assign mem[1185] = mem_1185_sv2v_reg;
  assign mem[1184] = mem_1184_sv2v_reg;
  assign mem[1183] = mem_1183_sv2v_reg;
  assign mem[1182] = mem_1182_sv2v_reg;
  assign mem[1181] = mem_1181_sv2v_reg;
  assign mem[1180] = mem_1180_sv2v_reg;
  assign mem[1179] = mem_1179_sv2v_reg;
  assign mem[1178] = mem_1178_sv2v_reg;
  assign mem[1177] = mem_1177_sv2v_reg;
  assign mem[1176] = mem_1176_sv2v_reg;
  assign mem[1175] = mem_1175_sv2v_reg;
  assign mem[1174] = mem_1174_sv2v_reg;
  assign mem[1173] = mem_1173_sv2v_reg;
  assign mem[1172] = mem_1172_sv2v_reg;
  assign mem[1171] = mem_1171_sv2v_reg;
  assign mem[1170] = mem_1170_sv2v_reg;
  assign mem[1169] = mem_1169_sv2v_reg;
  assign mem[1168] = mem_1168_sv2v_reg;
  assign mem[1167] = mem_1167_sv2v_reg;
  assign mem[1166] = mem_1166_sv2v_reg;
  assign mem[1165] = mem_1165_sv2v_reg;
  assign mem[1164] = mem_1164_sv2v_reg;
  assign mem[1163] = mem_1163_sv2v_reg;
  assign mem[1162] = mem_1162_sv2v_reg;
  assign mem[1161] = mem_1161_sv2v_reg;
  assign mem[1160] = mem_1160_sv2v_reg;
  assign mem[1159] = mem_1159_sv2v_reg;
  assign mem[1158] = mem_1158_sv2v_reg;
  assign mem[1157] = mem_1157_sv2v_reg;
  assign mem[1156] = mem_1156_sv2v_reg;
  assign mem[1155] = mem_1155_sv2v_reg;
  assign mem[1154] = mem_1154_sv2v_reg;
  assign mem[1153] = mem_1153_sv2v_reg;
  assign mem[1152] = mem_1152_sv2v_reg;
  assign mem[1151] = mem_1151_sv2v_reg;
  assign mem[1150] = mem_1150_sv2v_reg;
  assign mem[1149] = mem_1149_sv2v_reg;
  assign mem[1148] = mem_1148_sv2v_reg;
  assign mem[1147] = mem_1147_sv2v_reg;
  assign mem[1146] = mem_1146_sv2v_reg;
  assign mem[1145] = mem_1145_sv2v_reg;
  assign mem[1144] = mem_1144_sv2v_reg;
  assign mem[1143] = mem_1143_sv2v_reg;
  assign mem[1142] = mem_1142_sv2v_reg;
  assign mem[1141] = mem_1141_sv2v_reg;
  assign mem[1140] = mem_1140_sv2v_reg;
  assign mem[1139] = mem_1139_sv2v_reg;
  assign mem[1138] = mem_1138_sv2v_reg;
  assign mem[1137] = mem_1137_sv2v_reg;
  assign mem[1136] = mem_1136_sv2v_reg;
  assign mem[1135] = mem_1135_sv2v_reg;
  assign mem[1134] = mem_1134_sv2v_reg;
  assign mem[1133] = mem_1133_sv2v_reg;
  assign mem[1132] = mem_1132_sv2v_reg;
  assign mem[1131] = mem_1131_sv2v_reg;
  assign mem[1130] = mem_1130_sv2v_reg;
  assign mem[1129] = mem_1129_sv2v_reg;
  assign mem[1128] = mem_1128_sv2v_reg;
  assign mem[1127] = mem_1127_sv2v_reg;
  assign mem[1126] = mem_1126_sv2v_reg;
  assign mem[1125] = mem_1125_sv2v_reg;
  assign mem[1124] = mem_1124_sv2v_reg;
  assign mem[1123] = mem_1123_sv2v_reg;
  assign mem[1122] = mem_1122_sv2v_reg;
  assign mem[1121] = mem_1121_sv2v_reg;
  assign mem[1120] = mem_1120_sv2v_reg;
  assign mem[1119] = mem_1119_sv2v_reg;
  assign mem[1118] = mem_1118_sv2v_reg;
  assign mem[1117] = mem_1117_sv2v_reg;
  assign mem[1116] = mem_1116_sv2v_reg;
  assign mem[1115] = mem_1115_sv2v_reg;
  assign mem[1114] = mem_1114_sv2v_reg;
  assign mem[1113] = mem_1113_sv2v_reg;
  assign mem[1112] = mem_1112_sv2v_reg;
  assign mem[1111] = mem_1111_sv2v_reg;
  assign mem[1110] = mem_1110_sv2v_reg;
  assign mem[1109] = mem_1109_sv2v_reg;
  assign mem[1108] = mem_1108_sv2v_reg;
  assign mem[1107] = mem_1107_sv2v_reg;
  assign mem[1106] = mem_1106_sv2v_reg;
  assign mem[1105] = mem_1105_sv2v_reg;
  assign mem[1104] = mem_1104_sv2v_reg;
  assign mem[1103] = mem_1103_sv2v_reg;
  assign mem[1102] = mem_1102_sv2v_reg;
  assign mem[1101] = mem_1101_sv2v_reg;
  assign mem[1100] = mem_1100_sv2v_reg;
  assign mem[1099] = mem_1099_sv2v_reg;
  assign mem[1098] = mem_1098_sv2v_reg;
  assign mem[1097] = mem_1097_sv2v_reg;
  assign mem[1096] = mem_1096_sv2v_reg;
  assign mem[1095] = mem_1095_sv2v_reg;
  assign mem[1094] = mem_1094_sv2v_reg;
  assign mem[1093] = mem_1093_sv2v_reg;
  assign mem[1092] = mem_1092_sv2v_reg;
  assign mem[1091] = mem_1091_sv2v_reg;
  assign mem[1090] = mem_1090_sv2v_reg;
  assign mem[1089] = mem_1089_sv2v_reg;
  assign mem[1088] = mem_1088_sv2v_reg;
  assign mem[1087] = mem_1087_sv2v_reg;
  assign mem[1086] = mem_1086_sv2v_reg;
  assign mem[1085] = mem_1085_sv2v_reg;
  assign mem[1084] = mem_1084_sv2v_reg;
  assign mem[1083] = mem_1083_sv2v_reg;
  assign mem[1082] = mem_1082_sv2v_reg;
  assign mem[1081] = mem_1081_sv2v_reg;
  assign mem[1080] = mem_1080_sv2v_reg;
  assign mem[1079] = mem_1079_sv2v_reg;
  assign mem[1078] = mem_1078_sv2v_reg;
  assign mem[1077] = mem_1077_sv2v_reg;
  assign mem[1076] = mem_1076_sv2v_reg;
  assign mem[1075] = mem_1075_sv2v_reg;
  assign mem[1074] = mem_1074_sv2v_reg;
  assign mem[1073] = mem_1073_sv2v_reg;
  assign mem[1072] = mem_1072_sv2v_reg;
  assign mem[1071] = mem_1071_sv2v_reg;
  assign mem[1070] = mem_1070_sv2v_reg;
  assign mem[1069] = mem_1069_sv2v_reg;
  assign mem[1068] = mem_1068_sv2v_reg;
  assign mem[1067] = mem_1067_sv2v_reg;
  assign mem[1066] = mem_1066_sv2v_reg;
  assign mem[1065] = mem_1065_sv2v_reg;
  assign mem[1064] = mem_1064_sv2v_reg;
  assign mem[1063] = mem_1063_sv2v_reg;
  assign mem[1062] = mem_1062_sv2v_reg;
  assign mem[1061] = mem_1061_sv2v_reg;
  assign mem[1060] = mem_1060_sv2v_reg;
  assign mem[1059] = mem_1059_sv2v_reg;
  assign mem[1058] = mem_1058_sv2v_reg;
  assign mem[1057] = mem_1057_sv2v_reg;
  assign mem[1056] = mem_1056_sv2v_reg;
  assign mem[1055] = mem_1055_sv2v_reg;
  assign mem[1054] = mem_1054_sv2v_reg;
  assign mem[1053] = mem_1053_sv2v_reg;
  assign mem[1052] = mem_1052_sv2v_reg;
  assign mem[1051] = mem_1051_sv2v_reg;
  assign mem[1050] = mem_1050_sv2v_reg;
  assign mem[1049] = mem_1049_sv2v_reg;
  assign mem[1048] = mem_1048_sv2v_reg;
  assign mem[1047] = mem_1047_sv2v_reg;
  assign mem[1046] = mem_1046_sv2v_reg;
  assign mem[1045] = mem_1045_sv2v_reg;
  assign mem[1044] = mem_1044_sv2v_reg;
  assign mem[1043] = mem_1043_sv2v_reg;
  assign mem[1042] = mem_1042_sv2v_reg;
  assign mem[1041] = mem_1041_sv2v_reg;
  assign mem[1040] = mem_1040_sv2v_reg;
  assign mem[1039] = mem_1039_sv2v_reg;
  assign mem[1038] = mem_1038_sv2v_reg;
  assign mem[1037] = mem_1037_sv2v_reg;
  assign mem[1036] = mem_1036_sv2v_reg;
  assign mem[1035] = mem_1035_sv2v_reg;
  assign mem[1034] = mem_1034_sv2v_reg;
  assign mem[1033] = mem_1033_sv2v_reg;
  assign mem[1032] = mem_1032_sv2v_reg;
  assign mem[1031] = mem_1031_sv2v_reg;
  assign mem[1030] = mem_1030_sv2v_reg;
  assign mem[1029] = mem_1029_sv2v_reg;
  assign mem[1028] = mem_1028_sv2v_reg;
  assign mem[1027] = mem_1027_sv2v_reg;
  assign mem[1026] = mem_1026_sv2v_reg;
  assign mem[1025] = mem_1025_sv2v_reg;
  assign mem[1024] = mem_1024_sv2v_reg;
  assign mem[1023] = mem_1023_sv2v_reg;
  assign mem[1022] = mem_1022_sv2v_reg;
  assign mem[1021] = mem_1021_sv2v_reg;
  assign mem[1020] = mem_1020_sv2v_reg;
  assign mem[1019] = mem_1019_sv2v_reg;
  assign mem[1018] = mem_1018_sv2v_reg;
  assign mem[1017] = mem_1017_sv2v_reg;
  assign mem[1016] = mem_1016_sv2v_reg;
  assign mem[1015] = mem_1015_sv2v_reg;
  assign mem[1014] = mem_1014_sv2v_reg;
  assign mem[1013] = mem_1013_sv2v_reg;
  assign mem[1012] = mem_1012_sv2v_reg;
  assign mem[1011] = mem_1011_sv2v_reg;
  assign mem[1010] = mem_1010_sv2v_reg;
  assign mem[1009] = mem_1009_sv2v_reg;
  assign mem[1008] = mem_1008_sv2v_reg;
  assign mem[1007] = mem_1007_sv2v_reg;
  assign mem[1006] = mem_1006_sv2v_reg;
  assign mem[1005] = mem_1005_sv2v_reg;
  assign mem[1004] = mem_1004_sv2v_reg;
  assign mem[1003] = mem_1003_sv2v_reg;
  assign mem[1002] = mem_1002_sv2v_reg;
  assign mem[1001] = mem_1001_sv2v_reg;
  assign mem[1000] = mem_1000_sv2v_reg;
  assign mem[999] = mem_999_sv2v_reg;
  assign mem[998] = mem_998_sv2v_reg;
  assign mem[997] = mem_997_sv2v_reg;
  assign mem[996] = mem_996_sv2v_reg;
  assign mem[995] = mem_995_sv2v_reg;
  assign mem[994] = mem_994_sv2v_reg;
  assign mem[993] = mem_993_sv2v_reg;
  assign mem[992] = mem_992_sv2v_reg;
  assign mem[991] = mem_991_sv2v_reg;
  assign mem[990] = mem_990_sv2v_reg;
  assign mem[989] = mem_989_sv2v_reg;
  assign mem[988] = mem_988_sv2v_reg;
  assign mem[987] = mem_987_sv2v_reg;
  assign mem[986] = mem_986_sv2v_reg;
  assign mem[985] = mem_985_sv2v_reg;
  assign mem[984] = mem_984_sv2v_reg;
  assign mem[983] = mem_983_sv2v_reg;
  assign mem[982] = mem_982_sv2v_reg;
  assign mem[981] = mem_981_sv2v_reg;
  assign mem[980] = mem_980_sv2v_reg;
  assign mem[979] = mem_979_sv2v_reg;
  assign mem[978] = mem_978_sv2v_reg;
  assign mem[977] = mem_977_sv2v_reg;
  assign mem[976] = mem_976_sv2v_reg;
  assign mem[975] = mem_975_sv2v_reg;
  assign mem[974] = mem_974_sv2v_reg;
  assign mem[973] = mem_973_sv2v_reg;
  assign mem[972] = mem_972_sv2v_reg;
  assign mem[971] = mem_971_sv2v_reg;
  assign mem[970] = mem_970_sv2v_reg;
  assign mem[969] = mem_969_sv2v_reg;
  assign mem[968] = mem_968_sv2v_reg;
  assign mem[967] = mem_967_sv2v_reg;
  assign mem[966] = mem_966_sv2v_reg;
  assign mem[965] = mem_965_sv2v_reg;
  assign mem[964] = mem_964_sv2v_reg;
  assign mem[963] = mem_963_sv2v_reg;
  assign mem[962] = mem_962_sv2v_reg;
  assign mem[961] = mem_961_sv2v_reg;
  assign mem[960] = mem_960_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_6_sv2v_reg <= addr_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_5_sv2v_reg <= addr_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_4_sv2v_reg <= addr_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_3_sv2v_reg <= addr_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_2_sv2v_reg <= addr_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_1_sv2v_reg <= addr_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_0_sv2v_reg <= addr_i[0];
    end 
  end

  assign data_o[14] = (N159)? mem[14] : 
                      (N161)? mem[29] : 
                      (N163)? mem[44] : 
                      (N165)? mem[59] : 
                      (N167)? mem[74] : 
                      (N169)? mem[89] : 
                      (N171)? mem[104] : 
                      (N173)? mem[119] : 
                      (N175)? mem[134] : 
                      (N177)? mem[149] : 
                      (N179)? mem[164] : 
                      (N181)? mem[179] : 
                      (N183)? mem[194] : 
                      (N185)? mem[209] : 
                      (N187)? mem[224] : 
                      (N189)? mem[239] : 
                      (N191)? mem[254] : 
                      (N193)? mem[269] : 
                      (N195)? mem[284] : 
                      (N197)? mem[299] : 
                      (N199)? mem[314] : 
                      (N201)? mem[329] : 
                      (N203)? mem[344] : 
                      (N205)? mem[359] : 
                      (N207)? mem[374] : 
                      (N209)? mem[389] : 
                      (N211)? mem[404] : 
                      (N213)? mem[419] : 
                      (N215)? mem[434] : 
                      (N217)? mem[449] : 
                      (N219)? mem[464] : 
                      (N221)? mem[479] : 
                      (N223)? mem[494] : 
                      (N225)? mem[509] : 
                      (N227)? mem[524] : 
                      (N229)? mem[539] : 
                      (N231)? mem[554] : 
                      (N233)? mem[569] : 
                      (N235)? mem[584] : 
                      (N237)? mem[599] : 
                      (N239)? mem[614] : 
                      (N241)? mem[629] : 
                      (N243)? mem[644] : 
                      (N245)? mem[659] : 
                      (N247)? mem[674] : 
                      (N249)? mem[689] : 
                      (N251)? mem[704] : 
                      (N253)? mem[719] : 
                      (N255)? mem[734] : 
                      (N257)? mem[749] : 
                      (N259)? mem[764] : 
                      (N261)? mem[779] : 
                      (N263)? mem[794] : 
                      (N265)? mem[809] : 
                      (N267)? mem[824] : 
                      (N269)? mem[839] : 
                      (N271)? mem[854] : 
                      (N273)? mem[869] : 
                      (N275)? mem[884] : 
                      (N277)? mem[899] : 
                      (N279)? mem[914] : 
                      (N281)? mem[929] : 
                      (N283)? mem[944] : 
                      (N285)? mem[959] : 
                      (N160)? mem[974] : 
                      (N162)? mem[989] : 
                      (N164)? mem[1004] : 
                      (N166)? mem[1019] : 
                      (N168)? mem[1034] : 
                      (N170)? mem[1049] : 
                      (N172)? mem[1064] : 
                      (N174)? mem[1079] : 
                      (N176)? mem[1094] : 
                      (N178)? mem[1109] : 
                      (N180)? mem[1124] : 
                      (N182)? mem[1139] : 
                      (N184)? mem[1154] : 
                      (N186)? mem[1169] : 
                      (N188)? mem[1184] : 
                      (N190)? mem[1199] : 
                      (N192)? mem[1214] : 
                      (N194)? mem[1229] : 
                      (N196)? mem[1244] : 
                      (N198)? mem[1259] : 
                      (N200)? mem[1274] : 
                      (N202)? mem[1289] : 
                      (N204)? mem[1304] : 
                      (N206)? mem[1319] : 
                      (N208)? mem[1334] : 
                      (N210)? mem[1349] : 
                      (N212)? mem[1364] : 
                      (N214)? mem[1379] : 
                      (N216)? mem[1394] : 
                      (N218)? mem[1409] : 
                      (N220)? mem[1424] : 
                      (N222)? mem[1439] : 
                      (N224)? mem[1454] : 
                      (N226)? mem[1469] : 
                      (N228)? mem[1484] : 
                      (N230)? mem[1499] : 
                      (N232)? mem[1514] : 
                      (N234)? mem[1529] : 
                      (N236)? mem[1544] : 
                      (N238)? mem[1559] : 
                      (N240)? mem[1574] : 
                      (N242)? mem[1589] : 
                      (N244)? mem[1604] : 
                      (N246)? mem[1619] : 
                      (N248)? mem[1634] : 
                      (N250)? mem[1649] : 
                      (N252)? mem[1664] : 
                      (N254)? mem[1679] : 
                      (N256)? mem[1694] : 
                      (N258)? mem[1709] : 
                      (N260)? mem[1724] : 
                      (N262)? mem[1739] : 
                      (N264)? mem[1754] : 
                      (N266)? mem[1769] : 
                      (N268)? mem[1784] : 
                      (N270)? mem[1799] : 
                      (N272)? mem[1814] : 
                      (N274)? mem[1829] : 
                      (N276)? mem[1844] : 
                      (N278)? mem[1859] : 
                      (N280)? mem[1874] : 
                      (N282)? mem[1889] : 
                      (N284)? mem[1904] : 
                      (N286)? mem[1919] : 1'b0;
  assign data_o[13] = (N159)? mem[13] : 
                      (N161)? mem[28] : 
                      (N163)? mem[43] : 
                      (N165)? mem[58] : 
                      (N167)? mem[73] : 
                      (N169)? mem[88] : 
                      (N171)? mem[103] : 
                      (N173)? mem[118] : 
                      (N175)? mem[133] : 
                      (N177)? mem[148] : 
                      (N179)? mem[163] : 
                      (N181)? mem[178] : 
                      (N183)? mem[193] : 
                      (N185)? mem[208] : 
                      (N187)? mem[223] : 
                      (N189)? mem[238] : 
                      (N191)? mem[253] : 
                      (N193)? mem[268] : 
                      (N195)? mem[283] : 
                      (N197)? mem[298] : 
                      (N199)? mem[313] : 
                      (N201)? mem[328] : 
                      (N203)? mem[343] : 
                      (N205)? mem[358] : 
                      (N207)? mem[373] : 
                      (N209)? mem[388] : 
                      (N211)? mem[403] : 
                      (N213)? mem[418] : 
                      (N215)? mem[433] : 
                      (N217)? mem[448] : 
                      (N219)? mem[463] : 
                      (N221)? mem[478] : 
                      (N223)? mem[493] : 
                      (N225)? mem[508] : 
                      (N227)? mem[523] : 
                      (N229)? mem[538] : 
                      (N231)? mem[553] : 
                      (N233)? mem[568] : 
                      (N235)? mem[583] : 
                      (N237)? mem[598] : 
                      (N239)? mem[613] : 
                      (N241)? mem[628] : 
                      (N243)? mem[643] : 
                      (N245)? mem[658] : 
                      (N247)? mem[673] : 
                      (N249)? mem[688] : 
                      (N251)? mem[703] : 
                      (N253)? mem[718] : 
                      (N255)? mem[733] : 
                      (N257)? mem[748] : 
                      (N259)? mem[763] : 
                      (N261)? mem[778] : 
                      (N263)? mem[793] : 
                      (N265)? mem[808] : 
                      (N267)? mem[823] : 
                      (N269)? mem[838] : 
                      (N271)? mem[853] : 
                      (N273)? mem[868] : 
                      (N275)? mem[883] : 
                      (N277)? mem[898] : 
                      (N279)? mem[913] : 
                      (N281)? mem[928] : 
                      (N283)? mem[943] : 
                      (N285)? mem[958] : 
                      (N160)? mem[973] : 
                      (N162)? mem[988] : 
                      (N164)? mem[1003] : 
                      (N166)? mem[1018] : 
                      (N168)? mem[1033] : 
                      (N170)? mem[1048] : 
                      (N172)? mem[1063] : 
                      (N174)? mem[1078] : 
                      (N176)? mem[1093] : 
                      (N178)? mem[1108] : 
                      (N180)? mem[1123] : 
                      (N182)? mem[1138] : 
                      (N184)? mem[1153] : 
                      (N186)? mem[1168] : 
                      (N188)? mem[1183] : 
                      (N190)? mem[1198] : 
                      (N192)? mem[1213] : 
                      (N194)? mem[1228] : 
                      (N196)? mem[1243] : 
                      (N198)? mem[1258] : 
                      (N200)? mem[1273] : 
                      (N202)? mem[1288] : 
                      (N204)? mem[1303] : 
                      (N206)? mem[1318] : 
                      (N208)? mem[1333] : 
                      (N210)? mem[1348] : 
                      (N212)? mem[1363] : 
                      (N214)? mem[1378] : 
                      (N216)? mem[1393] : 
                      (N218)? mem[1408] : 
                      (N220)? mem[1423] : 
                      (N222)? mem[1438] : 
                      (N224)? mem[1453] : 
                      (N226)? mem[1468] : 
                      (N228)? mem[1483] : 
                      (N230)? mem[1498] : 
                      (N232)? mem[1513] : 
                      (N234)? mem[1528] : 
                      (N236)? mem[1543] : 
                      (N238)? mem[1558] : 
                      (N240)? mem[1573] : 
                      (N242)? mem[1588] : 
                      (N244)? mem[1603] : 
                      (N246)? mem[1618] : 
                      (N248)? mem[1633] : 
                      (N250)? mem[1648] : 
                      (N252)? mem[1663] : 
                      (N254)? mem[1678] : 
                      (N256)? mem[1693] : 
                      (N258)? mem[1708] : 
                      (N260)? mem[1723] : 
                      (N262)? mem[1738] : 
                      (N264)? mem[1753] : 
                      (N266)? mem[1768] : 
                      (N268)? mem[1783] : 
                      (N270)? mem[1798] : 
                      (N272)? mem[1813] : 
                      (N274)? mem[1828] : 
                      (N276)? mem[1843] : 
                      (N278)? mem[1858] : 
                      (N280)? mem[1873] : 
                      (N282)? mem[1888] : 
                      (N284)? mem[1903] : 
                      (N286)? mem[1918] : 1'b0;
  assign data_o[12] = (N159)? mem[12] : 
                      (N161)? mem[27] : 
                      (N163)? mem[42] : 
                      (N165)? mem[57] : 
                      (N167)? mem[72] : 
                      (N169)? mem[87] : 
                      (N171)? mem[102] : 
                      (N173)? mem[117] : 
                      (N175)? mem[132] : 
                      (N177)? mem[147] : 
                      (N179)? mem[162] : 
                      (N181)? mem[177] : 
                      (N183)? mem[192] : 
                      (N185)? mem[207] : 
                      (N187)? mem[222] : 
                      (N189)? mem[237] : 
                      (N191)? mem[252] : 
                      (N193)? mem[267] : 
                      (N195)? mem[282] : 
                      (N197)? mem[297] : 
                      (N199)? mem[312] : 
                      (N201)? mem[327] : 
                      (N203)? mem[342] : 
                      (N205)? mem[357] : 
                      (N207)? mem[372] : 
                      (N209)? mem[387] : 
                      (N211)? mem[402] : 
                      (N213)? mem[417] : 
                      (N215)? mem[432] : 
                      (N217)? mem[447] : 
                      (N219)? mem[462] : 
                      (N221)? mem[477] : 
                      (N223)? mem[492] : 
                      (N225)? mem[507] : 
                      (N227)? mem[522] : 
                      (N229)? mem[537] : 
                      (N231)? mem[552] : 
                      (N233)? mem[567] : 
                      (N235)? mem[582] : 
                      (N237)? mem[597] : 
                      (N239)? mem[612] : 
                      (N241)? mem[627] : 
                      (N243)? mem[642] : 
                      (N245)? mem[657] : 
                      (N247)? mem[672] : 
                      (N249)? mem[687] : 
                      (N251)? mem[702] : 
                      (N253)? mem[717] : 
                      (N255)? mem[732] : 
                      (N257)? mem[747] : 
                      (N259)? mem[762] : 
                      (N261)? mem[777] : 
                      (N263)? mem[792] : 
                      (N265)? mem[807] : 
                      (N267)? mem[822] : 
                      (N269)? mem[837] : 
                      (N271)? mem[852] : 
                      (N273)? mem[867] : 
                      (N275)? mem[882] : 
                      (N277)? mem[897] : 
                      (N279)? mem[912] : 
                      (N281)? mem[927] : 
                      (N283)? mem[942] : 
                      (N285)? mem[957] : 
                      (N160)? mem[972] : 
                      (N162)? mem[987] : 
                      (N164)? mem[1002] : 
                      (N166)? mem[1017] : 
                      (N168)? mem[1032] : 
                      (N170)? mem[1047] : 
                      (N172)? mem[1062] : 
                      (N174)? mem[1077] : 
                      (N176)? mem[1092] : 
                      (N178)? mem[1107] : 
                      (N180)? mem[1122] : 
                      (N182)? mem[1137] : 
                      (N184)? mem[1152] : 
                      (N186)? mem[1167] : 
                      (N188)? mem[1182] : 
                      (N190)? mem[1197] : 
                      (N192)? mem[1212] : 
                      (N194)? mem[1227] : 
                      (N196)? mem[1242] : 
                      (N198)? mem[1257] : 
                      (N200)? mem[1272] : 
                      (N202)? mem[1287] : 
                      (N204)? mem[1302] : 
                      (N206)? mem[1317] : 
                      (N208)? mem[1332] : 
                      (N210)? mem[1347] : 
                      (N212)? mem[1362] : 
                      (N214)? mem[1377] : 
                      (N216)? mem[1392] : 
                      (N218)? mem[1407] : 
                      (N220)? mem[1422] : 
                      (N222)? mem[1437] : 
                      (N224)? mem[1452] : 
                      (N226)? mem[1467] : 
                      (N228)? mem[1482] : 
                      (N230)? mem[1497] : 
                      (N232)? mem[1512] : 
                      (N234)? mem[1527] : 
                      (N236)? mem[1542] : 
                      (N238)? mem[1557] : 
                      (N240)? mem[1572] : 
                      (N242)? mem[1587] : 
                      (N244)? mem[1602] : 
                      (N246)? mem[1617] : 
                      (N248)? mem[1632] : 
                      (N250)? mem[1647] : 
                      (N252)? mem[1662] : 
                      (N254)? mem[1677] : 
                      (N256)? mem[1692] : 
                      (N258)? mem[1707] : 
                      (N260)? mem[1722] : 
                      (N262)? mem[1737] : 
                      (N264)? mem[1752] : 
                      (N266)? mem[1767] : 
                      (N268)? mem[1782] : 
                      (N270)? mem[1797] : 
                      (N272)? mem[1812] : 
                      (N274)? mem[1827] : 
                      (N276)? mem[1842] : 
                      (N278)? mem[1857] : 
                      (N280)? mem[1872] : 
                      (N282)? mem[1887] : 
                      (N284)? mem[1902] : 
                      (N286)? mem[1917] : 1'b0;
  assign data_o[11] = (N159)? mem[11] : 
                      (N161)? mem[26] : 
                      (N163)? mem[41] : 
                      (N165)? mem[56] : 
                      (N167)? mem[71] : 
                      (N169)? mem[86] : 
                      (N171)? mem[101] : 
                      (N173)? mem[116] : 
                      (N175)? mem[131] : 
                      (N177)? mem[146] : 
                      (N179)? mem[161] : 
                      (N181)? mem[176] : 
                      (N183)? mem[191] : 
                      (N185)? mem[206] : 
                      (N187)? mem[221] : 
                      (N189)? mem[236] : 
                      (N191)? mem[251] : 
                      (N193)? mem[266] : 
                      (N195)? mem[281] : 
                      (N197)? mem[296] : 
                      (N199)? mem[311] : 
                      (N201)? mem[326] : 
                      (N203)? mem[341] : 
                      (N205)? mem[356] : 
                      (N207)? mem[371] : 
                      (N209)? mem[386] : 
                      (N211)? mem[401] : 
                      (N213)? mem[416] : 
                      (N215)? mem[431] : 
                      (N217)? mem[446] : 
                      (N219)? mem[461] : 
                      (N221)? mem[476] : 
                      (N223)? mem[491] : 
                      (N225)? mem[506] : 
                      (N227)? mem[521] : 
                      (N229)? mem[536] : 
                      (N231)? mem[551] : 
                      (N233)? mem[566] : 
                      (N235)? mem[581] : 
                      (N237)? mem[596] : 
                      (N239)? mem[611] : 
                      (N241)? mem[626] : 
                      (N243)? mem[641] : 
                      (N245)? mem[656] : 
                      (N247)? mem[671] : 
                      (N249)? mem[686] : 
                      (N251)? mem[701] : 
                      (N253)? mem[716] : 
                      (N255)? mem[731] : 
                      (N257)? mem[746] : 
                      (N259)? mem[761] : 
                      (N261)? mem[776] : 
                      (N263)? mem[791] : 
                      (N265)? mem[806] : 
                      (N267)? mem[821] : 
                      (N269)? mem[836] : 
                      (N271)? mem[851] : 
                      (N273)? mem[866] : 
                      (N275)? mem[881] : 
                      (N277)? mem[896] : 
                      (N279)? mem[911] : 
                      (N281)? mem[926] : 
                      (N283)? mem[941] : 
                      (N285)? mem[956] : 
                      (N160)? mem[971] : 
                      (N162)? mem[986] : 
                      (N164)? mem[1001] : 
                      (N166)? mem[1016] : 
                      (N168)? mem[1031] : 
                      (N170)? mem[1046] : 
                      (N172)? mem[1061] : 
                      (N174)? mem[1076] : 
                      (N176)? mem[1091] : 
                      (N178)? mem[1106] : 
                      (N180)? mem[1121] : 
                      (N182)? mem[1136] : 
                      (N184)? mem[1151] : 
                      (N186)? mem[1166] : 
                      (N188)? mem[1181] : 
                      (N190)? mem[1196] : 
                      (N192)? mem[1211] : 
                      (N194)? mem[1226] : 
                      (N196)? mem[1241] : 
                      (N198)? mem[1256] : 
                      (N200)? mem[1271] : 
                      (N202)? mem[1286] : 
                      (N204)? mem[1301] : 
                      (N206)? mem[1316] : 
                      (N208)? mem[1331] : 
                      (N210)? mem[1346] : 
                      (N212)? mem[1361] : 
                      (N214)? mem[1376] : 
                      (N216)? mem[1391] : 
                      (N218)? mem[1406] : 
                      (N220)? mem[1421] : 
                      (N222)? mem[1436] : 
                      (N224)? mem[1451] : 
                      (N226)? mem[1466] : 
                      (N228)? mem[1481] : 
                      (N230)? mem[1496] : 
                      (N232)? mem[1511] : 
                      (N234)? mem[1526] : 
                      (N236)? mem[1541] : 
                      (N238)? mem[1556] : 
                      (N240)? mem[1571] : 
                      (N242)? mem[1586] : 
                      (N244)? mem[1601] : 
                      (N246)? mem[1616] : 
                      (N248)? mem[1631] : 
                      (N250)? mem[1646] : 
                      (N252)? mem[1661] : 
                      (N254)? mem[1676] : 
                      (N256)? mem[1691] : 
                      (N258)? mem[1706] : 
                      (N260)? mem[1721] : 
                      (N262)? mem[1736] : 
                      (N264)? mem[1751] : 
                      (N266)? mem[1766] : 
                      (N268)? mem[1781] : 
                      (N270)? mem[1796] : 
                      (N272)? mem[1811] : 
                      (N274)? mem[1826] : 
                      (N276)? mem[1841] : 
                      (N278)? mem[1856] : 
                      (N280)? mem[1871] : 
                      (N282)? mem[1886] : 
                      (N284)? mem[1901] : 
                      (N286)? mem[1916] : 1'b0;
  assign data_o[10] = (N159)? mem[10] : 
                      (N161)? mem[25] : 
                      (N163)? mem[40] : 
                      (N165)? mem[55] : 
                      (N167)? mem[70] : 
                      (N169)? mem[85] : 
                      (N171)? mem[100] : 
                      (N173)? mem[115] : 
                      (N175)? mem[130] : 
                      (N177)? mem[145] : 
                      (N179)? mem[160] : 
                      (N181)? mem[175] : 
                      (N183)? mem[190] : 
                      (N185)? mem[205] : 
                      (N187)? mem[220] : 
                      (N189)? mem[235] : 
                      (N191)? mem[250] : 
                      (N193)? mem[265] : 
                      (N195)? mem[280] : 
                      (N197)? mem[295] : 
                      (N199)? mem[310] : 
                      (N201)? mem[325] : 
                      (N203)? mem[340] : 
                      (N205)? mem[355] : 
                      (N207)? mem[370] : 
                      (N209)? mem[385] : 
                      (N211)? mem[400] : 
                      (N213)? mem[415] : 
                      (N215)? mem[430] : 
                      (N217)? mem[445] : 
                      (N219)? mem[460] : 
                      (N221)? mem[475] : 
                      (N223)? mem[490] : 
                      (N225)? mem[505] : 
                      (N227)? mem[520] : 
                      (N229)? mem[535] : 
                      (N231)? mem[550] : 
                      (N233)? mem[565] : 
                      (N235)? mem[580] : 
                      (N237)? mem[595] : 
                      (N239)? mem[610] : 
                      (N241)? mem[625] : 
                      (N243)? mem[640] : 
                      (N245)? mem[655] : 
                      (N247)? mem[670] : 
                      (N249)? mem[685] : 
                      (N251)? mem[700] : 
                      (N253)? mem[715] : 
                      (N255)? mem[730] : 
                      (N257)? mem[745] : 
                      (N259)? mem[760] : 
                      (N261)? mem[775] : 
                      (N263)? mem[790] : 
                      (N265)? mem[805] : 
                      (N267)? mem[820] : 
                      (N269)? mem[835] : 
                      (N271)? mem[850] : 
                      (N273)? mem[865] : 
                      (N275)? mem[880] : 
                      (N277)? mem[895] : 
                      (N279)? mem[910] : 
                      (N281)? mem[925] : 
                      (N283)? mem[940] : 
                      (N285)? mem[955] : 
                      (N160)? mem[970] : 
                      (N162)? mem[985] : 
                      (N164)? mem[1000] : 
                      (N166)? mem[1015] : 
                      (N168)? mem[1030] : 
                      (N170)? mem[1045] : 
                      (N172)? mem[1060] : 
                      (N174)? mem[1075] : 
                      (N176)? mem[1090] : 
                      (N178)? mem[1105] : 
                      (N180)? mem[1120] : 
                      (N182)? mem[1135] : 
                      (N184)? mem[1150] : 
                      (N186)? mem[1165] : 
                      (N188)? mem[1180] : 
                      (N190)? mem[1195] : 
                      (N192)? mem[1210] : 
                      (N194)? mem[1225] : 
                      (N196)? mem[1240] : 
                      (N198)? mem[1255] : 
                      (N200)? mem[1270] : 
                      (N202)? mem[1285] : 
                      (N204)? mem[1300] : 
                      (N206)? mem[1315] : 
                      (N208)? mem[1330] : 
                      (N210)? mem[1345] : 
                      (N212)? mem[1360] : 
                      (N214)? mem[1375] : 
                      (N216)? mem[1390] : 
                      (N218)? mem[1405] : 
                      (N220)? mem[1420] : 
                      (N222)? mem[1435] : 
                      (N224)? mem[1450] : 
                      (N226)? mem[1465] : 
                      (N228)? mem[1480] : 
                      (N230)? mem[1495] : 
                      (N232)? mem[1510] : 
                      (N234)? mem[1525] : 
                      (N236)? mem[1540] : 
                      (N238)? mem[1555] : 
                      (N240)? mem[1570] : 
                      (N242)? mem[1585] : 
                      (N244)? mem[1600] : 
                      (N246)? mem[1615] : 
                      (N248)? mem[1630] : 
                      (N250)? mem[1645] : 
                      (N252)? mem[1660] : 
                      (N254)? mem[1675] : 
                      (N256)? mem[1690] : 
                      (N258)? mem[1705] : 
                      (N260)? mem[1720] : 
                      (N262)? mem[1735] : 
                      (N264)? mem[1750] : 
                      (N266)? mem[1765] : 
                      (N268)? mem[1780] : 
                      (N270)? mem[1795] : 
                      (N272)? mem[1810] : 
                      (N274)? mem[1825] : 
                      (N276)? mem[1840] : 
                      (N278)? mem[1855] : 
                      (N280)? mem[1870] : 
                      (N282)? mem[1885] : 
                      (N284)? mem[1900] : 
                      (N286)? mem[1915] : 1'b0;
  assign data_o[9] = (N159)? mem[9] : 
                     (N161)? mem[24] : 
                     (N163)? mem[39] : 
                     (N165)? mem[54] : 
                     (N167)? mem[69] : 
                     (N169)? mem[84] : 
                     (N171)? mem[99] : 
                     (N173)? mem[114] : 
                     (N175)? mem[129] : 
                     (N177)? mem[144] : 
                     (N179)? mem[159] : 
                     (N181)? mem[174] : 
                     (N183)? mem[189] : 
                     (N185)? mem[204] : 
                     (N187)? mem[219] : 
                     (N189)? mem[234] : 
                     (N191)? mem[249] : 
                     (N193)? mem[264] : 
                     (N195)? mem[279] : 
                     (N197)? mem[294] : 
                     (N199)? mem[309] : 
                     (N201)? mem[324] : 
                     (N203)? mem[339] : 
                     (N205)? mem[354] : 
                     (N207)? mem[369] : 
                     (N209)? mem[384] : 
                     (N211)? mem[399] : 
                     (N213)? mem[414] : 
                     (N215)? mem[429] : 
                     (N217)? mem[444] : 
                     (N219)? mem[459] : 
                     (N221)? mem[474] : 
                     (N223)? mem[489] : 
                     (N225)? mem[504] : 
                     (N227)? mem[519] : 
                     (N229)? mem[534] : 
                     (N231)? mem[549] : 
                     (N233)? mem[564] : 
                     (N235)? mem[579] : 
                     (N237)? mem[594] : 
                     (N239)? mem[609] : 
                     (N241)? mem[624] : 
                     (N243)? mem[639] : 
                     (N245)? mem[654] : 
                     (N247)? mem[669] : 
                     (N249)? mem[684] : 
                     (N251)? mem[699] : 
                     (N253)? mem[714] : 
                     (N255)? mem[729] : 
                     (N257)? mem[744] : 
                     (N259)? mem[759] : 
                     (N261)? mem[774] : 
                     (N263)? mem[789] : 
                     (N265)? mem[804] : 
                     (N267)? mem[819] : 
                     (N269)? mem[834] : 
                     (N271)? mem[849] : 
                     (N273)? mem[864] : 
                     (N275)? mem[879] : 
                     (N277)? mem[894] : 
                     (N279)? mem[909] : 
                     (N281)? mem[924] : 
                     (N283)? mem[939] : 
                     (N285)? mem[954] : 
                     (N160)? mem[969] : 
                     (N162)? mem[984] : 
                     (N164)? mem[999] : 
                     (N166)? mem[1014] : 
                     (N168)? mem[1029] : 
                     (N170)? mem[1044] : 
                     (N172)? mem[1059] : 
                     (N174)? mem[1074] : 
                     (N176)? mem[1089] : 
                     (N178)? mem[1104] : 
                     (N180)? mem[1119] : 
                     (N182)? mem[1134] : 
                     (N184)? mem[1149] : 
                     (N186)? mem[1164] : 
                     (N188)? mem[1179] : 
                     (N190)? mem[1194] : 
                     (N192)? mem[1209] : 
                     (N194)? mem[1224] : 
                     (N196)? mem[1239] : 
                     (N198)? mem[1254] : 
                     (N200)? mem[1269] : 
                     (N202)? mem[1284] : 
                     (N204)? mem[1299] : 
                     (N206)? mem[1314] : 
                     (N208)? mem[1329] : 
                     (N210)? mem[1344] : 
                     (N212)? mem[1359] : 
                     (N214)? mem[1374] : 
                     (N216)? mem[1389] : 
                     (N218)? mem[1404] : 
                     (N220)? mem[1419] : 
                     (N222)? mem[1434] : 
                     (N224)? mem[1449] : 
                     (N226)? mem[1464] : 
                     (N228)? mem[1479] : 
                     (N230)? mem[1494] : 
                     (N232)? mem[1509] : 
                     (N234)? mem[1524] : 
                     (N236)? mem[1539] : 
                     (N238)? mem[1554] : 
                     (N240)? mem[1569] : 
                     (N242)? mem[1584] : 
                     (N244)? mem[1599] : 
                     (N246)? mem[1614] : 
                     (N248)? mem[1629] : 
                     (N250)? mem[1644] : 
                     (N252)? mem[1659] : 
                     (N254)? mem[1674] : 
                     (N256)? mem[1689] : 
                     (N258)? mem[1704] : 
                     (N260)? mem[1719] : 
                     (N262)? mem[1734] : 
                     (N264)? mem[1749] : 
                     (N266)? mem[1764] : 
                     (N268)? mem[1779] : 
                     (N270)? mem[1794] : 
                     (N272)? mem[1809] : 
                     (N274)? mem[1824] : 
                     (N276)? mem[1839] : 
                     (N278)? mem[1854] : 
                     (N280)? mem[1869] : 
                     (N282)? mem[1884] : 
                     (N284)? mem[1899] : 
                     (N286)? mem[1914] : 1'b0;
  assign data_o[8] = (N159)? mem[8] : 
                     (N161)? mem[23] : 
                     (N163)? mem[38] : 
                     (N165)? mem[53] : 
                     (N167)? mem[68] : 
                     (N169)? mem[83] : 
                     (N171)? mem[98] : 
                     (N173)? mem[113] : 
                     (N175)? mem[128] : 
                     (N177)? mem[143] : 
                     (N179)? mem[158] : 
                     (N181)? mem[173] : 
                     (N183)? mem[188] : 
                     (N185)? mem[203] : 
                     (N187)? mem[218] : 
                     (N189)? mem[233] : 
                     (N191)? mem[248] : 
                     (N193)? mem[263] : 
                     (N195)? mem[278] : 
                     (N197)? mem[293] : 
                     (N199)? mem[308] : 
                     (N201)? mem[323] : 
                     (N203)? mem[338] : 
                     (N205)? mem[353] : 
                     (N207)? mem[368] : 
                     (N209)? mem[383] : 
                     (N211)? mem[398] : 
                     (N213)? mem[413] : 
                     (N215)? mem[428] : 
                     (N217)? mem[443] : 
                     (N219)? mem[458] : 
                     (N221)? mem[473] : 
                     (N223)? mem[488] : 
                     (N225)? mem[503] : 
                     (N227)? mem[518] : 
                     (N229)? mem[533] : 
                     (N231)? mem[548] : 
                     (N233)? mem[563] : 
                     (N235)? mem[578] : 
                     (N237)? mem[593] : 
                     (N239)? mem[608] : 
                     (N241)? mem[623] : 
                     (N243)? mem[638] : 
                     (N245)? mem[653] : 
                     (N247)? mem[668] : 
                     (N249)? mem[683] : 
                     (N251)? mem[698] : 
                     (N253)? mem[713] : 
                     (N255)? mem[728] : 
                     (N257)? mem[743] : 
                     (N259)? mem[758] : 
                     (N261)? mem[773] : 
                     (N263)? mem[788] : 
                     (N265)? mem[803] : 
                     (N267)? mem[818] : 
                     (N269)? mem[833] : 
                     (N271)? mem[848] : 
                     (N273)? mem[863] : 
                     (N275)? mem[878] : 
                     (N277)? mem[893] : 
                     (N279)? mem[908] : 
                     (N281)? mem[923] : 
                     (N283)? mem[938] : 
                     (N285)? mem[953] : 
                     (N160)? mem[968] : 
                     (N162)? mem[983] : 
                     (N164)? mem[998] : 
                     (N166)? mem[1013] : 
                     (N168)? mem[1028] : 
                     (N170)? mem[1043] : 
                     (N172)? mem[1058] : 
                     (N174)? mem[1073] : 
                     (N176)? mem[1088] : 
                     (N178)? mem[1103] : 
                     (N180)? mem[1118] : 
                     (N182)? mem[1133] : 
                     (N184)? mem[1148] : 
                     (N186)? mem[1163] : 
                     (N188)? mem[1178] : 
                     (N190)? mem[1193] : 
                     (N192)? mem[1208] : 
                     (N194)? mem[1223] : 
                     (N196)? mem[1238] : 
                     (N198)? mem[1253] : 
                     (N200)? mem[1268] : 
                     (N202)? mem[1283] : 
                     (N204)? mem[1298] : 
                     (N206)? mem[1313] : 
                     (N208)? mem[1328] : 
                     (N210)? mem[1343] : 
                     (N212)? mem[1358] : 
                     (N214)? mem[1373] : 
                     (N216)? mem[1388] : 
                     (N218)? mem[1403] : 
                     (N220)? mem[1418] : 
                     (N222)? mem[1433] : 
                     (N224)? mem[1448] : 
                     (N226)? mem[1463] : 
                     (N228)? mem[1478] : 
                     (N230)? mem[1493] : 
                     (N232)? mem[1508] : 
                     (N234)? mem[1523] : 
                     (N236)? mem[1538] : 
                     (N238)? mem[1553] : 
                     (N240)? mem[1568] : 
                     (N242)? mem[1583] : 
                     (N244)? mem[1598] : 
                     (N246)? mem[1613] : 
                     (N248)? mem[1628] : 
                     (N250)? mem[1643] : 
                     (N252)? mem[1658] : 
                     (N254)? mem[1673] : 
                     (N256)? mem[1688] : 
                     (N258)? mem[1703] : 
                     (N260)? mem[1718] : 
                     (N262)? mem[1733] : 
                     (N264)? mem[1748] : 
                     (N266)? mem[1763] : 
                     (N268)? mem[1778] : 
                     (N270)? mem[1793] : 
                     (N272)? mem[1808] : 
                     (N274)? mem[1823] : 
                     (N276)? mem[1838] : 
                     (N278)? mem[1853] : 
                     (N280)? mem[1868] : 
                     (N282)? mem[1883] : 
                     (N284)? mem[1898] : 
                     (N286)? mem[1913] : 1'b0;
  assign data_o[7] = (N159)? mem[7] : 
                     (N161)? mem[22] : 
                     (N163)? mem[37] : 
                     (N165)? mem[52] : 
                     (N167)? mem[67] : 
                     (N169)? mem[82] : 
                     (N171)? mem[97] : 
                     (N173)? mem[112] : 
                     (N175)? mem[127] : 
                     (N177)? mem[142] : 
                     (N179)? mem[157] : 
                     (N181)? mem[172] : 
                     (N183)? mem[187] : 
                     (N185)? mem[202] : 
                     (N187)? mem[217] : 
                     (N189)? mem[232] : 
                     (N191)? mem[247] : 
                     (N193)? mem[262] : 
                     (N195)? mem[277] : 
                     (N197)? mem[292] : 
                     (N199)? mem[307] : 
                     (N201)? mem[322] : 
                     (N203)? mem[337] : 
                     (N205)? mem[352] : 
                     (N207)? mem[367] : 
                     (N209)? mem[382] : 
                     (N211)? mem[397] : 
                     (N213)? mem[412] : 
                     (N215)? mem[427] : 
                     (N217)? mem[442] : 
                     (N219)? mem[457] : 
                     (N221)? mem[472] : 
                     (N223)? mem[487] : 
                     (N225)? mem[502] : 
                     (N227)? mem[517] : 
                     (N229)? mem[532] : 
                     (N231)? mem[547] : 
                     (N233)? mem[562] : 
                     (N235)? mem[577] : 
                     (N237)? mem[592] : 
                     (N239)? mem[607] : 
                     (N241)? mem[622] : 
                     (N243)? mem[637] : 
                     (N245)? mem[652] : 
                     (N247)? mem[667] : 
                     (N249)? mem[682] : 
                     (N251)? mem[697] : 
                     (N253)? mem[712] : 
                     (N255)? mem[727] : 
                     (N257)? mem[742] : 
                     (N259)? mem[757] : 
                     (N261)? mem[772] : 
                     (N263)? mem[787] : 
                     (N265)? mem[802] : 
                     (N267)? mem[817] : 
                     (N269)? mem[832] : 
                     (N271)? mem[847] : 
                     (N273)? mem[862] : 
                     (N275)? mem[877] : 
                     (N277)? mem[892] : 
                     (N279)? mem[907] : 
                     (N281)? mem[922] : 
                     (N283)? mem[937] : 
                     (N285)? mem[952] : 
                     (N160)? mem[967] : 
                     (N162)? mem[982] : 
                     (N164)? mem[997] : 
                     (N166)? mem[1012] : 
                     (N168)? mem[1027] : 
                     (N170)? mem[1042] : 
                     (N172)? mem[1057] : 
                     (N174)? mem[1072] : 
                     (N176)? mem[1087] : 
                     (N178)? mem[1102] : 
                     (N180)? mem[1117] : 
                     (N182)? mem[1132] : 
                     (N184)? mem[1147] : 
                     (N186)? mem[1162] : 
                     (N188)? mem[1177] : 
                     (N190)? mem[1192] : 
                     (N192)? mem[1207] : 
                     (N194)? mem[1222] : 
                     (N196)? mem[1237] : 
                     (N198)? mem[1252] : 
                     (N200)? mem[1267] : 
                     (N202)? mem[1282] : 
                     (N204)? mem[1297] : 
                     (N206)? mem[1312] : 
                     (N208)? mem[1327] : 
                     (N210)? mem[1342] : 
                     (N212)? mem[1357] : 
                     (N214)? mem[1372] : 
                     (N216)? mem[1387] : 
                     (N218)? mem[1402] : 
                     (N220)? mem[1417] : 
                     (N222)? mem[1432] : 
                     (N224)? mem[1447] : 
                     (N226)? mem[1462] : 
                     (N228)? mem[1477] : 
                     (N230)? mem[1492] : 
                     (N232)? mem[1507] : 
                     (N234)? mem[1522] : 
                     (N236)? mem[1537] : 
                     (N238)? mem[1552] : 
                     (N240)? mem[1567] : 
                     (N242)? mem[1582] : 
                     (N244)? mem[1597] : 
                     (N246)? mem[1612] : 
                     (N248)? mem[1627] : 
                     (N250)? mem[1642] : 
                     (N252)? mem[1657] : 
                     (N254)? mem[1672] : 
                     (N256)? mem[1687] : 
                     (N258)? mem[1702] : 
                     (N260)? mem[1717] : 
                     (N262)? mem[1732] : 
                     (N264)? mem[1747] : 
                     (N266)? mem[1762] : 
                     (N268)? mem[1777] : 
                     (N270)? mem[1792] : 
                     (N272)? mem[1807] : 
                     (N274)? mem[1822] : 
                     (N276)? mem[1837] : 
                     (N278)? mem[1852] : 
                     (N280)? mem[1867] : 
                     (N282)? mem[1882] : 
                     (N284)? mem[1897] : 
                     (N286)? mem[1912] : 1'b0;
  assign data_o[6] = (N159)? mem[6] : 
                     (N161)? mem[21] : 
                     (N163)? mem[36] : 
                     (N165)? mem[51] : 
                     (N167)? mem[66] : 
                     (N169)? mem[81] : 
                     (N171)? mem[96] : 
                     (N173)? mem[111] : 
                     (N175)? mem[126] : 
                     (N177)? mem[141] : 
                     (N179)? mem[156] : 
                     (N181)? mem[171] : 
                     (N183)? mem[186] : 
                     (N185)? mem[201] : 
                     (N187)? mem[216] : 
                     (N189)? mem[231] : 
                     (N191)? mem[246] : 
                     (N193)? mem[261] : 
                     (N195)? mem[276] : 
                     (N197)? mem[291] : 
                     (N199)? mem[306] : 
                     (N201)? mem[321] : 
                     (N203)? mem[336] : 
                     (N205)? mem[351] : 
                     (N207)? mem[366] : 
                     (N209)? mem[381] : 
                     (N211)? mem[396] : 
                     (N213)? mem[411] : 
                     (N215)? mem[426] : 
                     (N217)? mem[441] : 
                     (N219)? mem[456] : 
                     (N221)? mem[471] : 
                     (N223)? mem[486] : 
                     (N225)? mem[501] : 
                     (N227)? mem[516] : 
                     (N229)? mem[531] : 
                     (N231)? mem[546] : 
                     (N233)? mem[561] : 
                     (N235)? mem[576] : 
                     (N237)? mem[591] : 
                     (N239)? mem[606] : 
                     (N241)? mem[621] : 
                     (N243)? mem[636] : 
                     (N245)? mem[651] : 
                     (N247)? mem[666] : 
                     (N249)? mem[681] : 
                     (N251)? mem[696] : 
                     (N253)? mem[711] : 
                     (N255)? mem[726] : 
                     (N257)? mem[741] : 
                     (N259)? mem[756] : 
                     (N261)? mem[771] : 
                     (N263)? mem[786] : 
                     (N265)? mem[801] : 
                     (N267)? mem[816] : 
                     (N269)? mem[831] : 
                     (N271)? mem[846] : 
                     (N273)? mem[861] : 
                     (N275)? mem[876] : 
                     (N277)? mem[891] : 
                     (N279)? mem[906] : 
                     (N281)? mem[921] : 
                     (N283)? mem[936] : 
                     (N285)? mem[951] : 
                     (N160)? mem[966] : 
                     (N162)? mem[981] : 
                     (N164)? mem[996] : 
                     (N166)? mem[1011] : 
                     (N168)? mem[1026] : 
                     (N170)? mem[1041] : 
                     (N172)? mem[1056] : 
                     (N174)? mem[1071] : 
                     (N176)? mem[1086] : 
                     (N178)? mem[1101] : 
                     (N180)? mem[1116] : 
                     (N182)? mem[1131] : 
                     (N184)? mem[1146] : 
                     (N186)? mem[1161] : 
                     (N188)? mem[1176] : 
                     (N190)? mem[1191] : 
                     (N192)? mem[1206] : 
                     (N194)? mem[1221] : 
                     (N196)? mem[1236] : 
                     (N198)? mem[1251] : 
                     (N200)? mem[1266] : 
                     (N202)? mem[1281] : 
                     (N204)? mem[1296] : 
                     (N206)? mem[1311] : 
                     (N208)? mem[1326] : 
                     (N210)? mem[1341] : 
                     (N212)? mem[1356] : 
                     (N214)? mem[1371] : 
                     (N216)? mem[1386] : 
                     (N218)? mem[1401] : 
                     (N220)? mem[1416] : 
                     (N222)? mem[1431] : 
                     (N224)? mem[1446] : 
                     (N226)? mem[1461] : 
                     (N228)? mem[1476] : 
                     (N230)? mem[1491] : 
                     (N232)? mem[1506] : 
                     (N234)? mem[1521] : 
                     (N236)? mem[1536] : 
                     (N238)? mem[1551] : 
                     (N240)? mem[1566] : 
                     (N242)? mem[1581] : 
                     (N244)? mem[1596] : 
                     (N246)? mem[1611] : 
                     (N248)? mem[1626] : 
                     (N250)? mem[1641] : 
                     (N252)? mem[1656] : 
                     (N254)? mem[1671] : 
                     (N256)? mem[1686] : 
                     (N258)? mem[1701] : 
                     (N260)? mem[1716] : 
                     (N262)? mem[1731] : 
                     (N264)? mem[1746] : 
                     (N266)? mem[1761] : 
                     (N268)? mem[1776] : 
                     (N270)? mem[1791] : 
                     (N272)? mem[1806] : 
                     (N274)? mem[1821] : 
                     (N276)? mem[1836] : 
                     (N278)? mem[1851] : 
                     (N280)? mem[1866] : 
                     (N282)? mem[1881] : 
                     (N284)? mem[1896] : 
                     (N286)? mem[1911] : 1'b0;
  assign data_o[5] = (N159)? mem[5] : 
                     (N161)? mem[20] : 
                     (N163)? mem[35] : 
                     (N165)? mem[50] : 
                     (N167)? mem[65] : 
                     (N169)? mem[80] : 
                     (N171)? mem[95] : 
                     (N173)? mem[110] : 
                     (N175)? mem[125] : 
                     (N177)? mem[140] : 
                     (N179)? mem[155] : 
                     (N181)? mem[170] : 
                     (N183)? mem[185] : 
                     (N185)? mem[200] : 
                     (N187)? mem[215] : 
                     (N189)? mem[230] : 
                     (N191)? mem[245] : 
                     (N193)? mem[260] : 
                     (N195)? mem[275] : 
                     (N197)? mem[290] : 
                     (N199)? mem[305] : 
                     (N201)? mem[320] : 
                     (N203)? mem[335] : 
                     (N205)? mem[350] : 
                     (N207)? mem[365] : 
                     (N209)? mem[380] : 
                     (N211)? mem[395] : 
                     (N213)? mem[410] : 
                     (N215)? mem[425] : 
                     (N217)? mem[440] : 
                     (N219)? mem[455] : 
                     (N221)? mem[470] : 
                     (N223)? mem[485] : 
                     (N225)? mem[500] : 
                     (N227)? mem[515] : 
                     (N229)? mem[530] : 
                     (N231)? mem[545] : 
                     (N233)? mem[560] : 
                     (N235)? mem[575] : 
                     (N237)? mem[590] : 
                     (N239)? mem[605] : 
                     (N241)? mem[620] : 
                     (N243)? mem[635] : 
                     (N245)? mem[650] : 
                     (N247)? mem[665] : 
                     (N249)? mem[680] : 
                     (N251)? mem[695] : 
                     (N253)? mem[710] : 
                     (N255)? mem[725] : 
                     (N257)? mem[740] : 
                     (N259)? mem[755] : 
                     (N261)? mem[770] : 
                     (N263)? mem[785] : 
                     (N265)? mem[800] : 
                     (N267)? mem[815] : 
                     (N269)? mem[830] : 
                     (N271)? mem[845] : 
                     (N273)? mem[860] : 
                     (N275)? mem[875] : 
                     (N277)? mem[890] : 
                     (N279)? mem[905] : 
                     (N281)? mem[920] : 
                     (N283)? mem[935] : 
                     (N285)? mem[950] : 
                     (N160)? mem[965] : 
                     (N162)? mem[980] : 
                     (N164)? mem[995] : 
                     (N166)? mem[1010] : 
                     (N168)? mem[1025] : 
                     (N170)? mem[1040] : 
                     (N172)? mem[1055] : 
                     (N174)? mem[1070] : 
                     (N176)? mem[1085] : 
                     (N178)? mem[1100] : 
                     (N180)? mem[1115] : 
                     (N182)? mem[1130] : 
                     (N184)? mem[1145] : 
                     (N186)? mem[1160] : 
                     (N188)? mem[1175] : 
                     (N190)? mem[1190] : 
                     (N192)? mem[1205] : 
                     (N194)? mem[1220] : 
                     (N196)? mem[1235] : 
                     (N198)? mem[1250] : 
                     (N200)? mem[1265] : 
                     (N202)? mem[1280] : 
                     (N204)? mem[1295] : 
                     (N206)? mem[1310] : 
                     (N208)? mem[1325] : 
                     (N210)? mem[1340] : 
                     (N212)? mem[1355] : 
                     (N214)? mem[1370] : 
                     (N216)? mem[1385] : 
                     (N218)? mem[1400] : 
                     (N220)? mem[1415] : 
                     (N222)? mem[1430] : 
                     (N224)? mem[1445] : 
                     (N226)? mem[1460] : 
                     (N228)? mem[1475] : 
                     (N230)? mem[1490] : 
                     (N232)? mem[1505] : 
                     (N234)? mem[1520] : 
                     (N236)? mem[1535] : 
                     (N238)? mem[1550] : 
                     (N240)? mem[1565] : 
                     (N242)? mem[1580] : 
                     (N244)? mem[1595] : 
                     (N246)? mem[1610] : 
                     (N248)? mem[1625] : 
                     (N250)? mem[1640] : 
                     (N252)? mem[1655] : 
                     (N254)? mem[1670] : 
                     (N256)? mem[1685] : 
                     (N258)? mem[1700] : 
                     (N260)? mem[1715] : 
                     (N262)? mem[1730] : 
                     (N264)? mem[1745] : 
                     (N266)? mem[1760] : 
                     (N268)? mem[1775] : 
                     (N270)? mem[1790] : 
                     (N272)? mem[1805] : 
                     (N274)? mem[1820] : 
                     (N276)? mem[1835] : 
                     (N278)? mem[1850] : 
                     (N280)? mem[1865] : 
                     (N282)? mem[1880] : 
                     (N284)? mem[1895] : 
                     (N286)? mem[1910] : 1'b0;
  assign data_o[4] = (N159)? mem[4] : 
                     (N161)? mem[19] : 
                     (N163)? mem[34] : 
                     (N165)? mem[49] : 
                     (N167)? mem[64] : 
                     (N169)? mem[79] : 
                     (N171)? mem[94] : 
                     (N173)? mem[109] : 
                     (N175)? mem[124] : 
                     (N177)? mem[139] : 
                     (N179)? mem[154] : 
                     (N181)? mem[169] : 
                     (N183)? mem[184] : 
                     (N185)? mem[199] : 
                     (N187)? mem[214] : 
                     (N189)? mem[229] : 
                     (N191)? mem[244] : 
                     (N193)? mem[259] : 
                     (N195)? mem[274] : 
                     (N197)? mem[289] : 
                     (N199)? mem[304] : 
                     (N201)? mem[319] : 
                     (N203)? mem[334] : 
                     (N205)? mem[349] : 
                     (N207)? mem[364] : 
                     (N209)? mem[379] : 
                     (N211)? mem[394] : 
                     (N213)? mem[409] : 
                     (N215)? mem[424] : 
                     (N217)? mem[439] : 
                     (N219)? mem[454] : 
                     (N221)? mem[469] : 
                     (N223)? mem[484] : 
                     (N225)? mem[499] : 
                     (N227)? mem[514] : 
                     (N229)? mem[529] : 
                     (N231)? mem[544] : 
                     (N233)? mem[559] : 
                     (N235)? mem[574] : 
                     (N237)? mem[589] : 
                     (N239)? mem[604] : 
                     (N241)? mem[619] : 
                     (N243)? mem[634] : 
                     (N245)? mem[649] : 
                     (N247)? mem[664] : 
                     (N249)? mem[679] : 
                     (N251)? mem[694] : 
                     (N253)? mem[709] : 
                     (N255)? mem[724] : 
                     (N257)? mem[739] : 
                     (N259)? mem[754] : 
                     (N261)? mem[769] : 
                     (N263)? mem[784] : 
                     (N265)? mem[799] : 
                     (N267)? mem[814] : 
                     (N269)? mem[829] : 
                     (N271)? mem[844] : 
                     (N273)? mem[859] : 
                     (N275)? mem[874] : 
                     (N277)? mem[889] : 
                     (N279)? mem[904] : 
                     (N281)? mem[919] : 
                     (N283)? mem[934] : 
                     (N285)? mem[949] : 
                     (N160)? mem[964] : 
                     (N162)? mem[979] : 
                     (N164)? mem[994] : 
                     (N166)? mem[1009] : 
                     (N168)? mem[1024] : 
                     (N170)? mem[1039] : 
                     (N172)? mem[1054] : 
                     (N174)? mem[1069] : 
                     (N176)? mem[1084] : 
                     (N178)? mem[1099] : 
                     (N180)? mem[1114] : 
                     (N182)? mem[1129] : 
                     (N184)? mem[1144] : 
                     (N186)? mem[1159] : 
                     (N188)? mem[1174] : 
                     (N190)? mem[1189] : 
                     (N192)? mem[1204] : 
                     (N194)? mem[1219] : 
                     (N196)? mem[1234] : 
                     (N198)? mem[1249] : 
                     (N200)? mem[1264] : 
                     (N202)? mem[1279] : 
                     (N204)? mem[1294] : 
                     (N206)? mem[1309] : 
                     (N208)? mem[1324] : 
                     (N210)? mem[1339] : 
                     (N212)? mem[1354] : 
                     (N214)? mem[1369] : 
                     (N216)? mem[1384] : 
                     (N218)? mem[1399] : 
                     (N220)? mem[1414] : 
                     (N222)? mem[1429] : 
                     (N224)? mem[1444] : 
                     (N226)? mem[1459] : 
                     (N228)? mem[1474] : 
                     (N230)? mem[1489] : 
                     (N232)? mem[1504] : 
                     (N234)? mem[1519] : 
                     (N236)? mem[1534] : 
                     (N238)? mem[1549] : 
                     (N240)? mem[1564] : 
                     (N242)? mem[1579] : 
                     (N244)? mem[1594] : 
                     (N246)? mem[1609] : 
                     (N248)? mem[1624] : 
                     (N250)? mem[1639] : 
                     (N252)? mem[1654] : 
                     (N254)? mem[1669] : 
                     (N256)? mem[1684] : 
                     (N258)? mem[1699] : 
                     (N260)? mem[1714] : 
                     (N262)? mem[1729] : 
                     (N264)? mem[1744] : 
                     (N266)? mem[1759] : 
                     (N268)? mem[1774] : 
                     (N270)? mem[1789] : 
                     (N272)? mem[1804] : 
                     (N274)? mem[1819] : 
                     (N276)? mem[1834] : 
                     (N278)? mem[1849] : 
                     (N280)? mem[1864] : 
                     (N282)? mem[1879] : 
                     (N284)? mem[1894] : 
                     (N286)? mem[1909] : 1'b0;
  assign data_o[3] = (N159)? mem[3] : 
                     (N161)? mem[18] : 
                     (N163)? mem[33] : 
                     (N165)? mem[48] : 
                     (N167)? mem[63] : 
                     (N169)? mem[78] : 
                     (N171)? mem[93] : 
                     (N173)? mem[108] : 
                     (N175)? mem[123] : 
                     (N177)? mem[138] : 
                     (N179)? mem[153] : 
                     (N181)? mem[168] : 
                     (N183)? mem[183] : 
                     (N185)? mem[198] : 
                     (N187)? mem[213] : 
                     (N189)? mem[228] : 
                     (N191)? mem[243] : 
                     (N193)? mem[258] : 
                     (N195)? mem[273] : 
                     (N197)? mem[288] : 
                     (N199)? mem[303] : 
                     (N201)? mem[318] : 
                     (N203)? mem[333] : 
                     (N205)? mem[348] : 
                     (N207)? mem[363] : 
                     (N209)? mem[378] : 
                     (N211)? mem[393] : 
                     (N213)? mem[408] : 
                     (N215)? mem[423] : 
                     (N217)? mem[438] : 
                     (N219)? mem[453] : 
                     (N221)? mem[468] : 
                     (N223)? mem[483] : 
                     (N225)? mem[498] : 
                     (N227)? mem[513] : 
                     (N229)? mem[528] : 
                     (N231)? mem[543] : 
                     (N233)? mem[558] : 
                     (N235)? mem[573] : 
                     (N237)? mem[588] : 
                     (N239)? mem[603] : 
                     (N241)? mem[618] : 
                     (N243)? mem[633] : 
                     (N245)? mem[648] : 
                     (N247)? mem[663] : 
                     (N249)? mem[678] : 
                     (N251)? mem[693] : 
                     (N253)? mem[708] : 
                     (N255)? mem[723] : 
                     (N257)? mem[738] : 
                     (N259)? mem[753] : 
                     (N261)? mem[768] : 
                     (N263)? mem[783] : 
                     (N265)? mem[798] : 
                     (N267)? mem[813] : 
                     (N269)? mem[828] : 
                     (N271)? mem[843] : 
                     (N273)? mem[858] : 
                     (N275)? mem[873] : 
                     (N277)? mem[888] : 
                     (N279)? mem[903] : 
                     (N281)? mem[918] : 
                     (N283)? mem[933] : 
                     (N285)? mem[948] : 
                     (N160)? mem[963] : 
                     (N162)? mem[978] : 
                     (N164)? mem[993] : 
                     (N166)? mem[1008] : 
                     (N168)? mem[1023] : 
                     (N170)? mem[1038] : 
                     (N172)? mem[1053] : 
                     (N174)? mem[1068] : 
                     (N176)? mem[1083] : 
                     (N178)? mem[1098] : 
                     (N180)? mem[1113] : 
                     (N182)? mem[1128] : 
                     (N184)? mem[1143] : 
                     (N186)? mem[1158] : 
                     (N188)? mem[1173] : 
                     (N190)? mem[1188] : 
                     (N192)? mem[1203] : 
                     (N194)? mem[1218] : 
                     (N196)? mem[1233] : 
                     (N198)? mem[1248] : 
                     (N200)? mem[1263] : 
                     (N202)? mem[1278] : 
                     (N204)? mem[1293] : 
                     (N206)? mem[1308] : 
                     (N208)? mem[1323] : 
                     (N210)? mem[1338] : 
                     (N212)? mem[1353] : 
                     (N214)? mem[1368] : 
                     (N216)? mem[1383] : 
                     (N218)? mem[1398] : 
                     (N220)? mem[1413] : 
                     (N222)? mem[1428] : 
                     (N224)? mem[1443] : 
                     (N226)? mem[1458] : 
                     (N228)? mem[1473] : 
                     (N230)? mem[1488] : 
                     (N232)? mem[1503] : 
                     (N234)? mem[1518] : 
                     (N236)? mem[1533] : 
                     (N238)? mem[1548] : 
                     (N240)? mem[1563] : 
                     (N242)? mem[1578] : 
                     (N244)? mem[1593] : 
                     (N246)? mem[1608] : 
                     (N248)? mem[1623] : 
                     (N250)? mem[1638] : 
                     (N252)? mem[1653] : 
                     (N254)? mem[1668] : 
                     (N256)? mem[1683] : 
                     (N258)? mem[1698] : 
                     (N260)? mem[1713] : 
                     (N262)? mem[1728] : 
                     (N264)? mem[1743] : 
                     (N266)? mem[1758] : 
                     (N268)? mem[1773] : 
                     (N270)? mem[1788] : 
                     (N272)? mem[1803] : 
                     (N274)? mem[1818] : 
                     (N276)? mem[1833] : 
                     (N278)? mem[1848] : 
                     (N280)? mem[1863] : 
                     (N282)? mem[1878] : 
                     (N284)? mem[1893] : 
                     (N286)? mem[1908] : 1'b0;
  assign data_o[2] = (N159)? mem[2] : 
                     (N161)? mem[17] : 
                     (N163)? mem[32] : 
                     (N165)? mem[47] : 
                     (N167)? mem[62] : 
                     (N169)? mem[77] : 
                     (N171)? mem[92] : 
                     (N173)? mem[107] : 
                     (N175)? mem[122] : 
                     (N177)? mem[137] : 
                     (N179)? mem[152] : 
                     (N181)? mem[167] : 
                     (N183)? mem[182] : 
                     (N185)? mem[197] : 
                     (N187)? mem[212] : 
                     (N189)? mem[227] : 
                     (N191)? mem[242] : 
                     (N193)? mem[257] : 
                     (N195)? mem[272] : 
                     (N197)? mem[287] : 
                     (N199)? mem[302] : 
                     (N201)? mem[317] : 
                     (N203)? mem[332] : 
                     (N205)? mem[347] : 
                     (N207)? mem[362] : 
                     (N209)? mem[377] : 
                     (N211)? mem[392] : 
                     (N213)? mem[407] : 
                     (N215)? mem[422] : 
                     (N217)? mem[437] : 
                     (N219)? mem[452] : 
                     (N221)? mem[467] : 
                     (N223)? mem[482] : 
                     (N225)? mem[497] : 
                     (N227)? mem[512] : 
                     (N229)? mem[527] : 
                     (N231)? mem[542] : 
                     (N233)? mem[557] : 
                     (N235)? mem[572] : 
                     (N237)? mem[587] : 
                     (N239)? mem[602] : 
                     (N241)? mem[617] : 
                     (N243)? mem[632] : 
                     (N245)? mem[647] : 
                     (N247)? mem[662] : 
                     (N249)? mem[677] : 
                     (N251)? mem[692] : 
                     (N253)? mem[707] : 
                     (N255)? mem[722] : 
                     (N257)? mem[737] : 
                     (N259)? mem[752] : 
                     (N261)? mem[767] : 
                     (N263)? mem[782] : 
                     (N265)? mem[797] : 
                     (N267)? mem[812] : 
                     (N269)? mem[827] : 
                     (N271)? mem[842] : 
                     (N273)? mem[857] : 
                     (N275)? mem[872] : 
                     (N277)? mem[887] : 
                     (N279)? mem[902] : 
                     (N281)? mem[917] : 
                     (N283)? mem[932] : 
                     (N285)? mem[947] : 
                     (N160)? mem[962] : 
                     (N162)? mem[977] : 
                     (N164)? mem[992] : 
                     (N166)? mem[1007] : 
                     (N168)? mem[1022] : 
                     (N170)? mem[1037] : 
                     (N172)? mem[1052] : 
                     (N174)? mem[1067] : 
                     (N176)? mem[1082] : 
                     (N178)? mem[1097] : 
                     (N180)? mem[1112] : 
                     (N182)? mem[1127] : 
                     (N184)? mem[1142] : 
                     (N186)? mem[1157] : 
                     (N188)? mem[1172] : 
                     (N190)? mem[1187] : 
                     (N192)? mem[1202] : 
                     (N194)? mem[1217] : 
                     (N196)? mem[1232] : 
                     (N198)? mem[1247] : 
                     (N200)? mem[1262] : 
                     (N202)? mem[1277] : 
                     (N204)? mem[1292] : 
                     (N206)? mem[1307] : 
                     (N208)? mem[1322] : 
                     (N210)? mem[1337] : 
                     (N212)? mem[1352] : 
                     (N214)? mem[1367] : 
                     (N216)? mem[1382] : 
                     (N218)? mem[1397] : 
                     (N220)? mem[1412] : 
                     (N222)? mem[1427] : 
                     (N224)? mem[1442] : 
                     (N226)? mem[1457] : 
                     (N228)? mem[1472] : 
                     (N230)? mem[1487] : 
                     (N232)? mem[1502] : 
                     (N234)? mem[1517] : 
                     (N236)? mem[1532] : 
                     (N238)? mem[1547] : 
                     (N240)? mem[1562] : 
                     (N242)? mem[1577] : 
                     (N244)? mem[1592] : 
                     (N246)? mem[1607] : 
                     (N248)? mem[1622] : 
                     (N250)? mem[1637] : 
                     (N252)? mem[1652] : 
                     (N254)? mem[1667] : 
                     (N256)? mem[1682] : 
                     (N258)? mem[1697] : 
                     (N260)? mem[1712] : 
                     (N262)? mem[1727] : 
                     (N264)? mem[1742] : 
                     (N266)? mem[1757] : 
                     (N268)? mem[1772] : 
                     (N270)? mem[1787] : 
                     (N272)? mem[1802] : 
                     (N274)? mem[1817] : 
                     (N276)? mem[1832] : 
                     (N278)? mem[1847] : 
                     (N280)? mem[1862] : 
                     (N282)? mem[1877] : 
                     (N284)? mem[1892] : 
                     (N286)? mem[1907] : 1'b0;
  assign data_o[1] = (N159)? mem[1] : 
                     (N161)? mem[16] : 
                     (N163)? mem[31] : 
                     (N165)? mem[46] : 
                     (N167)? mem[61] : 
                     (N169)? mem[76] : 
                     (N171)? mem[91] : 
                     (N173)? mem[106] : 
                     (N175)? mem[121] : 
                     (N177)? mem[136] : 
                     (N179)? mem[151] : 
                     (N181)? mem[166] : 
                     (N183)? mem[181] : 
                     (N185)? mem[196] : 
                     (N187)? mem[211] : 
                     (N189)? mem[226] : 
                     (N191)? mem[241] : 
                     (N193)? mem[256] : 
                     (N195)? mem[271] : 
                     (N197)? mem[286] : 
                     (N199)? mem[301] : 
                     (N201)? mem[316] : 
                     (N203)? mem[331] : 
                     (N205)? mem[346] : 
                     (N207)? mem[361] : 
                     (N209)? mem[376] : 
                     (N211)? mem[391] : 
                     (N213)? mem[406] : 
                     (N215)? mem[421] : 
                     (N217)? mem[436] : 
                     (N219)? mem[451] : 
                     (N221)? mem[466] : 
                     (N223)? mem[481] : 
                     (N225)? mem[496] : 
                     (N227)? mem[511] : 
                     (N229)? mem[526] : 
                     (N231)? mem[541] : 
                     (N233)? mem[556] : 
                     (N235)? mem[571] : 
                     (N237)? mem[586] : 
                     (N239)? mem[601] : 
                     (N241)? mem[616] : 
                     (N243)? mem[631] : 
                     (N245)? mem[646] : 
                     (N247)? mem[661] : 
                     (N249)? mem[676] : 
                     (N251)? mem[691] : 
                     (N253)? mem[706] : 
                     (N255)? mem[721] : 
                     (N257)? mem[736] : 
                     (N259)? mem[751] : 
                     (N261)? mem[766] : 
                     (N263)? mem[781] : 
                     (N265)? mem[796] : 
                     (N267)? mem[811] : 
                     (N269)? mem[826] : 
                     (N271)? mem[841] : 
                     (N273)? mem[856] : 
                     (N275)? mem[871] : 
                     (N277)? mem[886] : 
                     (N279)? mem[901] : 
                     (N281)? mem[916] : 
                     (N283)? mem[931] : 
                     (N285)? mem[946] : 
                     (N160)? mem[961] : 
                     (N162)? mem[976] : 
                     (N164)? mem[991] : 
                     (N166)? mem[1006] : 
                     (N168)? mem[1021] : 
                     (N170)? mem[1036] : 
                     (N172)? mem[1051] : 
                     (N174)? mem[1066] : 
                     (N176)? mem[1081] : 
                     (N178)? mem[1096] : 
                     (N180)? mem[1111] : 
                     (N182)? mem[1126] : 
                     (N184)? mem[1141] : 
                     (N186)? mem[1156] : 
                     (N188)? mem[1171] : 
                     (N190)? mem[1186] : 
                     (N192)? mem[1201] : 
                     (N194)? mem[1216] : 
                     (N196)? mem[1231] : 
                     (N198)? mem[1246] : 
                     (N200)? mem[1261] : 
                     (N202)? mem[1276] : 
                     (N204)? mem[1291] : 
                     (N206)? mem[1306] : 
                     (N208)? mem[1321] : 
                     (N210)? mem[1336] : 
                     (N212)? mem[1351] : 
                     (N214)? mem[1366] : 
                     (N216)? mem[1381] : 
                     (N218)? mem[1396] : 
                     (N220)? mem[1411] : 
                     (N222)? mem[1426] : 
                     (N224)? mem[1441] : 
                     (N226)? mem[1456] : 
                     (N228)? mem[1471] : 
                     (N230)? mem[1486] : 
                     (N232)? mem[1501] : 
                     (N234)? mem[1516] : 
                     (N236)? mem[1531] : 
                     (N238)? mem[1546] : 
                     (N240)? mem[1561] : 
                     (N242)? mem[1576] : 
                     (N244)? mem[1591] : 
                     (N246)? mem[1606] : 
                     (N248)? mem[1621] : 
                     (N250)? mem[1636] : 
                     (N252)? mem[1651] : 
                     (N254)? mem[1666] : 
                     (N256)? mem[1681] : 
                     (N258)? mem[1696] : 
                     (N260)? mem[1711] : 
                     (N262)? mem[1726] : 
                     (N264)? mem[1741] : 
                     (N266)? mem[1756] : 
                     (N268)? mem[1771] : 
                     (N270)? mem[1786] : 
                     (N272)? mem[1801] : 
                     (N274)? mem[1816] : 
                     (N276)? mem[1831] : 
                     (N278)? mem[1846] : 
                     (N280)? mem[1861] : 
                     (N282)? mem[1876] : 
                     (N284)? mem[1891] : 
                     (N286)? mem[1906] : 1'b0;
  assign data_o[0] = (N159)? mem[0] : 
                     (N161)? mem[15] : 
                     (N163)? mem[30] : 
                     (N165)? mem[45] : 
                     (N167)? mem[60] : 
                     (N169)? mem[75] : 
                     (N171)? mem[90] : 
                     (N173)? mem[105] : 
                     (N175)? mem[120] : 
                     (N177)? mem[135] : 
                     (N179)? mem[150] : 
                     (N181)? mem[165] : 
                     (N183)? mem[180] : 
                     (N185)? mem[195] : 
                     (N187)? mem[210] : 
                     (N189)? mem[225] : 
                     (N191)? mem[240] : 
                     (N193)? mem[255] : 
                     (N195)? mem[270] : 
                     (N197)? mem[285] : 
                     (N199)? mem[300] : 
                     (N201)? mem[315] : 
                     (N203)? mem[330] : 
                     (N205)? mem[345] : 
                     (N207)? mem[360] : 
                     (N209)? mem[375] : 
                     (N211)? mem[390] : 
                     (N213)? mem[405] : 
                     (N215)? mem[420] : 
                     (N217)? mem[435] : 
                     (N219)? mem[450] : 
                     (N221)? mem[465] : 
                     (N223)? mem[480] : 
                     (N225)? mem[495] : 
                     (N227)? mem[510] : 
                     (N229)? mem[525] : 
                     (N231)? mem[540] : 
                     (N233)? mem[555] : 
                     (N235)? mem[570] : 
                     (N237)? mem[585] : 
                     (N239)? mem[600] : 
                     (N241)? mem[615] : 
                     (N243)? mem[630] : 
                     (N245)? mem[645] : 
                     (N247)? mem[660] : 
                     (N249)? mem[675] : 
                     (N251)? mem[690] : 
                     (N253)? mem[705] : 
                     (N255)? mem[720] : 
                     (N257)? mem[735] : 
                     (N259)? mem[750] : 
                     (N261)? mem[765] : 
                     (N263)? mem[780] : 
                     (N265)? mem[795] : 
                     (N267)? mem[810] : 
                     (N269)? mem[825] : 
                     (N271)? mem[840] : 
                     (N273)? mem[855] : 
                     (N275)? mem[870] : 
                     (N277)? mem[885] : 
                     (N279)? mem[900] : 
                     (N281)? mem[915] : 
                     (N283)? mem[930] : 
                     (N285)? mem[945] : 
                     (N160)? mem[960] : 
                     (N162)? mem[975] : 
                     (N164)? mem[990] : 
                     (N166)? mem[1005] : 
                     (N168)? mem[1020] : 
                     (N170)? mem[1035] : 
                     (N172)? mem[1050] : 
                     (N174)? mem[1065] : 
                     (N176)? mem[1080] : 
                     (N178)? mem[1095] : 
                     (N180)? mem[1110] : 
                     (N182)? mem[1125] : 
                     (N184)? mem[1140] : 
                     (N186)? mem[1155] : 
                     (N188)? mem[1170] : 
                     (N190)? mem[1185] : 
                     (N192)? mem[1200] : 
                     (N194)? mem[1215] : 
                     (N196)? mem[1230] : 
                     (N198)? mem[1245] : 
                     (N200)? mem[1260] : 
                     (N202)? mem[1275] : 
                     (N204)? mem[1290] : 
                     (N206)? mem[1305] : 
                     (N208)? mem[1320] : 
                     (N210)? mem[1335] : 
                     (N212)? mem[1350] : 
                     (N214)? mem[1365] : 
                     (N216)? mem[1380] : 
                     (N218)? mem[1395] : 
                     (N220)? mem[1410] : 
                     (N222)? mem[1425] : 
                     (N224)? mem[1440] : 
                     (N226)? mem[1455] : 
                     (N228)? mem[1470] : 
                     (N230)? mem[1485] : 
                     (N232)? mem[1500] : 
                     (N234)? mem[1515] : 
                     (N236)? mem[1530] : 
                     (N238)? mem[1545] : 
                     (N240)? mem[1560] : 
                     (N242)? mem[1575] : 
                     (N244)? mem[1590] : 
                     (N246)? mem[1605] : 
                     (N248)? mem[1620] : 
                     (N250)? mem[1635] : 
                     (N252)? mem[1650] : 
                     (N254)? mem[1665] : 
                     (N256)? mem[1680] : 
                     (N258)? mem[1695] : 
                     (N260)? mem[1710] : 
                     (N262)? mem[1725] : 
                     (N264)? mem[1740] : 
                     (N266)? mem[1755] : 
                     (N268)? mem[1770] : 
                     (N270)? mem[1785] : 
                     (N272)? mem[1800] : 
                     (N274)? mem[1815] : 
                     (N276)? mem[1830] : 
                     (N278)? mem[1845] : 
                     (N280)? mem[1860] : 
                     (N282)? mem[1875] : 
                     (N284)? mem[1890] : 
                     (N286)? mem[1905] : 1'b0;

  always @(posedge clk_i) begin
    if(N4735) begin
      mem_1919_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4734) begin
      mem_1918_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4733) begin
      mem_1917_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4732) begin
      mem_1916_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4731) begin
      mem_1915_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4730) begin
      mem_1914_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4729) begin
      mem_1913_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4728) begin
      mem_1912_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4727) begin
      mem_1911_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4726) begin
      mem_1910_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4725) begin
      mem_1909_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4724) begin
      mem_1908_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4723) begin
      mem_1907_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4722) begin
      mem_1906_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4721) begin
      mem_1905_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4720) begin
      mem_1904_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4719) begin
      mem_1903_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4718) begin
      mem_1902_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4717) begin
      mem_1901_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4716) begin
      mem_1900_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4715) begin
      mem_1899_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4714) begin
      mem_1898_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4713) begin
      mem_1897_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4712) begin
      mem_1896_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4711) begin
      mem_1895_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4710) begin
      mem_1894_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4709) begin
      mem_1893_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4708) begin
      mem_1892_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4707) begin
      mem_1891_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4706) begin
      mem_1890_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4705) begin
      mem_1889_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4704) begin
      mem_1888_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4703) begin
      mem_1887_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4702) begin
      mem_1886_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4701) begin
      mem_1885_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4700) begin
      mem_1884_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4699) begin
      mem_1883_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4698) begin
      mem_1882_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4697) begin
      mem_1881_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4696) begin
      mem_1880_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4695) begin
      mem_1879_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4694) begin
      mem_1878_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4693) begin
      mem_1877_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4692) begin
      mem_1876_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4691) begin
      mem_1875_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4690) begin
      mem_1874_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4689) begin
      mem_1873_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4688) begin
      mem_1872_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4687) begin
      mem_1871_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4686) begin
      mem_1870_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4685) begin
      mem_1869_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4684) begin
      mem_1868_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4683) begin
      mem_1867_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4682) begin
      mem_1866_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4681) begin
      mem_1865_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4680) begin
      mem_1864_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4679) begin
      mem_1863_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4678) begin
      mem_1862_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4677) begin
      mem_1861_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4676) begin
      mem_1860_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4675) begin
      mem_1859_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4674) begin
      mem_1858_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4673) begin
      mem_1857_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4672) begin
      mem_1856_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4671) begin
      mem_1855_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4670) begin
      mem_1854_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4669) begin
      mem_1853_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4668) begin
      mem_1852_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4667) begin
      mem_1851_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4666) begin
      mem_1850_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4665) begin
      mem_1849_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4664) begin
      mem_1848_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4663) begin
      mem_1847_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4662) begin
      mem_1846_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4661) begin
      mem_1845_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4660) begin
      mem_1844_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4659) begin
      mem_1843_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4658) begin
      mem_1842_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4657) begin
      mem_1841_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4656) begin
      mem_1840_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4655) begin
      mem_1839_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4654) begin
      mem_1838_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4653) begin
      mem_1837_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4652) begin
      mem_1836_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4651) begin
      mem_1835_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4650) begin
      mem_1834_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4649) begin
      mem_1833_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4648) begin
      mem_1832_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4647) begin
      mem_1831_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4646) begin
      mem_1830_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4645) begin
      mem_1829_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4644) begin
      mem_1828_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4643) begin
      mem_1827_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4642) begin
      mem_1826_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4641) begin
      mem_1825_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4640) begin
      mem_1824_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4639) begin
      mem_1823_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4638) begin
      mem_1822_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4637) begin
      mem_1821_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4636) begin
      mem_1820_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4635) begin
      mem_1819_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4634) begin
      mem_1818_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4633) begin
      mem_1817_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4632) begin
      mem_1816_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4631) begin
      mem_1815_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4630) begin
      mem_1814_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4629) begin
      mem_1813_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4628) begin
      mem_1812_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4627) begin
      mem_1811_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4626) begin
      mem_1810_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4625) begin
      mem_1809_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4624) begin
      mem_1808_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4623) begin
      mem_1807_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4622) begin
      mem_1806_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4621) begin
      mem_1805_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4620) begin
      mem_1804_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4619) begin
      mem_1803_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4618) begin
      mem_1802_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4617) begin
      mem_1801_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4616) begin
      mem_1800_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4615) begin
      mem_1799_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4614) begin
      mem_1798_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4613) begin
      mem_1797_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4612) begin
      mem_1796_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4611) begin
      mem_1795_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4610) begin
      mem_1794_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4609) begin
      mem_1793_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4608) begin
      mem_1792_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4607) begin
      mem_1791_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4606) begin
      mem_1790_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4605) begin
      mem_1789_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4604) begin
      mem_1788_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4603) begin
      mem_1787_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4602) begin
      mem_1786_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4601) begin
      mem_1785_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4600) begin
      mem_1784_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4599) begin
      mem_1783_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4598) begin
      mem_1782_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4597) begin
      mem_1781_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4596) begin
      mem_1780_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4595) begin
      mem_1779_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4594) begin
      mem_1778_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4593) begin
      mem_1777_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4592) begin
      mem_1776_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4591) begin
      mem_1775_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4590) begin
      mem_1774_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4589) begin
      mem_1773_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4588) begin
      mem_1772_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4587) begin
      mem_1771_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4586) begin
      mem_1770_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4585) begin
      mem_1769_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4584) begin
      mem_1768_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4583) begin
      mem_1767_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4582) begin
      mem_1766_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4581) begin
      mem_1765_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4580) begin
      mem_1764_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4579) begin
      mem_1763_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4578) begin
      mem_1762_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4577) begin
      mem_1761_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4576) begin
      mem_1760_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4575) begin
      mem_1759_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4574) begin
      mem_1758_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4573) begin
      mem_1757_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4572) begin
      mem_1756_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4571) begin
      mem_1755_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4570) begin
      mem_1754_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4569) begin
      mem_1753_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4568) begin
      mem_1752_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4567) begin
      mem_1751_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4566) begin
      mem_1750_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4565) begin
      mem_1749_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4564) begin
      mem_1748_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4563) begin
      mem_1747_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4562) begin
      mem_1746_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4561) begin
      mem_1745_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4560) begin
      mem_1744_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4559) begin
      mem_1743_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4558) begin
      mem_1742_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4557) begin
      mem_1741_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4556) begin
      mem_1740_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4555) begin
      mem_1739_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4554) begin
      mem_1738_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4553) begin
      mem_1737_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4552) begin
      mem_1736_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4551) begin
      mem_1735_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4550) begin
      mem_1734_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4549) begin
      mem_1733_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4548) begin
      mem_1732_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4547) begin
      mem_1731_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4546) begin
      mem_1730_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4545) begin
      mem_1729_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4544) begin
      mem_1728_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4543) begin
      mem_1727_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4542) begin
      mem_1726_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4541) begin
      mem_1725_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4540) begin
      mem_1724_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4539) begin
      mem_1723_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4538) begin
      mem_1722_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4537) begin
      mem_1721_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4536) begin
      mem_1720_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4535) begin
      mem_1719_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4534) begin
      mem_1718_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4533) begin
      mem_1717_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4532) begin
      mem_1716_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4531) begin
      mem_1715_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4530) begin
      mem_1714_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4529) begin
      mem_1713_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4528) begin
      mem_1712_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4527) begin
      mem_1711_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4526) begin
      mem_1710_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4525) begin
      mem_1709_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4524) begin
      mem_1708_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4523) begin
      mem_1707_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4522) begin
      mem_1706_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4521) begin
      mem_1705_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4520) begin
      mem_1704_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4519) begin
      mem_1703_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4518) begin
      mem_1702_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4517) begin
      mem_1701_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4516) begin
      mem_1700_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4515) begin
      mem_1699_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4514) begin
      mem_1698_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4513) begin
      mem_1697_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4512) begin
      mem_1696_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4511) begin
      mem_1695_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4510) begin
      mem_1694_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4509) begin
      mem_1693_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4508) begin
      mem_1692_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4507) begin
      mem_1691_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4506) begin
      mem_1690_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4505) begin
      mem_1689_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4504) begin
      mem_1688_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4503) begin
      mem_1687_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4502) begin
      mem_1686_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4501) begin
      mem_1685_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4500) begin
      mem_1684_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4499) begin
      mem_1683_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4498) begin
      mem_1682_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4497) begin
      mem_1681_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4496) begin
      mem_1680_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4495) begin
      mem_1679_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4494) begin
      mem_1678_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4493) begin
      mem_1677_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4492) begin
      mem_1676_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4491) begin
      mem_1675_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4490) begin
      mem_1674_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4489) begin
      mem_1673_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4488) begin
      mem_1672_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4487) begin
      mem_1671_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4486) begin
      mem_1670_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4485) begin
      mem_1669_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4484) begin
      mem_1668_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4483) begin
      mem_1667_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4482) begin
      mem_1666_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4481) begin
      mem_1665_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4480) begin
      mem_1664_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4479) begin
      mem_1663_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4478) begin
      mem_1662_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4477) begin
      mem_1661_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4476) begin
      mem_1660_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4475) begin
      mem_1659_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4474) begin
      mem_1658_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4473) begin
      mem_1657_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4472) begin
      mem_1656_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4471) begin
      mem_1655_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4470) begin
      mem_1654_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4469) begin
      mem_1653_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4468) begin
      mem_1652_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4467) begin
      mem_1651_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4466) begin
      mem_1650_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4465) begin
      mem_1649_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4464) begin
      mem_1648_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4463) begin
      mem_1647_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4462) begin
      mem_1646_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4461) begin
      mem_1645_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4460) begin
      mem_1644_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4459) begin
      mem_1643_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4458) begin
      mem_1642_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4457) begin
      mem_1641_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4456) begin
      mem_1640_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4455) begin
      mem_1639_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4454) begin
      mem_1638_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4453) begin
      mem_1637_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4452) begin
      mem_1636_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4451) begin
      mem_1635_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4450) begin
      mem_1634_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4449) begin
      mem_1633_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4448) begin
      mem_1632_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4447) begin
      mem_1631_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4446) begin
      mem_1630_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4445) begin
      mem_1629_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4444) begin
      mem_1628_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4443) begin
      mem_1627_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4442) begin
      mem_1626_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4441) begin
      mem_1625_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4440) begin
      mem_1624_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4439) begin
      mem_1623_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4438) begin
      mem_1622_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4437) begin
      mem_1621_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4436) begin
      mem_1620_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4435) begin
      mem_1619_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4434) begin
      mem_1618_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4433) begin
      mem_1617_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4432) begin
      mem_1616_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4431) begin
      mem_1615_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4430) begin
      mem_1614_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4429) begin
      mem_1613_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4428) begin
      mem_1612_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4427) begin
      mem_1611_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4426) begin
      mem_1610_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4425) begin
      mem_1609_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4424) begin
      mem_1608_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4423) begin
      mem_1607_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4422) begin
      mem_1606_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4421) begin
      mem_1605_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4420) begin
      mem_1604_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4419) begin
      mem_1603_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4418) begin
      mem_1602_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4417) begin
      mem_1601_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4416) begin
      mem_1600_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4415) begin
      mem_1599_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4414) begin
      mem_1598_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4413) begin
      mem_1597_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4412) begin
      mem_1596_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4411) begin
      mem_1595_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4410) begin
      mem_1594_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4409) begin
      mem_1593_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4408) begin
      mem_1592_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4407) begin
      mem_1591_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4406) begin
      mem_1590_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4405) begin
      mem_1589_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4404) begin
      mem_1588_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4403) begin
      mem_1587_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4402) begin
      mem_1586_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4401) begin
      mem_1585_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4400) begin
      mem_1584_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4399) begin
      mem_1583_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4398) begin
      mem_1582_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4397) begin
      mem_1581_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4396) begin
      mem_1580_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4395) begin
      mem_1579_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4394) begin
      mem_1578_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4393) begin
      mem_1577_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4392) begin
      mem_1576_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4391) begin
      mem_1575_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4390) begin
      mem_1574_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4389) begin
      mem_1573_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4388) begin
      mem_1572_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4387) begin
      mem_1571_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4386) begin
      mem_1570_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4385) begin
      mem_1569_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4384) begin
      mem_1568_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4383) begin
      mem_1567_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4382) begin
      mem_1566_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4381) begin
      mem_1565_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4380) begin
      mem_1564_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4379) begin
      mem_1563_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4378) begin
      mem_1562_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4377) begin
      mem_1561_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4376) begin
      mem_1560_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4375) begin
      mem_1559_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4374) begin
      mem_1558_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4373) begin
      mem_1557_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4372) begin
      mem_1556_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4371) begin
      mem_1555_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4370) begin
      mem_1554_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4369) begin
      mem_1553_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4368) begin
      mem_1552_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4367) begin
      mem_1551_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4366) begin
      mem_1550_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4365) begin
      mem_1549_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4364) begin
      mem_1548_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4363) begin
      mem_1547_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4362) begin
      mem_1546_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4361) begin
      mem_1545_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4360) begin
      mem_1544_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4359) begin
      mem_1543_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4358) begin
      mem_1542_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4357) begin
      mem_1541_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4356) begin
      mem_1540_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4355) begin
      mem_1539_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4354) begin
      mem_1538_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4353) begin
      mem_1537_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4352) begin
      mem_1536_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4351) begin
      mem_1535_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4350) begin
      mem_1534_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4349) begin
      mem_1533_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4348) begin
      mem_1532_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4347) begin
      mem_1531_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4346) begin
      mem_1530_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4345) begin
      mem_1529_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4344) begin
      mem_1528_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4343) begin
      mem_1527_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4342) begin
      mem_1526_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4341) begin
      mem_1525_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4340) begin
      mem_1524_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4339) begin
      mem_1523_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4338) begin
      mem_1522_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4337) begin
      mem_1521_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4336) begin
      mem_1520_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4335) begin
      mem_1519_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4334) begin
      mem_1518_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4333) begin
      mem_1517_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4332) begin
      mem_1516_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4331) begin
      mem_1515_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4330) begin
      mem_1514_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4329) begin
      mem_1513_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4328) begin
      mem_1512_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4327) begin
      mem_1511_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4326) begin
      mem_1510_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4325) begin
      mem_1509_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4324) begin
      mem_1508_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4323) begin
      mem_1507_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4322) begin
      mem_1506_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4321) begin
      mem_1505_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4320) begin
      mem_1504_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4319) begin
      mem_1503_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4318) begin
      mem_1502_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4317) begin
      mem_1501_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4316) begin
      mem_1500_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4315) begin
      mem_1499_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4314) begin
      mem_1498_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4313) begin
      mem_1497_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4312) begin
      mem_1496_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4311) begin
      mem_1495_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4310) begin
      mem_1494_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4309) begin
      mem_1493_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4308) begin
      mem_1492_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4307) begin
      mem_1491_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4306) begin
      mem_1490_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4305) begin
      mem_1489_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4304) begin
      mem_1488_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4303) begin
      mem_1487_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4302) begin
      mem_1486_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4301) begin
      mem_1485_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4300) begin
      mem_1484_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4299) begin
      mem_1483_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4298) begin
      mem_1482_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4297) begin
      mem_1481_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4296) begin
      mem_1480_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4295) begin
      mem_1479_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4294) begin
      mem_1478_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4293) begin
      mem_1477_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4292) begin
      mem_1476_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4291) begin
      mem_1475_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4290) begin
      mem_1474_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4289) begin
      mem_1473_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4288) begin
      mem_1472_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4287) begin
      mem_1471_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4286) begin
      mem_1470_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4285) begin
      mem_1469_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4284) begin
      mem_1468_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4283) begin
      mem_1467_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4282) begin
      mem_1466_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4281) begin
      mem_1465_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4280) begin
      mem_1464_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4279) begin
      mem_1463_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4278) begin
      mem_1462_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4277) begin
      mem_1461_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4276) begin
      mem_1460_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4275) begin
      mem_1459_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4274) begin
      mem_1458_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4273) begin
      mem_1457_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4272) begin
      mem_1456_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4271) begin
      mem_1455_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4270) begin
      mem_1454_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4269) begin
      mem_1453_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4268) begin
      mem_1452_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4267) begin
      mem_1451_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4266) begin
      mem_1450_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4265) begin
      mem_1449_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4264) begin
      mem_1448_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4263) begin
      mem_1447_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4262) begin
      mem_1446_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4261) begin
      mem_1445_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4260) begin
      mem_1444_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4259) begin
      mem_1443_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4258) begin
      mem_1442_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4257) begin
      mem_1441_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4256) begin
      mem_1440_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4255) begin
      mem_1439_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4254) begin
      mem_1438_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4253) begin
      mem_1437_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4252) begin
      mem_1436_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4251) begin
      mem_1435_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4250) begin
      mem_1434_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4249) begin
      mem_1433_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4248) begin
      mem_1432_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4247) begin
      mem_1431_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4246) begin
      mem_1430_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4245) begin
      mem_1429_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4244) begin
      mem_1428_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4243) begin
      mem_1427_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4242) begin
      mem_1426_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4241) begin
      mem_1425_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4240) begin
      mem_1424_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4239) begin
      mem_1423_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4238) begin
      mem_1422_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4237) begin
      mem_1421_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4236) begin
      mem_1420_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4235) begin
      mem_1419_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4234) begin
      mem_1418_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4233) begin
      mem_1417_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4232) begin
      mem_1416_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4231) begin
      mem_1415_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4230) begin
      mem_1414_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4229) begin
      mem_1413_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4228) begin
      mem_1412_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4227) begin
      mem_1411_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4226) begin
      mem_1410_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4225) begin
      mem_1409_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4224) begin
      mem_1408_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4223) begin
      mem_1407_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4222) begin
      mem_1406_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4221) begin
      mem_1405_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4220) begin
      mem_1404_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4219) begin
      mem_1403_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4218) begin
      mem_1402_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4217) begin
      mem_1401_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4216) begin
      mem_1400_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4215) begin
      mem_1399_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4214) begin
      mem_1398_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4213) begin
      mem_1397_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4212) begin
      mem_1396_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4211) begin
      mem_1395_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4210) begin
      mem_1394_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4209) begin
      mem_1393_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4208) begin
      mem_1392_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4207) begin
      mem_1391_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4206) begin
      mem_1390_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4205) begin
      mem_1389_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4204) begin
      mem_1388_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4203) begin
      mem_1387_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4202) begin
      mem_1386_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4201) begin
      mem_1385_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4200) begin
      mem_1384_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4199) begin
      mem_1383_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4198) begin
      mem_1382_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4197) begin
      mem_1381_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4196) begin
      mem_1380_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4195) begin
      mem_1379_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4194) begin
      mem_1378_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4193) begin
      mem_1377_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4192) begin
      mem_1376_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4191) begin
      mem_1375_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4190) begin
      mem_1374_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4189) begin
      mem_1373_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4188) begin
      mem_1372_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4187) begin
      mem_1371_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4186) begin
      mem_1370_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4185) begin
      mem_1369_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4184) begin
      mem_1368_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4183) begin
      mem_1367_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4182) begin
      mem_1366_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4181) begin
      mem_1365_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4180) begin
      mem_1364_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4179) begin
      mem_1363_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4178) begin
      mem_1362_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4177) begin
      mem_1361_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4176) begin
      mem_1360_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4175) begin
      mem_1359_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4174) begin
      mem_1358_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4173) begin
      mem_1357_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4172) begin
      mem_1356_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4171) begin
      mem_1355_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4170) begin
      mem_1354_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4169) begin
      mem_1353_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4168) begin
      mem_1352_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4167) begin
      mem_1351_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4166) begin
      mem_1350_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4165) begin
      mem_1349_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4164) begin
      mem_1348_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4163) begin
      mem_1347_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4162) begin
      mem_1346_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4161) begin
      mem_1345_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4160) begin
      mem_1344_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4159) begin
      mem_1343_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4158) begin
      mem_1342_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4157) begin
      mem_1341_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4156) begin
      mem_1340_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4155) begin
      mem_1339_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4154) begin
      mem_1338_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4153) begin
      mem_1337_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4152) begin
      mem_1336_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4151) begin
      mem_1335_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4150) begin
      mem_1334_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4149) begin
      mem_1333_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4148) begin
      mem_1332_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4147) begin
      mem_1331_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4146) begin
      mem_1330_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4145) begin
      mem_1329_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4144) begin
      mem_1328_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4143) begin
      mem_1327_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4142) begin
      mem_1326_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4141) begin
      mem_1325_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4140) begin
      mem_1324_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4139) begin
      mem_1323_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4138) begin
      mem_1322_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4137) begin
      mem_1321_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4136) begin
      mem_1320_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4135) begin
      mem_1319_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4134) begin
      mem_1318_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4133) begin
      mem_1317_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4132) begin
      mem_1316_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4131) begin
      mem_1315_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4130) begin
      mem_1314_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4129) begin
      mem_1313_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4128) begin
      mem_1312_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4127) begin
      mem_1311_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4126) begin
      mem_1310_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4125) begin
      mem_1309_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4124) begin
      mem_1308_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4123) begin
      mem_1307_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4122) begin
      mem_1306_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4121) begin
      mem_1305_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4120) begin
      mem_1304_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4119) begin
      mem_1303_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4118) begin
      mem_1302_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4117) begin
      mem_1301_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4116) begin
      mem_1300_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4115) begin
      mem_1299_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4114) begin
      mem_1298_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4113) begin
      mem_1297_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4112) begin
      mem_1296_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4111) begin
      mem_1295_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4110) begin
      mem_1294_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4109) begin
      mem_1293_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4108) begin
      mem_1292_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4107) begin
      mem_1291_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4106) begin
      mem_1290_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4105) begin
      mem_1289_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4104) begin
      mem_1288_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4103) begin
      mem_1287_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4102) begin
      mem_1286_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4101) begin
      mem_1285_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4100) begin
      mem_1284_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4099) begin
      mem_1283_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4098) begin
      mem_1282_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4097) begin
      mem_1281_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4096) begin
      mem_1280_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4095) begin
      mem_1279_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4094) begin
      mem_1278_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4093) begin
      mem_1277_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4092) begin
      mem_1276_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4091) begin
      mem_1275_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4090) begin
      mem_1274_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4089) begin
      mem_1273_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4088) begin
      mem_1272_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4087) begin
      mem_1271_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4086) begin
      mem_1270_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4085) begin
      mem_1269_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4084) begin
      mem_1268_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4083) begin
      mem_1267_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4082) begin
      mem_1266_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4081) begin
      mem_1265_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4080) begin
      mem_1264_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4079) begin
      mem_1263_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4078) begin
      mem_1262_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4077) begin
      mem_1261_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4076) begin
      mem_1260_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4075) begin
      mem_1259_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4074) begin
      mem_1258_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4073) begin
      mem_1257_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4072) begin
      mem_1256_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4071) begin
      mem_1255_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4070) begin
      mem_1254_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4069) begin
      mem_1253_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4068) begin
      mem_1252_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4067) begin
      mem_1251_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4066) begin
      mem_1250_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4065) begin
      mem_1249_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4064) begin
      mem_1248_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4063) begin
      mem_1247_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4062) begin
      mem_1246_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4061) begin
      mem_1245_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4060) begin
      mem_1244_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4059) begin
      mem_1243_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4058) begin
      mem_1242_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4057) begin
      mem_1241_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4056) begin
      mem_1240_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4055) begin
      mem_1239_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4054) begin
      mem_1238_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4053) begin
      mem_1237_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4052) begin
      mem_1236_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4051) begin
      mem_1235_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4050) begin
      mem_1234_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4049) begin
      mem_1233_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4048) begin
      mem_1232_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4047) begin
      mem_1231_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4046) begin
      mem_1230_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4045) begin
      mem_1229_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4044) begin
      mem_1228_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4043) begin
      mem_1227_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4042) begin
      mem_1226_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4041) begin
      mem_1225_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4040) begin
      mem_1224_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4039) begin
      mem_1223_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4038) begin
      mem_1222_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4037) begin
      mem_1221_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4036) begin
      mem_1220_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4035) begin
      mem_1219_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4034) begin
      mem_1218_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4033) begin
      mem_1217_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4032) begin
      mem_1216_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4031) begin
      mem_1215_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4030) begin
      mem_1214_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4029) begin
      mem_1213_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4028) begin
      mem_1212_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4027) begin
      mem_1211_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4026) begin
      mem_1210_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4025) begin
      mem_1209_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4024) begin
      mem_1208_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4023) begin
      mem_1207_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4022) begin
      mem_1206_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4021) begin
      mem_1205_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4020) begin
      mem_1204_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4019) begin
      mem_1203_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4018) begin
      mem_1202_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4017) begin
      mem_1201_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4016) begin
      mem_1200_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4015) begin
      mem_1199_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N4014) begin
      mem_1198_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N4013) begin
      mem_1197_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N4012) begin
      mem_1196_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N4011) begin
      mem_1195_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N4010) begin
      mem_1194_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N4009) begin
      mem_1193_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N4008) begin
      mem_1192_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N4007) begin
      mem_1191_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N4006) begin
      mem_1190_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N4005) begin
      mem_1189_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N4004) begin
      mem_1188_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N4003) begin
      mem_1187_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N4002) begin
      mem_1186_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N4001) begin
      mem_1185_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N4000) begin
      mem_1184_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3999) begin
      mem_1183_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3998) begin
      mem_1182_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3997) begin
      mem_1181_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3996) begin
      mem_1180_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3995) begin
      mem_1179_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3994) begin
      mem_1178_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3993) begin
      mem_1177_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3992) begin
      mem_1176_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3991) begin
      mem_1175_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3990) begin
      mem_1174_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3989) begin
      mem_1173_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3988) begin
      mem_1172_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3987) begin
      mem_1171_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3986) begin
      mem_1170_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3985) begin
      mem_1169_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3984) begin
      mem_1168_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3983) begin
      mem_1167_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3982) begin
      mem_1166_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3981) begin
      mem_1165_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3980) begin
      mem_1164_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3979) begin
      mem_1163_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3978) begin
      mem_1162_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3977) begin
      mem_1161_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3976) begin
      mem_1160_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3975) begin
      mem_1159_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3974) begin
      mem_1158_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3973) begin
      mem_1157_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3972) begin
      mem_1156_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3971) begin
      mem_1155_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3970) begin
      mem_1154_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3969) begin
      mem_1153_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3968) begin
      mem_1152_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3967) begin
      mem_1151_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3966) begin
      mem_1150_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3965) begin
      mem_1149_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3964) begin
      mem_1148_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3963) begin
      mem_1147_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3962) begin
      mem_1146_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3961) begin
      mem_1145_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3960) begin
      mem_1144_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3959) begin
      mem_1143_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3958) begin
      mem_1142_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3957) begin
      mem_1141_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3956) begin
      mem_1140_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3955) begin
      mem_1139_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3954) begin
      mem_1138_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3953) begin
      mem_1137_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3952) begin
      mem_1136_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3951) begin
      mem_1135_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3950) begin
      mem_1134_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3949) begin
      mem_1133_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3948) begin
      mem_1132_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3947) begin
      mem_1131_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3946) begin
      mem_1130_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3945) begin
      mem_1129_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3944) begin
      mem_1128_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3943) begin
      mem_1127_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3942) begin
      mem_1126_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3941) begin
      mem_1125_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3940) begin
      mem_1124_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3939) begin
      mem_1123_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3938) begin
      mem_1122_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3937) begin
      mem_1121_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3936) begin
      mem_1120_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3935) begin
      mem_1119_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3934) begin
      mem_1118_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3933) begin
      mem_1117_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3932) begin
      mem_1116_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3931) begin
      mem_1115_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3930) begin
      mem_1114_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3929) begin
      mem_1113_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3928) begin
      mem_1112_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3927) begin
      mem_1111_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3926) begin
      mem_1110_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3925) begin
      mem_1109_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3924) begin
      mem_1108_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3923) begin
      mem_1107_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3922) begin
      mem_1106_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3921) begin
      mem_1105_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3920) begin
      mem_1104_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3919) begin
      mem_1103_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3918) begin
      mem_1102_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3917) begin
      mem_1101_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3916) begin
      mem_1100_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3915) begin
      mem_1099_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3914) begin
      mem_1098_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3913) begin
      mem_1097_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3912) begin
      mem_1096_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3911) begin
      mem_1095_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3910) begin
      mem_1094_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3909) begin
      mem_1093_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3908) begin
      mem_1092_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3907) begin
      mem_1091_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3906) begin
      mem_1090_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3905) begin
      mem_1089_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3904) begin
      mem_1088_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3903) begin
      mem_1087_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3902) begin
      mem_1086_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3901) begin
      mem_1085_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3900) begin
      mem_1084_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3899) begin
      mem_1083_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3898) begin
      mem_1082_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3897) begin
      mem_1081_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3896) begin
      mem_1080_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3895) begin
      mem_1079_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3894) begin
      mem_1078_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3893) begin
      mem_1077_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3892) begin
      mem_1076_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3891) begin
      mem_1075_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3890) begin
      mem_1074_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3889) begin
      mem_1073_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3888) begin
      mem_1072_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3887) begin
      mem_1071_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3886) begin
      mem_1070_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3885) begin
      mem_1069_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3884) begin
      mem_1068_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3883) begin
      mem_1067_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3882) begin
      mem_1066_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3881) begin
      mem_1065_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3880) begin
      mem_1064_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3879) begin
      mem_1063_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3878) begin
      mem_1062_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3877) begin
      mem_1061_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3876) begin
      mem_1060_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3875) begin
      mem_1059_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3874) begin
      mem_1058_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3873) begin
      mem_1057_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3872) begin
      mem_1056_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3871) begin
      mem_1055_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3870) begin
      mem_1054_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3869) begin
      mem_1053_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3868) begin
      mem_1052_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3867) begin
      mem_1051_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3866) begin
      mem_1050_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3865) begin
      mem_1049_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3864) begin
      mem_1048_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3863) begin
      mem_1047_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3862) begin
      mem_1046_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3861) begin
      mem_1045_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3860) begin
      mem_1044_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3859) begin
      mem_1043_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3858) begin
      mem_1042_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3857) begin
      mem_1041_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3856) begin
      mem_1040_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3855) begin
      mem_1039_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3854) begin
      mem_1038_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3853) begin
      mem_1037_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3852) begin
      mem_1036_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3851) begin
      mem_1035_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3850) begin
      mem_1034_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3849) begin
      mem_1033_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3848) begin
      mem_1032_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3847) begin
      mem_1031_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3846) begin
      mem_1030_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3845) begin
      mem_1029_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3844) begin
      mem_1028_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3843) begin
      mem_1027_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3842) begin
      mem_1026_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3841) begin
      mem_1025_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3840) begin
      mem_1024_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3839) begin
      mem_1023_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3838) begin
      mem_1022_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3837) begin
      mem_1021_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3836) begin
      mem_1020_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3835) begin
      mem_1019_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3834) begin
      mem_1018_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3833) begin
      mem_1017_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3832) begin
      mem_1016_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3831) begin
      mem_1015_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3830) begin
      mem_1014_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3829) begin
      mem_1013_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3828) begin
      mem_1012_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3827) begin
      mem_1011_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3826) begin
      mem_1010_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3825) begin
      mem_1009_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3824) begin
      mem_1008_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3823) begin
      mem_1007_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3822) begin
      mem_1006_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3821) begin
      mem_1005_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3820) begin
      mem_1004_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3819) begin
      mem_1003_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3818) begin
      mem_1002_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3817) begin
      mem_1001_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3816) begin
      mem_1000_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3815) begin
      mem_999_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3814) begin
      mem_998_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3813) begin
      mem_997_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3812) begin
      mem_996_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3811) begin
      mem_995_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3810) begin
      mem_994_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3809) begin
      mem_993_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3808) begin
      mem_992_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3807) begin
      mem_991_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3806) begin
      mem_990_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3805) begin
      mem_989_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3804) begin
      mem_988_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3803) begin
      mem_987_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3802) begin
      mem_986_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3801) begin
      mem_985_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3800) begin
      mem_984_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3799) begin
      mem_983_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3798) begin
      mem_982_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3797) begin
      mem_981_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3796) begin
      mem_980_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3795) begin
      mem_979_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3794) begin
      mem_978_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3793) begin
      mem_977_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3792) begin
      mem_976_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3791) begin
      mem_975_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3790) begin
      mem_974_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3789) begin
      mem_973_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3788) begin
      mem_972_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3787) begin
      mem_971_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3786) begin
      mem_970_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3785) begin
      mem_969_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3784) begin
      mem_968_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3783) begin
      mem_967_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3782) begin
      mem_966_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3781) begin
      mem_965_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3780) begin
      mem_964_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3779) begin
      mem_963_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3778) begin
      mem_962_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3777) begin
      mem_961_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3776) begin
      mem_960_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3775) begin
      mem_959_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3774) begin
      mem_958_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3773) begin
      mem_957_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3772) begin
      mem_956_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3771) begin
      mem_955_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3770) begin
      mem_954_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3769) begin
      mem_953_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3768) begin
      mem_952_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3767) begin
      mem_951_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3766) begin
      mem_950_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3765) begin
      mem_949_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3764) begin
      mem_948_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3763) begin
      mem_947_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3762) begin
      mem_946_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3761) begin
      mem_945_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3760) begin
      mem_944_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3759) begin
      mem_943_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3758) begin
      mem_942_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3757) begin
      mem_941_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3756) begin
      mem_940_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3755) begin
      mem_939_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3754) begin
      mem_938_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3753) begin
      mem_937_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3752) begin
      mem_936_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3751) begin
      mem_935_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3750) begin
      mem_934_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3749) begin
      mem_933_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3748) begin
      mem_932_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3747) begin
      mem_931_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3746) begin
      mem_930_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3745) begin
      mem_929_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3744) begin
      mem_928_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3743) begin
      mem_927_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3742) begin
      mem_926_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3741) begin
      mem_925_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3740) begin
      mem_924_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3739) begin
      mem_923_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3738) begin
      mem_922_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3737) begin
      mem_921_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3736) begin
      mem_920_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3735) begin
      mem_919_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3734) begin
      mem_918_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3733) begin
      mem_917_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3732) begin
      mem_916_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3731) begin
      mem_915_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3730) begin
      mem_914_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3729) begin
      mem_913_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3728) begin
      mem_912_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3727) begin
      mem_911_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3726) begin
      mem_910_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3725) begin
      mem_909_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3724) begin
      mem_908_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3723) begin
      mem_907_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3722) begin
      mem_906_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3721) begin
      mem_905_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3720) begin
      mem_904_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3719) begin
      mem_903_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3718) begin
      mem_902_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3717) begin
      mem_901_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3716) begin
      mem_900_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3715) begin
      mem_899_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3714) begin
      mem_898_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3713) begin
      mem_897_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3712) begin
      mem_896_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3711) begin
      mem_895_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3710) begin
      mem_894_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3709) begin
      mem_893_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3708) begin
      mem_892_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3707) begin
      mem_891_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3706) begin
      mem_890_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3705) begin
      mem_889_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3704) begin
      mem_888_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3703) begin
      mem_887_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3702) begin
      mem_886_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3701) begin
      mem_885_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3700) begin
      mem_884_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3699) begin
      mem_883_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3698) begin
      mem_882_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3697) begin
      mem_881_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3696) begin
      mem_880_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3695) begin
      mem_879_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3694) begin
      mem_878_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3693) begin
      mem_877_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3692) begin
      mem_876_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3691) begin
      mem_875_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3690) begin
      mem_874_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3689) begin
      mem_873_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3688) begin
      mem_872_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3687) begin
      mem_871_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3686) begin
      mem_870_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3685) begin
      mem_869_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3684) begin
      mem_868_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3683) begin
      mem_867_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3682) begin
      mem_866_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3681) begin
      mem_865_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3680) begin
      mem_864_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3679) begin
      mem_863_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3678) begin
      mem_862_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3677) begin
      mem_861_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3676) begin
      mem_860_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3675) begin
      mem_859_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3674) begin
      mem_858_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3673) begin
      mem_857_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3672) begin
      mem_856_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3671) begin
      mem_855_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3670) begin
      mem_854_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3669) begin
      mem_853_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3668) begin
      mem_852_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3667) begin
      mem_851_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3666) begin
      mem_850_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3665) begin
      mem_849_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3664) begin
      mem_848_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3663) begin
      mem_847_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3662) begin
      mem_846_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3661) begin
      mem_845_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3660) begin
      mem_844_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3659) begin
      mem_843_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3658) begin
      mem_842_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3657) begin
      mem_841_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3656) begin
      mem_840_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3655) begin
      mem_839_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3654) begin
      mem_838_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3653) begin
      mem_837_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3652) begin
      mem_836_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3651) begin
      mem_835_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3650) begin
      mem_834_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3649) begin
      mem_833_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3648) begin
      mem_832_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3647) begin
      mem_831_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3646) begin
      mem_830_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3645) begin
      mem_829_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3644) begin
      mem_828_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3643) begin
      mem_827_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3642) begin
      mem_826_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3641) begin
      mem_825_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3640) begin
      mem_824_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3639) begin
      mem_823_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3638) begin
      mem_822_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3637) begin
      mem_821_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3636) begin
      mem_820_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3635) begin
      mem_819_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3634) begin
      mem_818_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3633) begin
      mem_817_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3632) begin
      mem_816_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3631) begin
      mem_815_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3630) begin
      mem_814_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3629) begin
      mem_813_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3628) begin
      mem_812_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3627) begin
      mem_811_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3626) begin
      mem_810_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3625) begin
      mem_809_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3624) begin
      mem_808_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3623) begin
      mem_807_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3622) begin
      mem_806_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3621) begin
      mem_805_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3620) begin
      mem_804_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3619) begin
      mem_803_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3618) begin
      mem_802_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3617) begin
      mem_801_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3616) begin
      mem_800_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3615) begin
      mem_799_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3614) begin
      mem_798_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3613) begin
      mem_797_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3612) begin
      mem_796_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3611) begin
      mem_795_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3610) begin
      mem_794_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3609) begin
      mem_793_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3608) begin
      mem_792_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3607) begin
      mem_791_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3606) begin
      mem_790_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3605) begin
      mem_789_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3604) begin
      mem_788_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3603) begin
      mem_787_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3602) begin
      mem_786_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3601) begin
      mem_785_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3600) begin
      mem_784_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3599) begin
      mem_783_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3598) begin
      mem_782_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3597) begin
      mem_781_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3596) begin
      mem_780_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3595) begin
      mem_779_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3594) begin
      mem_778_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3593) begin
      mem_777_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3592) begin
      mem_776_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3591) begin
      mem_775_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3590) begin
      mem_774_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3589) begin
      mem_773_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3588) begin
      mem_772_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3587) begin
      mem_771_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3586) begin
      mem_770_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3585) begin
      mem_769_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3584) begin
      mem_768_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3583) begin
      mem_767_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3582) begin
      mem_766_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3581) begin
      mem_765_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3580) begin
      mem_764_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3579) begin
      mem_763_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3578) begin
      mem_762_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3577) begin
      mem_761_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3576) begin
      mem_760_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3575) begin
      mem_759_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3574) begin
      mem_758_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3573) begin
      mem_757_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3572) begin
      mem_756_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3571) begin
      mem_755_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3570) begin
      mem_754_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3569) begin
      mem_753_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3568) begin
      mem_752_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3567) begin
      mem_751_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3566) begin
      mem_750_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3565) begin
      mem_749_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3564) begin
      mem_748_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3563) begin
      mem_747_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3562) begin
      mem_746_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3561) begin
      mem_745_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3560) begin
      mem_744_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3559) begin
      mem_743_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3558) begin
      mem_742_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3557) begin
      mem_741_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3556) begin
      mem_740_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3555) begin
      mem_739_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3554) begin
      mem_738_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3553) begin
      mem_737_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3552) begin
      mem_736_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3551) begin
      mem_735_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3550) begin
      mem_734_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3549) begin
      mem_733_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3548) begin
      mem_732_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3547) begin
      mem_731_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3546) begin
      mem_730_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3545) begin
      mem_729_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3544) begin
      mem_728_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3543) begin
      mem_727_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3542) begin
      mem_726_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3541) begin
      mem_725_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3540) begin
      mem_724_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3539) begin
      mem_723_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3538) begin
      mem_722_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3537) begin
      mem_721_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3536) begin
      mem_720_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3535) begin
      mem_719_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3534) begin
      mem_718_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3533) begin
      mem_717_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3532) begin
      mem_716_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3531) begin
      mem_715_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3530) begin
      mem_714_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3529) begin
      mem_713_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3528) begin
      mem_712_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3527) begin
      mem_711_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3526) begin
      mem_710_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3525) begin
      mem_709_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3524) begin
      mem_708_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3523) begin
      mem_707_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3522) begin
      mem_706_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3521) begin
      mem_705_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3520) begin
      mem_704_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3519) begin
      mem_703_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3518) begin
      mem_702_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3517) begin
      mem_701_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3516) begin
      mem_700_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3515) begin
      mem_699_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3514) begin
      mem_698_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3513) begin
      mem_697_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3512) begin
      mem_696_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3511) begin
      mem_695_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3510) begin
      mem_694_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3509) begin
      mem_693_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3508) begin
      mem_692_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3507) begin
      mem_691_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3506) begin
      mem_690_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3505) begin
      mem_689_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3504) begin
      mem_688_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3503) begin
      mem_687_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3502) begin
      mem_686_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3501) begin
      mem_685_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3500) begin
      mem_684_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3499) begin
      mem_683_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3498) begin
      mem_682_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3497) begin
      mem_681_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3496) begin
      mem_680_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3495) begin
      mem_679_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3494) begin
      mem_678_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3493) begin
      mem_677_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3492) begin
      mem_676_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3491) begin
      mem_675_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3490) begin
      mem_674_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3489) begin
      mem_673_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3488) begin
      mem_672_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3487) begin
      mem_671_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3486) begin
      mem_670_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3485) begin
      mem_669_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3484) begin
      mem_668_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3483) begin
      mem_667_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3482) begin
      mem_666_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3481) begin
      mem_665_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3480) begin
      mem_664_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3479) begin
      mem_663_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3478) begin
      mem_662_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3477) begin
      mem_661_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3476) begin
      mem_660_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3475) begin
      mem_659_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3474) begin
      mem_658_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3473) begin
      mem_657_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3472) begin
      mem_656_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3471) begin
      mem_655_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3470) begin
      mem_654_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3469) begin
      mem_653_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3468) begin
      mem_652_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3467) begin
      mem_651_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3466) begin
      mem_650_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3465) begin
      mem_649_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3464) begin
      mem_648_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3463) begin
      mem_647_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3462) begin
      mem_646_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3461) begin
      mem_645_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3460) begin
      mem_644_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3459) begin
      mem_643_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3458) begin
      mem_642_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3457) begin
      mem_641_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3456) begin
      mem_640_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3455) begin
      mem_639_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3454) begin
      mem_638_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3453) begin
      mem_637_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3452) begin
      mem_636_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3451) begin
      mem_635_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3450) begin
      mem_634_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3449) begin
      mem_633_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3448) begin
      mem_632_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3447) begin
      mem_631_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3446) begin
      mem_630_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3445) begin
      mem_629_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3444) begin
      mem_628_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3443) begin
      mem_627_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3442) begin
      mem_626_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3441) begin
      mem_625_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3440) begin
      mem_624_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3439) begin
      mem_623_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3438) begin
      mem_622_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3437) begin
      mem_621_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3436) begin
      mem_620_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3435) begin
      mem_619_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3434) begin
      mem_618_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3433) begin
      mem_617_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3432) begin
      mem_616_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3431) begin
      mem_615_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3430) begin
      mem_614_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3429) begin
      mem_613_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3428) begin
      mem_612_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3427) begin
      mem_611_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3426) begin
      mem_610_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3425) begin
      mem_609_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3424) begin
      mem_608_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3423) begin
      mem_607_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3422) begin
      mem_606_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3421) begin
      mem_605_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3420) begin
      mem_604_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3419) begin
      mem_603_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3418) begin
      mem_602_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3417) begin
      mem_601_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3416) begin
      mem_600_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3415) begin
      mem_599_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3414) begin
      mem_598_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3413) begin
      mem_597_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3412) begin
      mem_596_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3411) begin
      mem_595_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3410) begin
      mem_594_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3409) begin
      mem_593_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3408) begin
      mem_592_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3407) begin
      mem_591_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3406) begin
      mem_590_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3405) begin
      mem_589_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3404) begin
      mem_588_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3403) begin
      mem_587_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3402) begin
      mem_586_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3401) begin
      mem_585_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3400) begin
      mem_584_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3399) begin
      mem_583_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3398) begin
      mem_582_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3397) begin
      mem_581_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3396) begin
      mem_580_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3395) begin
      mem_579_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3394) begin
      mem_578_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3393) begin
      mem_577_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3392) begin
      mem_576_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3391) begin
      mem_575_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3390) begin
      mem_574_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3389) begin
      mem_573_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3388) begin
      mem_572_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3387) begin
      mem_571_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3386) begin
      mem_570_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3385) begin
      mem_569_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3384) begin
      mem_568_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3383) begin
      mem_567_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3382) begin
      mem_566_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3381) begin
      mem_565_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3380) begin
      mem_564_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3379) begin
      mem_563_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3378) begin
      mem_562_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3377) begin
      mem_561_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3376) begin
      mem_560_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3375) begin
      mem_559_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3374) begin
      mem_558_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3373) begin
      mem_557_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3372) begin
      mem_556_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3371) begin
      mem_555_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3370) begin
      mem_554_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3369) begin
      mem_553_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3368) begin
      mem_552_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3367) begin
      mem_551_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3366) begin
      mem_550_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3365) begin
      mem_549_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3364) begin
      mem_548_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3363) begin
      mem_547_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3362) begin
      mem_546_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3361) begin
      mem_545_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3360) begin
      mem_544_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3359) begin
      mem_543_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3358) begin
      mem_542_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3357) begin
      mem_541_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3356) begin
      mem_540_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3355) begin
      mem_539_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3354) begin
      mem_538_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3353) begin
      mem_537_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3352) begin
      mem_536_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3351) begin
      mem_535_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3350) begin
      mem_534_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3349) begin
      mem_533_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3348) begin
      mem_532_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3347) begin
      mem_531_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3346) begin
      mem_530_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3345) begin
      mem_529_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3344) begin
      mem_528_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3343) begin
      mem_527_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3342) begin
      mem_526_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3341) begin
      mem_525_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3340) begin
      mem_524_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3339) begin
      mem_523_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3338) begin
      mem_522_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3337) begin
      mem_521_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3336) begin
      mem_520_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3335) begin
      mem_519_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3334) begin
      mem_518_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3333) begin
      mem_517_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3332) begin
      mem_516_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3331) begin
      mem_515_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3330) begin
      mem_514_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3329) begin
      mem_513_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3328) begin
      mem_512_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3327) begin
      mem_511_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3326) begin
      mem_510_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3325) begin
      mem_509_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3324) begin
      mem_508_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3323) begin
      mem_507_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3322) begin
      mem_506_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3321) begin
      mem_505_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3320) begin
      mem_504_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3319) begin
      mem_503_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3318) begin
      mem_502_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3317) begin
      mem_501_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3316) begin
      mem_500_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3315) begin
      mem_499_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3314) begin
      mem_498_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3313) begin
      mem_497_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3312) begin
      mem_496_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3311) begin
      mem_495_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3310) begin
      mem_494_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3309) begin
      mem_493_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3308) begin
      mem_492_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3307) begin
      mem_491_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3306) begin
      mem_490_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3305) begin
      mem_489_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3304) begin
      mem_488_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3303) begin
      mem_487_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3302) begin
      mem_486_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3301) begin
      mem_485_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3300) begin
      mem_484_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3299) begin
      mem_483_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3298) begin
      mem_482_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3297) begin
      mem_481_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3296) begin
      mem_480_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3295) begin
      mem_479_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3294) begin
      mem_478_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3293) begin
      mem_477_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3292) begin
      mem_476_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3291) begin
      mem_475_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3290) begin
      mem_474_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3289) begin
      mem_473_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3288) begin
      mem_472_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3287) begin
      mem_471_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3286) begin
      mem_470_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3285) begin
      mem_469_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3284) begin
      mem_468_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3283) begin
      mem_467_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3282) begin
      mem_466_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3281) begin
      mem_465_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3280) begin
      mem_464_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3279) begin
      mem_463_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3278) begin
      mem_462_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3277) begin
      mem_461_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3276) begin
      mem_460_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3275) begin
      mem_459_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3274) begin
      mem_458_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3273) begin
      mem_457_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3272) begin
      mem_456_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3271) begin
      mem_455_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3270) begin
      mem_454_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3269) begin
      mem_453_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3268) begin
      mem_452_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3267) begin
      mem_451_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3266) begin
      mem_450_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3265) begin
      mem_449_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3264) begin
      mem_448_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3263) begin
      mem_447_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3262) begin
      mem_446_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3261) begin
      mem_445_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3260) begin
      mem_444_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3259) begin
      mem_443_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3258) begin
      mem_442_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3257) begin
      mem_441_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3256) begin
      mem_440_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3255) begin
      mem_439_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3254) begin
      mem_438_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3253) begin
      mem_437_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3252) begin
      mem_436_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3251) begin
      mem_435_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3250) begin
      mem_434_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3249) begin
      mem_433_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3248) begin
      mem_432_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3247) begin
      mem_431_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3246) begin
      mem_430_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3245) begin
      mem_429_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3244) begin
      mem_428_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3243) begin
      mem_427_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3242) begin
      mem_426_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3241) begin
      mem_425_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3240) begin
      mem_424_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3239) begin
      mem_423_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3238) begin
      mem_422_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3237) begin
      mem_421_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3236) begin
      mem_420_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3235) begin
      mem_419_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3234) begin
      mem_418_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3233) begin
      mem_417_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3232) begin
      mem_416_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3231) begin
      mem_415_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3230) begin
      mem_414_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3229) begin
      mem_413_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3228) begin
      mem_412_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3227) begin
      mem_411_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3226) begin
      mem_410_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3225) begin
      mem_409_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3224) begin
      mem_408_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3223) begin
      mem_407_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3222) begin
      mem_406_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3221) begin
      mem_405_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3220) begin
      mem_404_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3219) begin
      mem_403_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3218) begin
      mem_402_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3217) begin
      mem_401_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3216) begin
      mem_400_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3215) begin
      mem_399_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3214) begin
      mem_398_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3213) begin
      mem_397_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3212) begin
      mem_396_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3211) begin
      mem_395_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3210) begin
      mem_394_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3209) begin
      mem_393_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3208) begin
      mem_392_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3207) begin
      mem_391_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3206) begin
      mem_390_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3205) begin
      mem_389_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3204) begin
      mem_388_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3203) begin
      mem_387_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3202) begin
      mem_386_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3201) begin
      mem_385_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3200) begin
      mem_384_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3199) begin
      mem_383_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3198) begin
      mem_382_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3197) begin
      mem_381_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3196) begin
      mem_380_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3195) begin
      mem_379_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3194) begin
      mem_378_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3193) begin
      mem_377_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3192) begin
      mem_376_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3191) begin
      mem_375_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3190) begin
      mem_374_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3189) begin
      mem_373_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3188) begin
      mem_372_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3187) begin
      mem_371_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3186) begin
      mem_370_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3185) begin
      mem_369_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3184) begin
      mem_368_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3183) begin
      mem_367_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3182) begin
      mem_366_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3181) begin
      mem_365_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3180) begin
      mem_364_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3179) begin
      mem_363_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3178) begin
      mem_362_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3177) begin
      mem_361_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3176) begin
      mem_360_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3175) begin
      mem_359_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3174) begin
      mem_358_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3173) begin
      mem_357_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3172) begin
      mem_356_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3171) begin
      mem_355_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3170) begin
      mem_354_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3169) begin
      mem_353_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3168) begin
      mem_352_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3167) begin
      mem_351_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3166) begin
      mem_350_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3165) begin
      mem_349_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3164) begin
      mem_348_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3163) begin
      mem_347_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3162) begin
      mem_346_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3161) begin
      mem_345_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3160) begin
      mem_344_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3159) begin
      mem_343_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3158) begin
      mem_342_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3157) begin
      mem_341_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3156) begin
      mem_340_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3155) begin
      mem_339_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3154) begin
      mem_338_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3153) begin
      mem_337_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3152) begin
      mem_336_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3151) begin
      mem_335_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3150) begin
      mem_334_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3149) begin
      mem_333_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3148) begin
      mem_332_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3147) begin
      mem_331_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3146) begin
      mem_330_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3145) begin
      mem_329_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3144) begin
      mem_328_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3143) begin
      mem_327_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3142) begin
      mem_326_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3141) begin
      mem_325_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3140) begin
      mem_324_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3139) begin
      mem_323_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3138) begin
      mem_322_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3137) begin
      mem_321_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3136) begin
      mem_320_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3135) begin
      mem_319_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3134) begin
      mem_318_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3133) begin
      mem_317_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3132) begin
      mem_316_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3131) begin
      mem_315_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3130) begin
      mem_314_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3129) begin
      mem_313_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3128) begin
      mem_312_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3127) begin
      mem_311_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3126) begin
      mem_310_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3125) begin
      mem_309_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3124) begin
      mem_308_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3123) begin
      mem_307_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3122) begin
      mem_306_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3121) begin
      mem_305_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3120) begin
      mem_304_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3119) begin
      mem_303_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3118) begin
      mem_302_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3117) begin
      mem_301_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3116) begin
      mem_300_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3115) begin
      mem_299_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3114) begin
      mem_298_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3113) begin
      mem_297_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3112) begin
      mem_296_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3111) begin
      mem_295_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3110) begin
      mem_294_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3109) begin
      mem_293_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3108) begin
      mem_292_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3107) begin
      mem_291_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3106) begin
      mem_290_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3105) begin
      mem_289_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3104) begin
      mem_288_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3103) begin
      mem_287_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3102) begin
      mem_286_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3101) begin
      mem_285_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3100) begin
      mem_284_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3099) begin
      mem_283_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3098) begin
      mem_282_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3097) begin
      mem_281_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3096) begin
      mem_280_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3095) begin
      mem_279_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3094) begin
      mem_278_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3093) begin
      mem_277_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3092) begin
      mem_276_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3091) begin
      mem_275_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3090) begin
      mem_274_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3089) begin
      mem_273_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3088) begin
      mem_272_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3087) begin
      mem_271_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3086) begin
      mem_270_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3085) begin
      mem_269_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3084) begin
      mem_268_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3083) begin
      mem_267_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3082) begin
      mem_266_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3081) begin
      mem_265_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3080) begin
      mem_264_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3079) begin
      mem_263_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3078) begin
      mem_262_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3077) begin
      mem_261_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3076) begin
      mem_260_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3075) begin
      mem_259_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3074) begin
      mem_258_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3073) begin
      mem_257_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3072) begin
      mem_256_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3071) begin
      mem_255_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3070) begin
      mem_254_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3069) begin
      mem_253_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3068) begin
      mem_252_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3067) begin
      mem_251_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3066) begin
      mem_250_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3065) begin
      mem_249_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3064) begin
      mem_248_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3063) begin
      mem_247_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3062) begin
      mem_246_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3061) begin
      mem_245_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3060) begin
      mem_244_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3059) begin
      mem_243_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3058) begin
      mem_242_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3057) begin
      mem_241_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3056) begin
      mem_240_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3055) begin
      mem_239_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3054) begin
      mem_238_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3053) begin
      mem_237_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3052) begin
      mem_236_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3051) begin
      mem_235_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3050) begin
      mem_234_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3049) begin
      mem_233_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3048) begin
      mem_232_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3047) begin
      mem_231_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3046) begin
      mem_230_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3045) begin
      mem_229_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3044) begin
      mem_228_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3043) begin
      mem_227_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3042) begin
      mem_226_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3041) begin
      mem_225_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3040) begin
      mem_224_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3039) begin
      mem_223_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3038) begin
      mem_222_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3037) begin
      mem_221_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3036) begin
      mem_220_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3035) begin
      mem_219_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3034) begin
      mem_218_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3033) begin
      mem_217_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3032) begin
      mem_216_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3031) begin
      mem_215_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3030) begin
      mem_214_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3029) begin
      mem_213_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3028) begin
      mem_212_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3027) begin
      mem_211_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3026) begin
      mem_210_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3025) begin
      mem_209_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3024) begin
      mem_208_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3023) begin
      mem_207_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3022) begin
      mem_206_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3021) begin
      mem_205_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3020) begin
      mem_204_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3019) begin
      mem_203_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3018) begin
      mem_202_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3017) begin
      mem_201_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3016) begin
      mem_200_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3015) begin
      mem_199_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N3014) begin
      mem_198_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N3013) begin
      mem_197_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N3012) begin
      mem_196_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N3011) begin
      mem_195_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N3010) begin
      mem_194_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N3009) begin
      mem_193_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N3008) begin
      mem_192_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N3007) begin
      mem_191_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N3006) begin
      mem_190_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N3005) begin
      mem_189_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N3004) begin
      mem_188_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N3003) begin
      mem_187_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N3002) begin
      mem_186_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N3001) begin
      mem_185_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N3000) begin
      mem_184_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2999) begin
      mem_183_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2998) begin
      mem_182_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2997) begin
      mem_181_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2996) begin
      mem_180_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2995) begin
      mem_179_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2994) begin
      mem_178_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2993) begin
      mem_177_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2992) begin
      mem_176_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2991) begin
      mem_175_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2990) begin
      mem_174_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2989) begin
      mem_173_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2988) begin
      mem_172_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2987) begin
      mem_171_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2986) begin
      mem_170_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2985) begin
      mem_169_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2984) begin
      mem_168_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2983) begin
      mem_167_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2982) begin
      mem_166_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2981) begin
      mem_165_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2980) begin
      mem_164_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2979) begin
      mem_163_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2978) begin
      mem_162_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2977) begin
      mem_161_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2976) begin
      mem_160_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2975) begin
      mem_159_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2974) begin
      mem_158_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2973) begin
      mem_157_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2972) begin
      mem_156_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2971) begin
      mem_155_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2970) begin
      mem_154_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2969) begin
      mem_153_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2968) begin
      mem_152_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2967) begin
      mem_151_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2966) begin
      mem_150_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2965) begin
      mem_149_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2964) begin
      mem_148_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2963) begin
      mem_147_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2962) begin
      mem_146_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2961) begin
      mem_145_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2960) begin
      mem_144_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2959) begin
      mem_143_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2958) begin
      mem_142_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2957) begin
      mem_141_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2956) begin
      mem_140_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2955) begin
      mem_139_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2954) begin
      mem_138_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2953) begin
      mem_137_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2952) begin
      mem_136_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2951) begin
      mem_135_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2950) begin
      mem_134_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2949) begin
      mem_133_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2948) begin
      mem_132_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2947) begin
      mem_131_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2946) begin
      mem_130_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2945) begin
      mem_129_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2944) begin
      mem_128_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2943) begin
      mem_127_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2942) begin
      mem_126_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2941) begin
      mem_125_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2940) begin
      mem_124_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2939) begin
      mem_123_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2938) begin
      mem_122_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2937) begin
      mem_121_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2936) begin
      mem_120_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2935) begin
      mem_119_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2934) begin
      mem_118_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2933) begin
      mem_117_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2932) begin
      mem_116_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2931) begin
      mem_115_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2930) begin
      mem_114_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2929) begin
      mem_113_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2928) begin
      mem_112_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2927) begin
      mem_111_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2926) begin
      mem_110_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2925) begin
      mem_109_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2924) begin
      mem_108_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2923) begin
      mem_107_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2922) begin
      mem_106_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2921) begin
      mem_105_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2920) begin
      mem_104_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2919) begin
      mem_103_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2918) begin
      mem_102_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2917) begin
      mem_101_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2916) begin
      mem_100_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2915) begin
      mem_99_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2914) begin
      mem_98_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2913) begin
      mem_97_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2912) begin
      mem_96_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2911) begin
      mem_95_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2910) begin
      mem_94_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2909) begin
      mem_93_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2908) begin
      mem_92_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2907) begin
      mem_91_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2906) begin
      mem_90_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2905) begin
      mem_89_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2904) begin
      mem_88_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2903) begin
      mem_87_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2902) begin
      mem_86_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2901) begin
      mem_85_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2900) begin
      mem_84_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2899) begin
      mem_83_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2898) begin
      mem_82_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2897) begin
      mem_81_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2896) begin
      mem_80_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2895) begin
      mem_79_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2894) begin
      mem_78_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2893) begin
      mem_77_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2892) begin
      mem_76_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2891) begin
      mem_75_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2890) begin
      mem_74_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2889) begin
      mem_73_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2888) begin
      mem_72_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2887) begin
      mem_71_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2886) begin
      mem_70_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2885) begin
      mem_69_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2884) begin
      mem_68_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2883) begin
      mem_67_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2882) begin
      mem_66_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2881) begin
      mem_65_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2880) begin
      mem_64_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2879) begin
      mem_63_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2878) begin
      mem_62_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2877) begin
      mem_61_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2876) begin
      mem_60_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2875) begin
      mem_59_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2874) begin
      mem_58_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2873) begin
      mem_57_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2872) begin
      mem_56_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2871) begin
      mem_55_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2870) begin
      mem_54_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2869) begin
      mem_53_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2868) begin
      mem_52_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2867) begin
      mem_51_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2866) begin
      mem_50_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2865) begin
      mem_49_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2864) begin
      mem_48_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2863) begin
      mem_47_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2862) begin
      mem_46_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2861) begin
      mem_45_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2860) begin
      mem_44_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2859) begin
      mem_43_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2858) begin
      mem_42_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2857) begin
      mem_41_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2856) begin
      mem_40_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2855) begin
      mem_39_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2854) begin
      mem_38_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2853) begin
      mem_37_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2852) begin
      mem_36_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2851) begin
      mem_35_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2850) begin
      mem_34_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2849) begin
      mem_33_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2848) begin
      mem_32_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2847) begin
      mem_31_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2846) begin
      mem_30_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2845) begin
      mem_29_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2844) begin
      mem_28_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2843) begin
      mem_27_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2842) begin
      mem_26_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2841) begin
      mem_25_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2840) begin
      mem_24_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2839) begin
      mem_23_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2838) begin
      mem_22_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2837) begin
      mem_21_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2836) begin
      mem_20_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2835) begin
      mem_19_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2834) begin
      mem_18_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2833) begin
      mem_17_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2832) begin
      mem_16_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2831) begin
      mem_15_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N2830) begin
      mem_14_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(N2829) begin
      mem_13_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(N2828) begin
      mem_12_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(N2827) begin
      mem_11_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(N2826) begin
      mem_10_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(N2825) begin
      mem_9_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(N2824) begin
      mem_8_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(N2823) begin
      mem_7_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(N2822) begin
      mem_6_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N2821) begin
      mem_5_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N2820) begin
      mem_4_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N2819) begin
      mem_3_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N2818) begin
      mem_2_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N2817) begin
      mem_1_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N2816) begin
      mem_0_sv2v_reg <= data_i[0];
    end 
  end

  assign N4736 = addr_i[6] & N4769;
  assign N4737 = addr_i[6] & N4770;
  assign N4738 = addr_i[6] & N4771;
  assign N595 = N4736 & N4789;
  assign N594 = N4736 & N4790;
  assign N593 = N4736 & N4791;
  assign N592 = N4736 & N4792;
  assign N591 = N4736 & N4793;
  assign N590 = N4736 & N4794;
  assign N589 = N4736 & N4795;
  assign N588 = N4736 & N4796;
  assign N587 = N4736 & N4797;
  assign N586 = N4736 & N4798;
  assign N585 = N4736 & N4799;
  assign N584 = N4736 & N4800;
  assign N583 = N4736 & N4801;
  assign N582 = N4736 & N4802;
  assign N581 = N4736 & N4803;
  assign N580 = N4736 & N4804;
  assign N579 = N4737 & N4789;
  assign N578 = N4737 & N4790;
  assign N577 = N4737 & N4791;
  assign N576 = N4737 & N4792;
  assign N575 = N4737 & N4793;
  assign N574 = N4737 & N4794;
  assign N573 = N4737 & N4795;
  assign N572 = N4737 & N4796;
  assign N571 = N4737 & N4797;
  assign N570 = N4737 & N4798;
  assign N569 = N4737 & N4799;
  assign N568 = N4737 & N4800;
  assign N567 = N4737 & N4801;
  assign N566 = N4737 & N4802;
  assign N565 = N4737 & N4803;
  assign N564 = N4737 & N4804;
  assign N563 = N4738 & N4789;
  assign N562 = N4738 & N4790;
  assign N561 = N4738 & N4791;
  assign N560 = N4738 & N4792;
  assign N559 = N4738 & N4793;
  assign N558 = N4738 & N4794;
  assign N557 = N4738 & N4795;
  assign N556 = N4738 & N4796;
  assign N555 = N4738 & N4797;
  assign N554 = N4738 & N4798;
  assign N553 = N4738 & N4799;
  assign N552 = N4738 & N4800;
  assign N551 = N4738 & N4801;
  assign N550 = N4738 & N4802;
  assign N549 = N4738 & N4803;
  assign N548 = N4738 & N4804;
  assign N4739 = addr_i[6] & N4769;
  assign N4740 = addr_i[6] & N4770;
  assign N4741 = addr_i[6] & N4771;
  assign N1417 = N4739 & N4789;
  assign N1416 = N4739 & N4790;
  assign N1415 = N4739 & N4791;
  assign N1414 = N4739 & N4792;
  assign N1413 = N4739 & N4793;
  assign N1412 = N4739 & N4794;
  assign N1411 = N4739 & N4795;
  assign N1410 = N4739 & N4796;
  assign N1409 = N4739 & N4797;
  assign N1408 = N4739 & N4798;
  assign N1407 = N4739 & N4799;
  assign N1406 = N4739 & N4800;
  assign N1405 = N4739 & N4801;
  assign N1404 = N4739 & N4802;
  assign N1403 = N4739 & N4803;
  assign N1402 = N4739 & N4804;
  assign N1401 = N4740 & N4789;
  assign N1400 = N4740 & N4790;
  assign N1399 = N4740 & N4791;
  assign N1398 = N4740 & N4792;
  assign N1397 = N4740 & N4793;
  assign N1396 = N4740 & N4794;
  assign N1395 = N4740 & N4795;
  assign N1394 = N4740 & N4796;
  assign N1393 = N4740 & N4797;
  assign N1392 = N4740 & N4798;
  assign N1391 = N4740 & N4799;
  assign N1390 = N4740 & N4800;
  assign N1389 = N4740 & N4801;
  assign N1388 = N4740 & N4802;
  assign N1387 = N4740 & N4803;
  assign N1386 = N4740 & N4804;
  assign N1385 = N4741 & N4789;
  assign N1384 = N4741 & N4790;
  assign N1383 = N4741 & N4791;
  assign N1382 = N4741 & N4792;
  assign N1381 = N4741 & N4793;
  assign N1380 = N4741 & N4794;
  assign N1379 = N4741 & N4795;
  assign N1378 = N4741 & N4796;
  assign N1377 = N4741 & N4797;
  assign N1376 = N4741 & N4798;
  assign N1375 = N4741 & N4799;
  assign N1374 = N4741 & N4800;
  assign N1373 = N4741 & N4801;
  assign N1372 = N4741 & N4802;
  assign N1371 = N4741 & N4803;
  assign N1370 = N4741 & N4804;
  assign N1626 = N4747 & N4789;
  assign N1625 = N4747 & N4790;
  assign N1624 = N4747 & N4791;
  assign N1623 = N4747 & N4792;
  assign N1622 = N4747 & N4793;
  assign N1621 = N4747 & N4794;
  assign N1620 = N4747 & N4795;
  assign N1619 = N4747 & N4796;
  assign N1618 = N4747 & N4797;
  assign N1617 = N4747 & N4798;
  assign N1616 = N4747 & N4799;
  assign N1615 = N4747 & N4800;
  assign N1614 = N4747 & N4801;
  assign N1613 = N4747 & N4802;
  assign N1612 = N4747 & N4803;
  assign N1611 = N4747 & N4804;
  assign N1610 = N4748 & N4789;
  assign N1609 = N4748 & N4790;
  assign N1608 = N4748 & N4791;
  assign N1607 = N4748 & N4792;
  assign N1606 = N4748 & N4793;
  assign N1605 = N4748 & N4794;
  assign N1604 = N4748 & N4795;
  assign N1603 = N4748 & N4796;
  assign N1602 = N4748 & N4797;
  assign N1601 = N4748 & N4798;
  assign N1600 = N4748 & N4799;
  assign N1599 = N4748 & N4800;
  assign N1598 = N4748 & N4801;
  assign N1597 = N4748 & N4802;
  assign N1596 = N4748 & N4803;
  assign N1595 = N4748 & N4804;
  assign N1594 = N4749 & N4789;
  assign N1593 = N4749 & N4790;
  assign N1592 = N4749 & N4791;
  assign N1591 = N4749 & N4792;
  assign N1590 = N4749 & N4793;
  assign N1589 = N4749 & N4794;
  assign N1588 = N4749 & N4795;
  assign N1587 = N4749 & N4796;
  assign N1586 = N4749 & N4797;
  assign N1585 = N4749 & N4798;
  assign N1584 = N4749 & N4799;
  assign N1583 = N4749 & N4800;
  assign N1582 = N4749 & N4801;
  assign N1581 = N4749 & N4802;
  assign N1580 = N4749 & N4803;
  assign N1579 = N4749 & N4804;
  assign N1578 = N4750 & N4789;
  assign N1577 = N4750 & N4790;
  assign N1576 = N4750 & N4791;
  assign N1575 = N4750 & N4792;
  assign N1574 = N4750 & N4793;
  assign N1573 = N4750 & N4794;
  assign N1572 = N4750 & N4795;
  assign N1571 = N4750 & N4796;
  assign N1570 = N4750 & N4797;
  assign N1569 = N4750 & N4798;
  assign N1568 = N4750 & N4799;
  assign N1567 = N4750 & N4800;
  assign N1566 = N4750 & N4801;
  assign N1565 = N4750 & N4802;
  assign N1564 = N4750 & N4803;
  assign N1563 = N4750 & N4804;
  assign N1562 = N4751 & N4789;
  assign N1561 = N4751 & N4790;
  assign N1560 = N4751 & N4791;
  assign N1559 = N4751 & N4792;
  assign N1558 = N4751 & N4793;
  assign N1557 = N4751 & N4794;
  assign N1556 = N4751 & N4795;
  assign N1555 = N4751 & N4796;
  assign N1554 = N4751 & N4797;
  assign N1553 = N4751 & N4798;
  assign N1552 = N4751 & N4799;
  assign N1551 = N4751 & N4800;
  assign N1550 = N4751 & N4801;
  assign N1549 = N4751 & N4802;
  assign N1548 = N4751 & N4803;
  assign N1547 = N4751 & N4804;
  assign N1835 = N4742 & N4789;
  assign N1834 = N4742 & N4790;
  assign N1833 = N4742 & N4791;
  assign N1832 = N4742 & N4792;
  assign N1831 = N4742 & N4793;
  assign N1830 = N4742 & N4794;
  assign N1829 = N4742 & N4795;
  assign N1828 = N4742 & N4796;
  assign N1827 = N4742 & N4797;
  assign N1826 = N4742 & N4798;
  assign N1825 = N4742 & N4799;
  assign N1824 = N4742 & N4800;
  assign N1823 = N4742 & N4801;
  assign N1822 = N4742 & N4802;
  assign N1821 = N4742 & N4803;
  assign N1820 = N4742 & N4804;
  assign N1819 = N4743 & N4789;
  assign N1818 = N4743 & N4790;
  assign N1817 = N4743 & N4791;
  assign N1816 = N4743 & N4792;
  assign N1815 = N4743 & N4793;
  assign N1814 = N4743 & N4794;
  assign N1813 = N4743 & N4795;
  assign N1812 = N4743 & N4796;
  assign N1811 = N4743 & N4797;
  assign N1810 = N4743 & N4798;
  assign N1809 = N4743 & N4799;
  assign N1808 = N4743 & N4800;
  assign N1807 = N4743 & N4801;
  assign N1806 = N4743 & N4802;
  assign N1805 = N4743 & N4803;
  assign N1804 = N4743 & N4804;
  assign N1803 = N4744 & N4789;
  assign N1802 = N4744 & N4790;
  assign N1801 = N4744 & N4791;
  assign N1800 = N4744 & N4792;
  assign N1799 = N4744 & N4793;
  assign N1798 = N4744 & N4794;
  assign N1797 = N4744 & N4795;
  assign N1796 = N4744 & N4796;
  assign N1795 = N4744 & N4797;
  assign N1794 = N4744 & N4798;
  assign N1793 = N4744 & N4799;
  assign N1792 = N4744 & N4800;
  assign N1791 = N4744 & N4801;
  assign N1790 = N4744 & N4802;
  assign N1789 = N4744 & N4803;
  assign N1788 = N4744 & N4804;
  assign N1787 = N4745 & N4789;
  assign N1786 = N4745 & N4790;
  assign N1785 = N4745 & N4791;
  assign N1784 = N4745 & N4792;
  assign N1783 = N4745 & N4793;
  assign N1782 = N4745 & N4794;
  assign N1781 = N4745 & N4795;
  assign N1780 = N4745 & N4796;
  assign N1779 = N4745 & N4797;
  assign N1778 = N4745 & N4798;
  assign N1777 = N4745 & N4799;
  assign N1776 = N4745 & N4800;
  assign N1775 = N4745 & N4801;
  assign N1774 = N4745 & N4802;
  assign N1773 = N4745 & N4803;
  assign N1772 = N4745 & N4804;
  assign N1771 = N4746 & N4789;
  assign N1770 = N4746 & N4790;
  assign N1769 = N4746 & N4791;
  assign N1768 = N4746 & N4792;
  assign N1767 = N4746 & N4793;
  assign N1766 = N4746 & N4794;
  assign N1765 = N4746 & N4795;
  assign N1764 = N4746 & N4796;
  assign N1763 = N4746 & N4797;
  assign N1762 = N4746 & N4798;
  assign N1761 = N4746 & N4799;
  assign N1760 = N4746 & N4800;
  assign N1759 = N4746 & N4801;
  assign N1758 = N4746 & N4802;
  assign N1757 = N4746 & N4803;
  assign N1756 = N4746 & N4804;
  assign N4742 = addr_i[6] & N4772;
  assign N4743 = N4768 & N4769;
  assign N4744 = N4768 & N4770;
  assign N4745 = N4768 & N4771;
  assign N4746 = N4768 & N4772;
  assign N2173 = N4742 & N4752;
  assign N2172 = N4742 & N4753;
  assign N2171 = N4742 & N4754;
  assign N2170 = N4742 & N4755;
  assign N2169 = N4742 & N4756;
  assign N2168 = N4742 & N4757;
  assign N2167 = N4742 & N4758;
  assign N2166 = N4742 & N4759;
  assign N2165 = N4742 & N4760;
  assign N2164 = N4742 & N4761;
  assign N2163 = N4742 & N4762;
  assign N2162 = N4742 & N4763;
  assign N2161 = N4742 & N4764;
  assign N2160 = N4742 & N4765;
  assign N2159 = N4742 & N4766;
  assign N2158 = N4742 & N4767;
  assign N2157 = N4743 & N4752;
  assign N2156 = N4743 & N4753;
  assign N2155 = N4743 & N4754;
  assign N2154 = N4743 & N4755;
  assign N2153 = N4743 & N4756;
  assign N2152 = N4743 & N4757;
  assign N2151 = N4743 & N4758;
  assign N2150 = N4743 & N4759;
  assign N2149 = N4743 & N4760;
  assign N2148 = N4743 & N4761;
  assign N2147 = N4743 & N4762;
  assign N2146 = N4743 & N4763;
  assign N2145 = N4743 & N4764;
  assign N2144 = N4743 & N4765;
  assign N2143 = N4743 & N4766;
  assign N2142 = N4743 & N4767;
  assign N2141 = N4744 & N4752;
  assign N2140 = N4744 & N4753;
  assign N2139 = N4744 & N4754;
  assign N2138 = N4744 & N4755;
  assign N2137 = N4744 & N4756;
  assign N2136 = N4744 & N4757;
  assign N2135 = N4744 & N4758;
  assign N2134 = N4744 & N4759;
  assign N2133 = N4744 & N4760;
  assign N2132 = N4744 & N4761;
  assign N2131 = N4744 & N4762;
  assign N2130 = N4744 & N4763;
  assign N2129 = N4744 & N4764;
  assign N2128 = N4744 & N4765;
  assign N2127 = N4744 & N4766;
  assign N2126 = N4744 & N4767;
  assign N2125 = N4745 & N4752;
  assign N2124 = N4745 & N4753;
  assign N2123 = N4745 & N4754;
  assign N2122 = N4745 & N4755;
  assign N2121 = N4745 & N4756;
  assign N2120 = N4745 & N4757;
  assign N2119 = N4745 & N4758;
  assign N2118 = N4745 & N4759;
  assign N2117 = N4745 & N4760;
  assign N2116 = N4745 & N4761;
  assign N2115 = N4745 & N4762;
  assign N2114 = N4745 & N4763;
  assign N2113 = N4745 & N4764;
  assign N2112 = N4745 & N4765;
  assign N2111 = N4745 & N4766;
  assign N2110 = N4745 & N4767;
  assign N2109 = N4746 & N4752;
  assign N2108 = N4746 & N4753;
  assign N2107 = N4746 & N4754;
  assign N2106 = N4746 & N4755;
  assign N2105 = N4746 & N4756;
  assign N2104 = N4746 & N4757;
  assign N2103 = N4746 & N4758;
  assign N2102 = N4746 & N4759;
  assign N2101 = N4746 & N4760;
  assign N2100 = N4746 & N4761;
  assign N2099 = N4746 & N4762;
  assign N2098 = N4746 & N4763;
  assign N2097 = N4746 & N4764;
  assign N2096 = N4746 & N4765;
  assign N2095 = N4746 & N4766;
  assign N2094 = N4746 & N4767;
  assign N4747 = addr_i[6] & N4772;
  assign N4748 = N4768 & N4769;
  assign N4749 = N4768 & N4770;
  assign N4750 = N4768 & N4771;
  assign N4751 = N4768 & N4772;
  assign N4752 = N4781 & N4785;
  assign N4753 = N4781 & N4786;
  assign N4754 = N4781 & N4787;
  assign N4755 = N4781 & N4788;
  assign N4756 = N4782 & N4785;
  assign N4757 = N4782 & N4786;
  assign N4758 = N4782 & N4787;
  assign N4759 = N4782 & N4788;
  assign N4760 = N4783 & N4785;
  assign N4761 = N4783 & N4786;
  assign N4762 = N4783 & N4787;
  assign N4763 = N4783 & N4788;
  assign N4764 = N4784 & N4785;
  assign N4765 = N4784 & N4786;
  assign N4766 = N4784 & N4787;
  assign N4767 = N4784 & N4788;
  assign N2430 = N4773 & N4752;
  assign N2429 = N4773 & N4753;
  assign N2428 = N4773 & N4754;
  assign N2427 = N4773 & N4755;
  assign N2426 = N4773 & N4756;
  assign N2425 = N4773 & N4757;
  assign N2424 = N4773 & N4758;
  assign N2423 = N4773 & N4759;
  assign N2422 = N4773 & N4760;
  assign N2421 = N4773 & N4761;
  assign N2420 = N4773 & N4762;
  assign N2419 = N4773 & N4763;
  assign N2418 = N4773 & N4764;
  assign N2417 = N4773 & N4765;
  assign N2416 = N4773 & N4766;
  assign N2415 = N4773 & N4767;
  assign N2414 = N4774 & N4752;
  assign N2413 = N4774 & N4753;
  assign N2412 = N4774 & N4754;
  assign N2411 = N4774 & N4755;
  assign N2410 = N4774 & N4756;
  assign N2409 = N4774 & N4757;
  assign N2408 = N4774 & N4758;
  assign N2407 = N4774 & N4759;
  assign N2406 = N4774 & N4760;
  assign N2405 = N4774 & N4761;
  assign N2404 = N4774 & N4762;
  assign N2403 = N4774 & N4763;
  assign N2402 = N4774 & N4764;
  assign N2401 = N4774 & N4765;
  assign N2400 = N4774 & N4766;
  assign N2399 = N4774 & N4767;
  assign N2398 = N4775 & N4752;
  assign N2397 = N4775 & N4753;
  assign N2396 = N4775 & N4754;
  assign N2395 = N4775 & N4755;
  assign N2394 = N4775 & N4756;
  assign N2393 = N4775 & N4757;
  assign N2392 = N4775 & N4758;
  assign N2391 = N4775 & N4759;
  assign N2390 = N4775 & N4760;
  assign N2389 = N4775 & N4761;
  assign N2388 = N4775 & N4762;
  assign N2387 = N4775 & N4763;
  assign N2386 = N4775 & N4764;
  assign N2385 = N4775 & N4765;
  assign N2384 = N4775 & N4766;
  assign N2383 = N4775 & N4767;
  assign N2382 = N4747 & N4752;
  assign N2381 = N4747 & N4753;
  assign N2380 = N4747 & N4754;
  assign N2379 = N4747 & N4755;
  assign N2378 = N4747 & N4756;
  assign N2377 = N4747 & N4757;
  assign N2376 = N4747 & N4758;
  assign N2375 = N4747 & N4759;
  assign N2374 = N4747 & N4760;
  assign N2373 = N4747 & N4761;
  assign N2372 = N4747 & N4762;
  assign N2371 = N4747 & N4763;
  assign N2370 = N4747 & N4764;
  assign N2369 = N4747 & N4765;
  assign N2368 = N4747 & N4766;
  assign N2367 = N4747 & N4767;
  assign N2366 = N4748 & N4752;
  assign N2365 = N4748 & N4753;
  assign N2364 = N4748 & N4754;
  assign N2363 = N4748 & N4755;
  assign N2362 = N4748 & N4756;
  assign N2361 = N4748 & N4757;
  assign N2360 = N4748 & N4758;
  assign N2359 = N4748 & N4759;
  assign N2358 = N4748 & N4760;
  assign N2357 = N4748 & N4761;
  assign N2356 = N4748 & N4762;
  assign N2355 = N4748 & N4763;
  assign N2354 = N4748 & N4764;
  assign N2353 = N4748 & N4765;
  assign N2352 = N4748 & N4766;
  assign N2351 = N4748 & N4767;
  assign N2350 = N4749 & N4752;
  assign N2349 = N4749 & N4753;
  assign N2348 = N4749 & N4754;
  assign N2347 = N4749 & N4755;
  assign N2346 = N4749 & N4756;
  assign N2345 = N4749 & N4757;
  assign N2344 = N4749 & N4758;
  assign N2343 = N4749 & N4759;
  assign N2342 = N4749 & N4760;
  assign N2341 = N4749 & N4761;
  assign N2340 = N4749 & N4762;
  assign N2339 = N4749 & N4763;
  assign N2338 = N4749 & N4764;
  assign N2337 = N4749 & N4765;
  assign N2336 = N4749 & N4766;
  assign N2335 = N4749 & N4767;
  assign N2334 = N4750 & N4752;
  assign N2333 = N4750 & N4753;
  assign N2332 = N4750 & N4754;
  assign N2331 = N4750 & N4755;
  assign N2330 = N4750 & N4756;
  assign N2329 = N4750 & N4757;
  assign N2328 = N4750 & N4758;
  assign N2327 = N4750 & N4759;
  assign N2326 = N4750 & N4760;
  assign N2325 = N4750 & N4761;
  assign N2324 = N4750 & N4762;
  assign N2323 = N4750 & N4763;
  assign N2322 = N4750 & N4764;
  assign N2321 = N4750 & N4765;
  assign N2320 = N4750 & N4766;
  assign N2319 = N4750 & N4767;
  assign N2318 = N4751 & N4752;
  assign N2317 = N4751 & N4753;
  assign N2316 = N4751 & N4754;
  assign N2315 = N4751 & N4755;
  assign N2314 = N4751 & N4756;
  assign N2313 = N4751 & N4757;
  assign N2312 = N4751 & N4758;
  assign N2311 = N4751 & N4759;
  assign N2310 = N4751 & N4760;
  assign N2309 = N4751 & N4761;
  assign N2308 = N4751 & N4762;
  assign N2307 = N4751 & N4763;
  assign N2306 = N4751 & N4764;
  assign N2305 = N4751 & N4765;
  assign N2304 = N4751 & N4766;
  assign N2303 = N4751 & N4767;
  assign N4768 = ~addr_i[6];
  assign N4769 = addr_i[4] & addr_i[5];
  assign N4770 = N0 & addr_i[5];
  assign N0 = ~addr_i[4];
  assign N4771 = addr_i[4] & N1;
  assign N1 = ~addr_i[5];
  assign N4772 = N2 & N3;
  assign N2 = ~addr_i[4];
  assign N3 = ~addr_i[5];
  assign N4773 = addr_i[6] & N4769;
  assign N4774 = addr_i[6] & N4770;
  assign N4775 = addr_i[6] & N4771;
  assign N4776 = addr_i[6] & N4772;
  assign N4777 = N4768 & N4769;
  assign N4778 = N4768 & N4770;
  assign N4779 = N4768 & N4771;
  assign N4780 = N4768 & N4772;
  assign N4781 = addr_i[2] & addr_i[3];
  assign N4782 = N4 & addr_i[3];
  assign N4 = ~addr_i[2];
  assign N4783 = addr_i[2] & N5;
  assign N5 = ~addr_i[3];
  assign N4784 = N6 & N7;
  assign N6 = ~addr_i[2];
  assign N7 = ~addr_i[3];
  assign N4785 = addr_i[0] & addr_i[1];
  assign N4786 = N8 & addr_i[1];
  assign N8 = ~addr_i[0];
  assign N4787 = addr_i[0] & N9;
  assign N9 = ~addr_i[1];
  assign N4788 = N10 & N11;
  assign N10 = ~addr_i[0];
  assign N11 = ~addr_i[1];
  assign N4789 = N4781 & N4785;
  assign N4790 = N4781 & N4786;
  assign N4791 = N4781 & N4787;
  assign N4792 = N4781 & N4788;
  assign N4793 = N4782 & N4785;
  assign N4794 = N4782 & N4786;
  assign N4795 = N4782 & N4787;
  assign N4796 = N4782 & N4788;
  assign N4797 = N4783 & N4785;
  assign N4798 = N4783 & N4786;
  assign N4799 = N4783 & N4787;
  assign N4800 = N4783 & N4788;
  assign N4801 = N4784 & N4785;
  assign N4802 = N4784 & N4786;
  assign N4803 = N4784 & N4787;
  assign N4804 = N4784 & N4788;
  assign N2687 = N4773 & N4789;
  assign N2686 = N4773 & N4790;
  assign N2685 = N4773 & N4791;
  assign N2684 = N4773 & N4792;
  assign N2683 = N4773 & N4793;
  assign N2682 = N4773 & N4794;
  assign N2681 = N4773 & N4795;
  assign N2680 = N4773 & N4796;
  assign N2679 = N4773 & N4797;
  assign N2678 = N4773 & N4798;
  assign N2677 = N4773 & N4799;
  assign N2676 = N4773 & N4800;
  assign N2675 = N4773 & N4801;
  assign N2674 = N4773 & N4802;
  assign N2673 = N4773 & N4803;
  assign N2672 = N4773 & N4804;
  assign N2671 = N4774 & N4789;
  assign N2670 = N4774 & N4790;
  assign N2669 = N4774 & N4791;
  assign N2668 = N4774 & N4792;
  assign N2667 = N4774 & N4793;
  assign N2666 = N4774 & N4794;
  assign N2665 = N4774 & N4795;
  assign N2664 = N4774 & N4796;
  assign N2663 = N4774 & N4797;
  assign N2662 = N4774 & N4798;
  assign N2661 = N4774 & N4799;
  assign N2660 = N4774 & N4800;
  assign N2659 = N4774 & N4801;
  assign N2658 = N4774 & N4802;
  assign N2657 = N4774 & N4803;
  assign N2656 = N4774 & N4804;
  assign N2655 = N4775 & N4789;
  assign N2654 = N4775 & N4790;
  assign N2653 = N4775 & N4791;
  assign N2652 = N4775 & N4792;
  assign N2651 = N4775 & N4793;
  assign N2650 = N4775 & N4794;
  assign N2649 = N4775 & N4795;
  assign N2648 = N4775 & N4796;
  assign N2647 = N4775 & N4797;
  assign N2646 = N4775 & N4798;
  assign N2645 = N4775 & N4799;
  assign N2644 = N4775 & N4800;
  assign N2643 = N4775 & N4801;
  assign N2642 = N4775 & N4802;
  assign N2641 = N4775 & N4803;
  assign N2640 = N4775 & N4804;
  assign N2639 = N4776 & N4789;
  assign N2638 = N4776 & N4790;
  assign N2637 = N4776 & N4791;
  assign N2636 = N4776 & N4792;
  assign N2635 = N4776 & N4793;
  assign N2634 = N4776 & N4794;
  assign N2633 = N4776 & N4795;
  assign N2632 = N4776 & N4796;
  assign N2631 = N4776 & N4797;
  assign N2630 = N4776 & N4798;
  assign N2629 = N4776 & N4799;
  assign N2628 = N4776 & N4800;
  assign N2627 = N4776 & N4801;
  assign N2626 = N4776 & N4802;
  assign N2625 = N4776 & N4803;
  assign N2624 = N4776 & N4804;
  assign N2623 = N4777 & N4789;
  assign N2622 = N4777 & N4790;
  assign N2621 = N4777 & N4791;
  assign N2620 = N4777 & N4792;
  assign N2619 = N4777 & N4793;
  assign N2618 = N4777 & N4794;
  assign N2617 = N4777 & N4795;
  assign N2616 = N4777 & N4796;
  assign N2615 = N4777 & N4797;
  assign N2614 = N4777 & N4798;
  assign N2613 = N4777 & N4799;
  assign N2612 = N4777 & N4800;
  assign N2611 = N4777 & N4801;
  assign N2610 = N4777 & N4802;
  assign N2609 = N4777 & N4803;
  assign N2608 = N4777 & N4804;
  assign N2607 = N4778 & N4789;
  assign N2606 = N4778 & N4790;
  assign N2605 = N4778 & N4791;
  assign N2604 = N4778 & N4792;
  assign N2603 = N4778 & N4793;
  assign N2602 = N4778 & N4794;
  assign N2601 = N4778 & N4795;
  assign N2600 = N4778 & N4796;
  assign N2599 = N4778 & N4797;
  assign N2598 = N4778 & N4798;
  assign N2597 = N4778 & N4799;
  assign N2596 = N4778 & N4800;
  assign N2595 = N4778 & N4801;
  assign N2594 = N4778 & N4802;
  assign N2593 = N4778 & N4803;
  assign N2592 = N4778 & N4804;
  assign N2591 = N4779 & N4789;
  assign N2590 = N4779 & N4790;
  assign N2589 = N4779 & N4791;
  assign N2588 = N4779 & N4792;
  assign N2587 = N4779 & N4793;
  assign N2586 = N4779 & N4794;
  assign N2585 = N4779 & N4795;
  assign N2584 = N4779 & N4796;
  assign N2583 = N4779 & N4797;
  assign N2582 = N4779 & N4798;
  assign N2581 = N4779 & N4799;
  assign N2580 = N4779 & N4800;
  assign N2579 = N4779 & N4801;
  assign N2578 = N4779 & N4802;
  assign N2577 = N4779 & N4803;
  assign N2576 = N4779 & N4804;
  assign N2575 = N4780 & N4789;
  assign N2574 = N4780 & N4790;
  assign N2573 = N4780 & N4791;
  assign N2572 = N4780 & N4792;
  assign N2571 = N4780 & N4793;
  assign N2570 = N4780 & N4794;
  assign N2569 = N4780 & N4795;
  assign N2568 = N4780 & N4796;
  assign N2567 = N4780 & N4797;
  assign N2566 = N4780 & N4798;
  assign N2565 = N4780 & N4799;
  assign N2564 = N4780 & N4800;
  assign N2563 = N4780 & N4801;
  assign N2562 = N4780 & N4802;
  assign N2561 = N4780 & N4803;
  assign N2560 = N4780 & N4804;
  assign { N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290 } = (N12)? { N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N289)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[0];
  assign { N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419 } = (N13)? { N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N418)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[1];
  assign { N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596 } = (N14)? { N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N547)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[2];
  assign { N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725 } = (N15)? { N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N724)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = w_mask_i[3];
  assign { N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854 } = (N16)? { N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N853)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_mask_i[4];
  assign { N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983 } = (N17)? { N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             (N982)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = w_mask_i[5];
  assign { N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112 } = (N18)? { N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1111)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = w_mask_i[6];
  assign { N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241 } = (N19)? { N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1240)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = w_mask_i[7];
  assign { N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418 } = (N20)? { N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1369)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = w_mask_i[8];
  assign { N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627 } = (N21)? { N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1546)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = w_mask_i[9];
  assign { N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836 } = (N22)? { N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1755)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = w_mask_i[10];
  assign { N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965 } = (N23)? { N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1964)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = w_mask_i[11];
  assign { N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174 } = (N24)? { N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2093)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N24 = w_mask_i[12];
  assign { N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431 } = (N25)? { N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2302)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = w_mask_i[13];
  assign { N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688 } = (N26)? { N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2559)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = w_mask_i[14];
  assign { N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073, N4072, N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251, N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N3226, N3225, N3224, N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816 } = (N27)? { N2815, N2558, N2301, N2092, N1963, N1754, N1545, N1368, N1239, N1110, N981, N852, N723, N546, N417, N2814, N2557, N2300, N2091, N1962, N1753, N1544, N1367, N1238, N1109, N980, N851, N722, N545, N416, N2813, N2556, N2299, N2090, N1961, N1752, N1543, N1366, N1237, N1108, N979, N850, N721, N544, N415, N2812, N2555, N2298, N2089, N1960, N1751, N1542, N1365, N1236, N1107, N978, N849, N720, N543, N414, N2811, N2554, N2297, N2088, N1959, N1750, N1541, N1364, N1235, N1106, N977, N848, N719, N542, N413, N2810, N2553, N2296, N2087, N1958, N1749, N1540, N1363, N1234, N1105, N976, N847, N718, N541, N412, N2809, N2552, N2295, N2086, N1957, N1748, N1539, N1362, N1233, N1104, N975, N846, N717, N540, N411, N2808, N2551, N2294, N2085, N1956, N1747, N1538, N1361, N1232, N1103, N974, N845, N716, N539, N410, N2807, N2550, N2293, N2084, N1955, N1746, N1537, N1360, N1231, N1102, N973, N844, N715, N538, N409, N2806, N2549, N2292, N2083, N1954, N1745, N1536, N1359, N1230, N1101, N972, N843, N714, N537, N408, N2805, N2548, N2291, N2082, N1953, N1744, N1535, N1358, N1229, N1100, N971, N842, N713, N536, N407, N2804, N2547, N2290, N2081, N1952, N1743, N1534, N1357, N1228, N1099, N970, N841, N712, N535, N406, N2803, N2546, N2289, N2080, N1951, N1742, N1533, N1356, N1227, N1098, N969, N840, N711, N534, N405, N2802, N2545, N2288, N2079, N1950, N1741, N1532, N1355, N1226, N1097, N968, N839, N710, N533, N404, N2801, N2544, N2287, N2078, N1949, N1740, N1531, N1354, N1225, N1096, N967, N838, N709, N532, N403, N2800, N2543, N2286, N2077, N1948, N1739, N1530, N1353, N1224, N1095, N966, N837, N708, N531, N402, N2799, N2542, N2285, N2076, N1947, N1738, N1529, N1352, N1223, N1094, N965, N836, N707, N530, N401, N2798, N2541, N2284, N2075, N1946, N1737, N1528, N1351, N1222, N1093, N964, N835, N706, N529, N400, N2797, N2540, N2283, N2074, N1945, N1736, N1527, N1350, N1221, N1092, N963, N834, N705, N528, N399, N2796, N2539, N2282, N2073, N1944, N1735, N1526, N1349, N1220, N1091, N962, N833, N704, N527, N398, N2795, N2538, N2281, N2072, N1943, N1734, N1525, N1348, N1219, N1090, N961, N832, N703, N526, N397, N2794, N2537, N2280, N2071, N1942, N1733, N1524, N1347, N1218, N1089, N960, N831, N702, N525, N396, N2793, N2536, N2279, N2070, N1941, N1732, N1523, N1346, N1217, N1088, N959, N830, N701, N524, N395, N2792, N2535, N2278, N2069, N1940, N1731, N1522, N1345, N1216, N1087, N958, N829, N700, N523, N394, N2791, N2534, N2277, N2068, N1939, N1730, N1521, N1344, N1215, N1086, N957, N828, N699, N522, N393, N2790, N2533, N2276, N2067, N1938, N1729, N1520, N1343, N1214, N1085, N956, N827, N698, N521, N392, N2789, N2532, N2275, N2066, N1937, N1728, N1519, N1342, N1213, N1084, N955, N826, N697, N520, N391, N2788, N2531, N2274, N2065, N1936, N1727, N1518, N1341, N1212, N1083, N954, N825, N696, N519, N390, N2787, N2530, N2273, N2064, N1935, N1726, N1517, N1340, N1211, N1082, N953, N824, N695, N518, N389, N2786, N2529, N2272, N2063, N1934, N1725, N1516, N1339, N1210, N1081, N952, N823, N694, N517, N388, N2785, N2528, N2271, N2062, N1933, N1724, N1515, N1338, N1209, N1080, N951, N822, N693, N516, N387, N2784, N2527, N2270, N2061, N1932, N1723, N1514, N1337, N1208, N1079, N950, N821, N692, N515, N386, N2783, N2526, N2269, N2060, N1931, N1722, N1513, N1336, N1207, N1078, N949, N820, N691, N514, N385, N2782, N2525, N2268, N2059, N1930, N1721, N1512, N1335, N1206, N1077, N948, N819, N690, N513, N384, N2781, N2524, N2267, N2058, N1929, N1720, N1511, N1334, N1205, N1076, N947, N818, N689, N512, N383, N2780, N2523, N2266, N2057, N1928, N1719, N1510, N1333, N1204, N1075, N946, N817, N688, N511, N382, N2779, N2522, N2265, N2056, N1927, N1718, N1509, N1332, N1203, N1074, N945, N816, N687, N510, N381, N2778, N2521, N2264, N2055, N1926, N1717, N1508, N1331, N1202, N1073, N944, N815, N686, N509, N380, N2777, N2520, N2263, N2054, N1925, N1716, N1507, N1330, N1201, N1072, N943, N814, N685, N508, N379, N2776, N2519, N2262, N2053, N1924, N1715, N1506, N1329, N1200, N1071, N942, N813, N684, N507, N378, N2775, N2518, N2261, N2052, N1923, N1714, N1505, N1328, N1199, N1070, N941, N812, N683, N506, N377, N2774, N2517, N2260, N2051, N1922, N1713, N1504, N1327, N1198, N1069, N940, N811, N682, N505, N376, N2773, N2516, N2259, N2050, N1921, N1712, N1503, N1326, N1197, N1068, N939, N810, N681, N504, N375, N2772, N2515, N2258, N2049, N1920, N1711, N1502, N1325, N1196, N1067, N938, N809, N680, N503, N374, N2771, N2514, N2257, N2048, N1919, N1710, N1501, N1324, N1195, N1066, N937, N808, N679, N502, N373, N2770, N2513, N2256, N2047, N1918, N1709, N1500, N1323, N1194, N1065, N936, N807, N678, N501, N372, N2769, N2512, N2255, N2046, N1917, N1708, N1499, N1322, N1193, N1064, N935, N806, N677, N500, N371, N2768, N2511, N2254, N2045, N1916, N1707, N1498, N1321, N1192, N1063, N934, N805, N676, N499, N370, N2767, N2510, N2253, N2044, N1915, N1706, N1497, N1320, N1191, N1062, N933, N804, N675, N498, N369, N2766, N2509, N2252, N2043, N1914, N1705, N1496, N1319, N1190, N1061, N932, N803, N674, N497, N368, N2765, N2508, N2251, N2042, N1913, N1704, N1495, N1318, N1189, N1060, N931, N802, N673, N496, N367, N2764, N2507, N2250, N2041, N1912, N1703, N1494, N1317, N1188, N1059, N930, N801, N672, N495, N366, N2763, N2506, N2249, N2040, N1911, N1702, N1493, N1316, N1187, N1058, N929, N800, N671, N494, N365, N2762, N2505, N2248, N2039, N1910, N1701, N1492, N1315, N1186, N1057, N928, N799, N670, N493, N364, N2761, N2504, N2247, N2038, N1909, N1700, N1491, N1314, N1185, N1056, N927, N798, N669, N492, N363, N2760, N2503, N2246, N2037, N1908, N1699, N1490, N1313, N1184, N1055, N926, N797, N668, N491, N362, N2759, N2502, N2245, N2036, N1907, N1698, N1489, N1312, N1183, N1054, N925, N796, N667, N490, N361, N2758, N2501, N2244, N2035, N1906, N1697, N1488, N1311, N1182, N1053, N924, N795, N666, N489, N360, N2757, N2500, N2243, N2034, N1905, N1696, N1487, N1310, N1181, N1052, N923, N794, N665, N488, N359, N2756, N2499, N2242, N2033, N1904, N1695, N1486, N1309, N1180, N1051, N922, N793, N664, N487, N358, N2755, N2498, N2241, N2032, N1903, N1694, N1485, N1308, N1179, N1050, N921, N792, N663, N486, N357, N2754, N2497, N2240, N2031, N1902, N1693, N1484, N1307, N1178, N1049, N920, N791, N662, N485, N356, N2753, N2496, N2239, N2030, N1901, N1692, N1483, N1306, N1177, N1048, N919, N790, N661, N484, N355, N2752, N2495, N2238, N2029, N1900, N1691, N1482, N1305, N1176, N1047, N918, N789, N660, N483, N354, N2751, N2494, N2237, N2028, N1899, N1690, N1481, N1304, N1175, N1046, N917, N788, N659, N482, N353, N2750, N2493, N2236, N2027, N1898, N1689, N1480, N1303, N1174, N1045, N916, N787, N658, N481, N352, N2749, N2492, N2235, N2026, N1897, N1688, N1479, N1302, N1173, N1044, N915, N786, N657, N480, N351, N2748, N2491, N2234, N2025, N1896, N1687, N1478, N1301, N1172, N1043, N914, N785, N656, N479, N350, N2747, N2490, N2233, N2024, N1895, N1686, N1477, N1300, N1171, N1042, N913, N784, N655, N478, N349, N2746, N2489, N2232, N2023, N1894, N1685, N1476, N1299, N1170, N1041, N912, N783, N654, N477, N348, N2745, N2488, N2231, N2022, N1893, N1684, N1475, N1298, N1169, N1040, N911, N782, N653, N476, N347, N2744, N2487, N2230, N2021, N1892, N1683, N1474, N1297, N1168, N1039, N910, N781, N652, N475, N346, N2743, N2486, N2229, N2020, N1891, N1682, N1473, N1296, N1167, N1038, N909, N780, N651, N474, N345, N2742, N2485, N2228, N2019, N1890, N1681, N1472, N1295, N1166, N1037, N908, N779, N650, N473, N344, N2741, N2484, N2227, N2018, N1889, N1680, N1471, N1294, N1165, N1036, N907, N778, N649, N472, N343, N2740, N2483, N2226, N2017, N1888, N1679, N1470, N1293, N1164, N1035, N906, N777, N648, N471, N342, N2739, N2482, N2225, N2016, N1887, N1678, N1469, N1292, N1163, N1034, N905, N776, N647, N470, N341, N2738, N2481, N2224, N2015, N1886, N1677, N1468, N1291, N1162, N1033, N904, N775, N646, N469, N340, N2737, N2480, N2223, N2014, N1885, N1676, N1467, N1290, N1161, N1032, N903, N774, N645, N468, N339, N2736, N2479, N2222, N2013, N1884, N1675, N1466, N1289, N1160, N1031, N902, N773, N644, N467, N338, N2735, N2478, N2221, N2012, N1883, N1674, N1465, N1288, N1159, N1030, N901, N772, N643, N466, N337, N2734, N2477, N2220, N2011, N1882, N1673, N1464, N1287, N1158, N1029, N900, N771, N642, N465, N336, N2733, N2476, N2219, N2010, N1881, N1672, N1463, N1286, N1157, N1028, N899, N770, N641, N464, N335, N2732, N2475, N2218, N2009, N1880, N1671, N1462, N1285, N1156, N1027, N898, N769, N640, N463, N334, N2731, N2474, N2217, N2008, N1879, N1670, N1461, N1284, N1155, N1026, N897, N768, N639, N462, N333, N2730, N2473, N2216, N2007, N1878, N1669, N1460, N1283, N1154, N1025, N896, N767, N638, N461, N332, N2729, N2472, N2215, N2006, N1877, N1668, N1459, N1282, N1153, N1024, N895, N766, N637, N460, N331, N2728, N2471, N2214, N2005, N1876, N1667, N1458, N1281, N1152, N1023, N894, N765, N636, N459, N330, N2727, N2470, N2213, N2004, N1875, N1666, N1457, N1280, N1151, N1022, N893, N764, N635, N458, N329, N2726, N2469, N2212, N2003, N1874, N1665, N1456, N1279, N1150, N1021, N892, N763, N634, N457, N328, N2725, N2468, N2211, N2002, N1873, N1664, N1455, N1278, N1149, N1020, N891, N762, N633, N456, N327, N2724, N2467, N2210, N2001, N1872, N1663, N1454, N1277, N1148, N1019, N890, N761, N632, N455, N326, N2723, N2466, N2209, N2000, N1871, N1662, N1453, N1276, N1147, N1018, N889, N760, N631, N454, N325, N2722, N2465, N2208, N1999, N1870, N1661, N1452, N1275, N1146, N1017, N888, N759, N630, N453, N324, N2721, N2464, N2207, N1998, N1869, N1660, N1451, N1274, N1145, N1016, N887, N758, N629, N452, N323, N2720, N2463, N2206, N1997, N1868, N1659, N1450, N1273, N1144, N1015, N886, N757, N628, N451, N322, N2719, N2462, N2205, N1996, N1867, N1658, N1449, N1272, N1143, N1014, N885, N756, N627, N450, N321, N2718, N2461, N2204, N1995, N1866, N1657, N1448, N1271, N1142, N1013, N884, N755, N626, N449, N320, N2717, N2460, N2203, N1994, N1865, N1656, N1447, N1270, N1141, N1012, N883, N754, N625, N448, N319, N2716, N2459, N2202, N1993, N1864, N1655, N1446, N1269, N1140, N1011, N882, N753, N624, N447, N318, N2715, N2458, N2201, N1992, N1863, N1654, N1445, N1268, N1139, N1010, N881, N752, N623, N446, N317, N2714, N2457, N2200, N1991, N1862, N1653, N1444, N1267, N1138, N1009, N880, N751, N622, N445, N316, N2713, N2456, N2199, N1990, N1861, N1652, N1443, N1266, N1137, N1008, N879, N750, N621, N444, N315, N2712, N2455, N2198, N1989, N1860, N1651, N1442, N1265, N1136, N1007, N878, N749, N620, N443, N314, N2711, N2454, N2197, N1988, N1859, N1650, N1441, N1264, N1135, N1006, N877, N748, N619, N442, N313, N2710, N2453, N2196, N1987, N1858, N1649, N1440, N1263, N1134, N1005, N876, N747, N618, N441, N312, N2709, N2452, N2195, N1986, N1857, N1648, N1439, N1262, N1133, N1004, N875, N746, N617, N440, N311, N2708, N2451, N2194, N1985, N1856, N1647, N1438, N1261, N1132, N1003, N874, N745, N616, N439, N310, N2707, N2450, N2193, N1984, N1855, N1646, N1437, N1260, N1131, N1002, N873, N744, N615, N438, N309, N2706, N2449, N2192, N1983, N1854, N1645, N1436, N1259, N1130, N1001, N872, N743, N614, N437, N308, N2705, N2448, N2191, N1982, N1853, N1644, N1435, N1258, N1129, N1000, N871, N742, N613, N436, N307, N2704, N2447, N2190, N1981, N1852, N1643, N1434, N1257, N1128, N999, N870, N741, N612, N435, N306, N2703, N2446, N2189, N1980, N1851, N1642, N1433, N1256, N1127, N998, N869, N740, N611, N434, N305, N2702, N2445, N2188, N1979, N1850, N1641, N1432, N1255, N1126, N997, N868, N739, N610, N433, N304, N2701, N2444, N2187, N1978, N1849, N1640, N1431, N1254, N1125, N996, N867, N738, N609, N432, N303, N2700, N2443, N2186, N1977, N1848, N1639, N1430, N1253, N1124, N995, N866, N737, N608, N431, N302, N2699, N2442, N2185, N1976, N1847, N1638, N1429, N1252, N1123, N994, N865, N736, N607, N430, N301, N2698, N2441, N2184, N1975, N1846, N1637, N1428, N1251, N1122, N993, N864, N735, N606, N429, N300, N2697, N2440, N2183, N1974, N1845, N1636, N1427, N1250, N1121, N992, N863, N734, N605, N428, N299, N2696, N2439, N2182, N1973, N1844, N1635, N1426, N1249, N1120, N991, N862, N733, N604, N427, N298, N2695, N2438, N2181, N1972, N1843, N1634, N1425, N1248, N1119, N990, N861, N732, N603, N426, N297, N2694, N2437, N2180, N1971, N1842, N1633, N1424, N1247, N1118, N989, N860, N731, N602, N425, N296, N2693, N2436, N2179, N1970, N1841, N1632, N1423, N1246, N1117, N988, N859, N730, N601, N424, N295, N2692, N2435, N2178, N1969, N1840, N1631, N1422, N1245, N1116, N987, N858, N729, N600, N423, N294, N2691, N2434, N2177, N1968, N1839, N1630, N1421, N1244, N1115, N986, N857, N728, N599, N422, N293, N2690, N2433, N2176, N1967, N1838, N1629, N1420, N1243, N1114, N985, N856, N727, N598, N421, N292, N2689, N2432, N2175, N1966, N1837, N1628, N1419, N1242, N1113, N984, N855, N726, N597, N420, N291, N2688, N2431, N2174, N1965, N1836, N1627, N1418, N1241, N1112, N983, N854, N725, N596, N419, N290 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N288)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N27 = N287;
  assign N28 = ~addr_r[0];
  assign N29 = ~addr_r[1];
  assign N30 = N28 & N29;
  assign N31 = N28 & addr_r[1];
  assign N32 = addr_r[0] & N29;
  assign N33 = addr_r[0] & addr_r[1];
  assign N34 = ~addr_r[2];
  assign N35 = N30 & N34;
  assign N36 = N30 & addr_r[2];
  assign N37 = N32 & N34;
  assign N38 = N32 & addr_r[2];
  assign N39 = N31 & N34;
  assign N40 = N31 & addr_r[2];
  assign N41 = N33 & N34;
  assign N42 = N33 & addr_r[2];
  assign N43 = ~addr_r[3];
  assign N44 = N35 & N43;
  assign N45 = N35 & addr_r[3];
  assign N46 = N37 & N43;
  assign N47 = N37 & addr_r[3];
  assign N48 = N39 & N43;
  assign N49 = N39 & addr_r[3];
  assign N50 = N41 & N43;
  assign N51 = N41 & addr_r[3];
  assign N52 = N36 & N43;
  assign N53 = N36 & addr_r[3];
  assign N54 = N38 & N43;
  assign N55 = N38 & addr_r[3];
  assign N56 = N40 & N43;
  assign N57 = N40 & addr_r[3];
  assign N58 = N42 & N43;
  assign N59 = N42 & addr_r[3];
  assign N60 = ~addr_r[4];
  assign N61 = N44 & N60;
  assign N62 = N44 & addr_r[4];
  assign N63 = N46 & N60;
  assign N64 = N46 & addr_r[4];
  assign N65 = N48 & N60;
  assign N66 = N48 & addr_r[4];
  assign N67 = N50 & N60;
  assign N68 = N50 & addr_r[4];
  assign N69 = N52 & N60;
  assign N70 = N52 & addr_r[4];
  assign N71 = N54 & N60;
  assign N72 = N54 & addr_r[4];
  assign N73 = N56 & N60;
  assign N74 = N56 & addr_r[4];
  assign N75 = N58 & N60;
  assign N76 = N58 & addr_r[4];
  assign N77 = N45 & N60;
  assign N78 = N45 & addr_r[4];
  assign N79 = N47 & N60;
  assign N80 = N47 & addr_r[4];
  assign N81 = N49 & N60;
  assign N82 = N49 & addr_r[4];
  assign N83 = N51 & N60;
  assign N84 = N51 & addr_r[4];
  assign N85 = N53 & N60;
  assign N86 = N53 & addr_r[4];
  assign N87 = N55 & N60;
  assign N88 = N55 & addr_r[4];
  assign N89 = N57 & N60;
  assign N90 = N57 & addr_r[4];
  assign N91 = N59 & N60;
  assign N92 = N59 & addr_r[4];
  assign N93 = ~addr_r[5];
  assign N94 = N61 & N93;
  assign N95 = N61 & addr_r[5];
  assign N96 = N63 & N93;
  assign N97 = N63 & addr_r[5];
  assign N98 = N65 & N93;
  assign N99 = N65 & addr_r[5];
  assign N100 = N67 & N93;
  assign N101 = N67 & addr_r[5];
  assign N102 = N69 & N93;
  assign N103 = N69 & addr_r[5];
  assign N104 = N71 & N93;
  assign N105 = N71 & addr_r[5];
  assign N106 = N73 & N93;
  assign N107 = N73 & addr_r[5];
  assign N108 = N75 & N93;
  assign N109 = N75 & addr_r[5];
  assign N110 = N77 & N93;
  assign N111 = N77 & addr_r[5];
  assign N112 = N79 & N93;
  assign N113 = N79 & addr_r[5];
  assign N114 = N81 & N93;
  assign N115 = N81 & addr_r[5];
  assign N116 = N83 & N93;
  assign N117 = N83 & addr_r[5];
  assign N118 = N85 & N93;
  assign N119 = N85 & addr_r[5];
  assign N120 = N87 & N93;
  assign N121 = N87 & addr_r[5];
  assign N122 = N89 & N93;
  assign N123 = N89 & addr_r[5];
  assign N124 = N91 & N93;
  assign N125 = N91 & addr_r[5];
  assign N126 = N62 & N93;
  assign N127 = N62 & addr_r[5];
  assign N128 = N64 & N93;
  assign N129 = N64 & addr_r[5];
  assign N130 = N66 & N93;
  assign N131 = N66 & addr_r[5];
  assign N132 = N68 & N93;
  assign N133 = N68 & addr_r[5];
  assign N134 = N70 & N93;
  assign N135 = N70 & addr_r[5];
  assign N136 = N72 & N93;
  assign N137 = N72 & addr_r[5];
  assign N138 = N74 & N93;
  assign N139 = N74 & addr_r[5];
  assign N140 = N76 & N93;
  assign N141 = N76 & addr_r[5];
  assign N142 = N78 & N93;
  assign N143 = N78 & addr_r[5];
  assign N144 = N80 & N93;
  assign N145 = N80 & addr_r[5];
  assign N146 = N82 & N93;
  assign N147 = N82 & addr_r[5];
  assign N148 = N84 & N93;
  assign N149 = N84 & addr_r[5];
  assign N150 = N86 & N93;
  assign N151 = N86 & addr_r[5];
  assign N152 = N88 & N93;
  assign N153 = N88 & addr_r[5];
  assign N154 = N90 & N93;
  assign N155 = N90 & addr_r[5];
  assign N156 = N92 & N93;
  assign N157 = N92 & addr_r[5];
  assign N158 = ~addr_r[6];
  assign N159 = N94 & N158;
  assign N160 = N94 & addr_r[6];
  assign N161 = N96 & N158;
  assign N162 = N96 & addr_r[6];
  assign N163 = N98 & N158;
  assign N164 = N98 & addr_r[6];
  assign N165 = N100 & N158;
  assign N166 = N100 & addr_r[6];
  assign N167 = N102 & N158;
  assign N168 = N102 & addr_r[6];
  assign N169 = N104 & N158;
  assign N170 = N104 & addr_r[6];
  assign N171 = N106 & N158;
  assign N172 = N106 & addr_r[6];
  assign N173 = N108 & N158;
  assign N174 = N108 & addr_r[6];
  assign N175 = N110 & N158;
  assign N176 = N110 & addr_r[6];
  assign N177 = N112 & N158;
  assign N178 = N112 & addr_r[6];
  assign N179 = N114 & N158;
  assign N180 = N114 & addr_r[6];
  assign N181 = N116 & N158;
  assign N182 = N116 & addr_r[6];
  assign N183 = N118 & N158;
  assign N184 = N118 & addr_r[6];
  assign N185 = N120 & N158;
  assign N186 = N120 & addr_r[6];
  assign N187 = N122 & N158;
  assign N188 = N122 & addr_r[6];
  assign N189 = N124 & N158;
  assign N190 = N124 & addr_r[6];
  assign N191 = N126 & N158;
  assign N192 = N126 & addr_r[6];
  assign N193 = N128 & N158;
  assign N194 = N128 & addr_r[6];
  assign N195 = N130 & N158;
  assign N196 = N130 & addr_r[6];
  assign N197 = N132 & N158;
  assign N198 = N132 & addr_r[6];
  assign N199 = N134 & N158;
  assign N200 = N134 & addr_r[6];
  assign N201 = N136 & N158;
  assign N202 = N136 & addr_r[6];
  assign N203 = N138 & N158;
  assign N204 = N138 & addr_r[6];
  assign N205 = N140 & N158;
  assign N206 = N140 & addr_r[6];
  assign N207 = N142 & N158;
  assign N208 = N142 & addr_r[6];
  assign N209 = N144 & N158;
  assign N210 = N144 & addr_r[6];
  assign N211 = N146 & N158;
  assign N212 = N146 & addr_r[6];
  assign N213 = N148 & N158;
  assign N214 = N148 & addr_r[6];
  assign N215 = N150 & N158;
  assign N216 = N150 & addr_r[6];
  assign N217 = N152 & N158;
  assign N218 = N152 & addr_r[6];
  assign N219 = N154 & N158;
  assign N220 = N154 & addr_r[6];
  assign N221 = N156 & N158;
  assign N222 = N156 & addr_r[6];
  assign N223 = N95 & N158;
  assign N224 = N95 & addr_r[6];
  assign N225 = N97 & N158;
  assign N226 = N97 & addr_r[6];
  assign N227 = N99 & N158;
  assign N228 = N99 & addr_r[6];
  assign N229 = N101 & N158;
  assign N230 = N101 & addr_r[6];
  assign N231 = N103 & N158;
  assign N232 = N103 & addr_r[6];
  assign N233 = N105 & N158;
  assign N234 = N105 & addr_r[6];
  assign N235 = N107 & N158;
  assign N236 = N107 & addr_r[6];
  assign N237 = N109 & N158;
  assign N238 = N109 & addr_r[6];
  assign N239 = N111 & N158;
  assign N240 = N111 & addr_r[6];
  assign N241 = N113 & N158;
  assign N242 = N113 & addr_r[6];
  assign N243 = N115 & N158;
  assign N244 = N115 & addr_r[6];
  assign N245 = N117 & N158;
  assign N246 = N117 & addr_r[6];
  assign N247 = N119 & N158;
  assign N248 = N119 & addr_r[6];
  assign N249 = N121 & N158;
  assign N250 = N121 & addr_r[6];
  assign N251 = N123 & N158;
  assign N252 = N123 & addr_r[6];
  assign N253 = N125 & N158;
  assign N254 = N125 & addr_r[6];
  assign N255 = N127 & N158;
  assign N256 = N127 & addr_r[6];
  assign N257 = N129 & N158;
  assign N258 = N129 & addr_r[6];
  assign N259 = N131 & N158;
  assign N260 = N131 & addr_r[6];
  assign N261 = N133 & N158;
  assign N262 = N133 & addr_r[6];
  assign N263 = N135 & N158;
  assign N264 = N135 & addr_r[6];
  assign N265 = N137 & N158;
  assign N266 = N137 & addr_r[6];
  assign N267 = N139 & N158;
  assign N268 = N139 & addr_r[6];
  assign N269 = N141 & N158;
  assign N270 = N141 & addr_r[6];
  assign N271 = N143 & N158;
  assign N272 = N143 & addr_r[6];
  assign N273 = N145 & N158;
  assign N274 = N145 & addr_r[6];
  assign N275 = N147 & N158;
  assign N276 = N147 & addr_r[6];
  assign N277 = N149 & N158;
  assign N278 = N149 & addr_r[6];
  assign N279 = N151 & N158;
  assign N280 = N151 & addr_r[6];
  assign N281 = N153 & N158;
  assign N282 = N153 & addr_r[6];
  assign N283 = N155 & N158;
  assign N284 = N155 & addr_r[6];
  assign N285 = N157 & N158;
  assign N286 = N157 & addr_r[6];
  assign N287 = v_i & w_i;
  assign N288 = ~N287;
  assign N289 = ~w_mask_i[0];
  assign N418 = ~w_mask_i[1];
  assign N547 = ~w_mask_i[2];
  assign N724 = ~w_mask_i[3];
  assign N853 = ~w_mask_i[4];
  assign N982 = ~w_mask_i[5];
  assign N1111 = ~w_mask_i[6];
  assign N1240 = ~w_mask_i[7];
  assign N1369 = ~w_mask_i[8];
  assign N1546 = ~w_mask_i[9];
  assign N1755 = ~w_mask_i[10];
  assign N1964 = ~w_mask_i[11];
  assign N2093 = ~w_mask_i[12];
  assign N2302 = ~w_mask_i[13];
  assign N2559 = ~w_mask_i[14];

endmodule