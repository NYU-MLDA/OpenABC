module decode1_0_bf8b4530d8d246dd74ac53a13471bba17941dff7(clk, rst, stall_in, flush_in, \f_in.valid , \f_in.stop_mark , \f_in.fetch_failed , \f_in.nia , \f_in.insn , \f_in.big_endian , \f_in.next_predicted , \f_in.next_pred_ntaken , busy_out, flush_out, \f_out.redirect , \f_out.redirect_nia , \d_out.valid , \d_out.stop_mark , \d_out.nia , \d_out.insn , \d_out.ispr1 , \d_out.ispr2 , \d_out.ispro , \d_out.decode , \d_out.br_pred , \d_out.big_endian , log_out);
  wire _000_;
  wire [164:0] _001_;
  wire _002_;
  wire [46:0] _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire [164:0] _009_;
  wire [46:0] _010_;
  wire [164:0] _011_;
  wire _012_;
  wire [163:0] _013_;
  wire [46:0] _014_;
  wire [46:0] _015_;
  wire _016_;
  wire [163:0] _017_;
  wire _018_;
  wire [163:0] _019_;
  wire [46:0] _020_;
  wire [46:0] _021_;
  wire [164:0] _022_;
  wire [164:0] _023_;
  wire [46:0] _024_;
  wire [46:0] _025_;
  wire [86:0] _026_;
  reg [164:0] _027_;
  reg [164:0] _028_;
  reg [46:0] _029_;
  reg [46:0] _030_;
  reg [86:0] _031_;
  wire [5:0] _032_;
  wire [10:0] _033_;
  wire _034_;
  wire [5:0] _035_;
  wire _036_;
  wire [9:0] _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire [6:0] _055_;
  wire [4:0] _056_;
  wire [4:0] _057_;
  wire [6:0] _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire [6:0] _076_;
  wire [4:0] _077_;
  wire [4:0] _078_;
  wire [6:0] _079_;
  wire [9:0] _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire [1:0] _090_;
  wire _091_;
  wire [1:0] _092_;
  wire [1:0] _093_;
  wire [1:0] _094_;
  wire [1:0] _095_;
  wire [9:0] _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire [6:0] _105_;
  wire [6:0] _106_;
  wire [6:0] _107_;
  wire _108_;
  wire [6:0] _109_;
  wire _110_;
  wire [9:0] _111_;
  wire _112_;
  wire [2:0] _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire [6:0] _119_;
  wire [6:0] _120_;
  wire [6:0] _121_;
  wire _122_;
  wire _123_;
  wire [6:0] _124_;
  wire [6:0] _125_;
  wire [13:0] _126_;
  wire [6:0] _127_;
  wire _128_;
  wire [31:0] _129_;
  wire _130_;
  wire [44:0] _131_;
  wire _132_;
  wire [3:0] _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire [1:0] _138_;
  wire _139_;
  wire [4:0] _140_;
  wire _141_;
  wire [9:0] _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire [1:0] _148_;
  wire _149_;
  wire _150_;
  wire [8:0] _151_;
  wire [4:0] _152_;
  wire [43:0] _153_;
  wire _154_;
  wire [6:0] _155_;
  wire [6:0] _156_;
  wire [6:0] _157_;
  wire [43:0] _158_;
  wire _159_;
  wire _160_;
  wire [1:0] _161_;
  wire [41:0] _162_;
  wire [1:0] _163_;
  wire [23:0] _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire [44:0] _169_;
  wire [61:0] _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire [61:0] _180_;
  wire [1:0] _181_;
  wire [1:0] _182_;
  wire _183_;
  wire _184_;
  wire [1:0] _185_;
  wire [38:0] _186_;
  wire _187_;
  wire [2815:0] _188_;
  wire [43:0] _189_;
  wire [2047:0] _190_;
  wire _191_;
  wire [2815:0] _192_;
  wire [43:0] _193_;
  wire [45055:0] _194_;
  wire [43:0] _195_;
  wire [1023:0] _196_;
  wire _197_;
  wire [351:0] _198_;
  wire [43:0] _199_;
  wire [703:0] _200_;
  wire [43:0] _201_;
  wire [175:0] _202_;
  wire [43:0] _203_;
  wire [1407:0] _204_;
  wire [43:0] _205_;
  wire [175:0] _206_;
  wire [43:0] _207_;
  wire [22527:0] _208_;
  wire [43:0] _209_;
  wire [747:0] _210_;
  wire [43:0] _211_;
  wire [86:0] br;
  wire [86:0] br_in;
  output busy_out;
  wire busy_out;
  input clk;
  wire clk;
  output \d_out.big_endian ;
  wire \d_out.big_endian ;
  output \d_out.br_pred ;
  wire \d_out.br_pred ;
  output [43:0] \d_out.decode ;
  wire [43:0] \d_out.decode ;
  output [31:0] \d_out.insn ;
  wire [31:0] \d_out.insn ;
  output [6:0] \d_out.ispr1 ;
  wire [6:0] \d_out.ispr1 ;
  output [6:0] \d_out.ispr2 ;
  wire [6:0] \d_out.ispr2 ;
  output [6:0] \d_out.ispro ;
  wire [6:0] \d_out.ispro ;
  output [63:0] \d_out.nia ;
  wire [63:0] \d_out.nia ;
  output \d_out.stop_mark ;
  wire \d_out.stop_mark ;
  output \d_out.valid ;
  wire \d_out.valid ;
  input \f_in.big_endian ;
  wire \f_in.big_endian ;
  input \f_in.fetch_failed ;
  wire \f_in.fetch_failed ;
  input [31:0] \f_in.insn ;
  wire [31:0] \f_in.insn ;
  input \f_in.next_pred_ntaken ;
  wire \f_in.next_pred_ntaken ;
  input \f_in.next_predicted ;
  wire \f_in.next_predicted ;
  input [63:0] \f_in.nia ;
  wire [63:0] \f_in.nia ;
  input \f_in.stop_mark ;
  wire \f_in.stop_mark ;
  input \f_in.valid ;
  wire \f_in.valid ;
  output \f_out.redirect ;
  wire \f_out.redirect ;
  output [63:0] \f_out.redirect_nia ;
  wire [63:0] \f_out.redirect_nia ;
  input flush_in;
  wire flush_in;
  output flush_out;
  wire flush_out;
  output [12:0] log_out;
  wire [12:0] log_out;
  wire [164:0] r;
  wire [46:0] ri;
  wire [46:0] ri_in;
  wire [164:0] rin;
  input rst;
  wire rst;
  wire [164:0] s;
  wire [46:0] si;
  input stall_in;
  wire stall_in;
  reg [43:0] \8046  [63:0];
  initial begin
    \8046 [0] = 44'h00000000000;
    \8046 [1] = 44'h00000000000;
    \8046 [2] = 44'h00000000000;
    \8046 [3] = 44'h00000000000;
    \8046 [4] = 44'h00000000000;
    \8046 [5] = 44'h00000000000;
    \8046 [6] = 44'h00000000000;
    \8046 [7] = 44'h8008008a4fa;
    \8046 [8] = 44'h00480143506;
    \8046 [9] = 44'h00080043506;
    \8046 [10] = 44'h01460143506;
    \8046 [11] = 44'h01060043506;
    \8046 [12] = 44'hc04802034fe;
    \8046 [13] = 44'h000802034fe;
    \8046 [14] = 44'hc14602034fe;
    \8046 [15] = 44'h010602034fe;
    \8046 [16] = 44'h00000000000;
    \8046 [17] = 44'h00000000000;
    \8046 [18] = 44'h00440113502;
    \8046 [19] = 44'h00040013502;
    \8046 [20] = 44'hc06400834fa;
    \8046 [21] = 44'h002400834fa;
    \8046 [22] = 44'hc04400834fa;
    \8046 [23] = 44'h000400834fa;
    \8046 [24] = 44'h00420113502;
    \8046 [25] = 44'h00020013502;
    \8046 [26] = 44'h00460113502;
    \8046 [27] = 44'h00060013502;
    \8046 [28] = 44'hc04200834fa;
    \8046 [29] = 44'h000200834fa;
    \8046 [30] = 44'hc04600834fa;
    \8046 [31] = 44'h000600834fa;
    \8046 [32] = 44'h00000000000;
    \8046 [33] = 44'h00000000000;
    \8046 [34] = 44'h04000115019;
    \8046 [35] = 44'h04000112019;
    \8046 [36] = 44'h000001151d1;
    \8046 [37] = 44'h000001121d1;
    \8046 [38] = 44'h00000115161;
    \8046 [39] = 44'h00000112161;
    \8046 [40] = 44'h09000111181;
    \8046 [41] = 44'h00000000000;
    \8046 [42] = 44'h0900011d181;
    \8046 [43] = 44'h0900011d381;
    \8046 [44] = 44'h00000000000;
    \8046 [45] = 44'h10000186029;
    \8046 [46] = 44'h00000000199;
    \8046 [47] = 44'h10000587631;
    \8046 [48] = 44'h00000084411;
    \8046 [49] = 44'h00000083411;
    \8046 [50] = 44'h04010083211;
    \8046 [51] = 44'h00010083211;
    \8046 [52] = 44'h0200d803249;
    \8046 [53] = 44'h0000d802249;
    \8046 [54] = 44'h00000000000;
    \8046 [55] = 44'h0001d083211;
    \8046 [56] = 44'h02000083349;
    \8046 [57] = 44'h00000000000;
    \8046 [58] = 44'h00000000000;
    \8046 [59] = 44'h00000000000;
    \8046 [60] = 44'h010000033c9;
    \8046 [61] = 44'h000000033c9;
    \8046 [62] = 44'h00000000000;
    \8046 [63] = 44'h20000000021;
  end
  assign _189_ = \8046 [_032_];
  reg [0:0] \8048  [2047:0];
  initial begin
    \8048 [0] = 1'h0;
    \8048 [1] = 1'h0;
    \8048 [2] = 1'h0;
    \8048 [3] = 1'h0;
    \8048 [4] = 1'h0;
    \8048 [5] = 1'h0;
    \8048 [6] = 1'h0;
    \8048 [7] = 1'h0;
    \8048 [8] = 1'h0;
    \8048 [9] = 1'h0;
    \8048 [10] = 1'h0;
    \8048 [11] = 1'h0;
    \8048 [12] = 1'h0;
    \8048 [13] = 1'h0;
    \8048 [14] = 1'h0;
    \8048 [15] = 1'h0;
    \8048 [16] = 1'h0;
    \8048 [17] = 1'h0;
    \8048 [18] = 1'h0;
    \8048 [19] = 1'h0;
    \8048 [20] = 1'h0;
    \8048 [21] = 1'h0;
    \8048 [22] = 1'h0;
    \8048 [23] = 1'h0;
    \8048 [24] = 1'h0;
    \8048 [25] = 1'h0;
    \8048 [26] = 1'h0;
    \8048 [27] = 1'h0;
    \8048 [28] = 1'h0;
    \8048 [29] = 1'h0;
    \8048 [30] = 1'h0;
    \8048 [31] = 1'h0;
    \8048 [32] = 1'h0;
    \8048 [33] = 1'h0;
    \8048 [34] = 1'h0;
    \8048 [35] = 1'h0;
    \8048 [36] = 1'h0;
    \8048 [37] = 1'h0;
    \8048 [38] = 1'h0;
    \8048 [39] = 1'h0;
    \8048 [40] = 1'h0;
    \8048 [41] = 1'h0;
    \8048 [42] = 1'h0;
    \8048 [43] = 1'h0;
    \8048 [44] = 1'h0;
    \8048 [45] = 1'h0;
    \8048 [46] = 1'h0;
    \8048 [47] = 1'h0;
    \8048 [48] = 1'h0;
    \8048 [49] = 1'h0;
    \8048 [50] = 1'h0;
    \8048 [51] = 1'h0;
    \8048 [52] = 1'h0;
    \8048 [53] = 1'h0;
    \8048 [54] = 1'h0;
    \8048 [55] = 1'h0;
    \8048 [56] = 1'h0;
    \8048 [57] = 1'h0;
    \8048 [58] = 1'h0;
    \8048 [59] = 1'h0;
    \8048 [60] = 1'h0;
    \8048 [61] = 1'h0;
    \8048 [62] = 1'h0;
    \8048 [63] = 1'h0;
    \8048 [64] = 1'h0;
    \8048 [65] = 1'h0;
    \8048 [66] = 1'h0;
    \8048 [67] = 1'h0;
    \8048 [68] = 1'h0;
    \8048 [69] = 1'h0;
    \8048 [70] = 1'h0;
    \8048 [71] = 1'h0;
    \8048 [72] = 1'h0;
    \8048 [73] = 1'h0;
    \8048 [74] = 1'h0;
    \8048 [75] = 1'h0;
    \8048 [76] = 1'h0;
    \8048 [77] = 1'h0;
    \8048 [78] = 1'h0;
    \8048 [79] = 1'h0;
    \8048 [80] = 1'h0;
    \8048 [81] = 1'h0;
    \8048 [82] = 1'h0;
    \8048 [83] = 1'h0;
    \8048 [84] = 1'h0;
    \8048 [85] = 1'h0;
    \8048 [86] = 1'h0;
    \8048 [87] = 1'h0;
    \8048 [88] = 1'h0;
    \8048 [89] = 1'h0;
    \8048 [90] = 1'h0;
    \8048 [91] = 1'h0;
    \8048 [92] = 1'h0;
    \8048 [93] = 1'h0;
    \8048 [94] = 1'h0;
    \8048 [95] = 1'h0;
    \8048 [96] = 1'h0;
    \8048 [97] = 1'h0;
    \8048 [98] = 1'h0;
    \8048 [99] = 1'h0;
    \8048 [100] = 1'h0;
    \8048 [101] = 1'h0;
    \8048 [102] = 1'h0;
    \8048 [103] = 1'h0;
    \8048 [104] = 1'h0;
    \8048 [105] = 1'h0;
    \8048 [106] = 1'h0;
    \8048 [107] = 1'h0;
    \8048 [108] = 1'h0;
    \8048 [109] = 1'h0;
    \8048 [110] = 1'h0;
    \8048 [111] = 1'h0;
    \8048 [112] = 1'h0;
    \8048 [113] = 1'h0;
    \8048 [114] = 1'h0;
    \8048 [115] = 1'h0;
    \8048 [116] = 1'h0;
    \8048 [117] = 1'h0;
    \8048 [118] = 1'h0;
    \8048 [119] = 1'h0;
    \8048 [120] = 1'h0;
    \8048 [121] = 1'h0;
    \8048 [122] = 1'h0;
    \8048 [123] = 1'h0;
    \8048 [124] = 1'h0;
    \8048 [125] = 1'h0;
    \8048 [126] = 1'h0;
    \8048 [127] = 1'h0;
    \8048 [128] = 1'h0;
    \8048 [129] = 1'h0;
    \8048 [130] = 1'h0;
    \8048 [131] = 1'h0;
    \8048 [132] = 1'h0;
    \8048 [133] = 1'h0;
    \8048 [134] = 1'h0;
    \8048 [135] = 1'h0;
    \8048 [136] = 1'h0;
    \8048 [137] = 1'h0;
    \8048 [138] = 1'h0;
    \8048 [139] = 1'h0;
    \8048 [140] = 1'h0;
    \8048 [141] = 1'h0;
    \8048 [142] = 1'h0;
    \8048 [143] = 1'h0;
    \8048 [144] = 1'h0;
    \8048 [145] = 1'h0;
    \8048 [146] = 1'h0;
    \8048 [147] = 1'h0;
    \8048 [148] = 1'h0;
    \8048 [149] = 1'h0;
    \8048 [150] = 1'h0;
    \8048 [151] = 1'h0;
    \8048 [152] = 1'h0;
    \8048 [153] = 1'h0;
    \8048 [154] = 1'h0;
    \8048 [155] = 1'h0;
    \8048 [156] = 1'h0;
    \8048 [157] = 1'h0;
    \8048 [158] = 1'h0;
    \8048 [159] = 1'h0;
    \8048 [160] = 1'h0;
    \8048 [161] = 1'h0;
    \8048 [162] = 1'h0;
    \8048 [163] = 1'h0;
    \8048 [164] = 1'h0;
    \8048 [165] = 1'h0;
    \8048 [166] = 1'h0;
    \8048 [167] = 1'h0;
    \8048 [168] = 1'h0;
    \8048 [169] = 1'h0;
    \8048 [170] = 1'h0;
    \8048 [171] = 1'h0;
    \8048 [172] = 1'h0;
    \8048 [173] = 1'h0;
    \8048 [174] = 1'h0;
    \8048 [175] = 1'h0;
    \8048 [176] = 1'h0;
    \8048 [177] = 1'h0;
    \8048 [178] = 1'h0;
    \8048 [179] = 1'h0;
    \8048 [180] = 1'h0;
    \8048 [181] = 1'h0;
    \8048 [182] = 1'h0;
    \8048 [183] = 1'h0;
    \8048 [184] = 1'h0;
    \8048 [185] = 1'h0;
    \8048 [186] = 1'h0;
    \8048 [187] = 1'h0;
    \8048 [188] = 1'h0;
    \8048 [189] = 1'h0;
    \8048 [190] = 1'h0;
    \8048 [191] = 1'h0;
    \8048 [192] = 1'h0;
    \8048 [193] = 1'h0;
    \8048 [194] = 1'h0;
    \8048 [195] = 1'h0;
    \8048 [196] = 1'h0;
    \8048 [197] = 1'h0;
    \8048 [198] = 1'h0;
    \8048 [199] = 1'h0;
    \8048 [200] = 1'h0;
    \8048 [201] = 1'h0;
    \8048 [202] = 1'h0;
    \8048 [203] = 1'h0;
    \8048 [204] = 1'h0;
    \8048 [205] = 1'h0;
    \8048 [206] = 1'h0;
    \8048 [207] = 1'h0;
    \8048 [208] = 1'h0;
    \8048 [209] = 1'h0;
    \8048 [210] = 1'h0;
    \8048 [211] = 1'h0;
    \8048 [212] = 1'h0;
    \8048 [213] = 1'h0;
    \8048 [214] = 1'h0;
    \8048 [215] = 1'h0;
    \8048 [216] = 1'h0;
    \8048 [217] = 1'h0;
    \8048 [218] = 1'h0;
    \8048 [219] = 1'h0;
    \8048 [220] = 1'h0;
    \8048 [221] = 1'h0;
    \8048 [222] = 1'h0;
    \8048 [223] = 1'h0;
    \8048 [224] = 1'h0;
    \8048 [225] = 1'h0;
    \8048 [226] = 1'h0;
    \8048 [227] = 1'h0;
    \8048 [228] = 1'h0;
    \8048 [229] = 1'h0;
    \8048 [230] = 1'h0;
    \8048 [231] = 1'h0;
    \8048 [232] = 1'h0;
    \8048 [233] = 1'h0;
    \8048 [234] = 1'h0;
    \8048 [235] = 1'h0;
    \8048 [236] = 1'h0;
    \8048 [237] = 1'h0;
    \8048 [238] = 1'h0;
    \8048 [239] = 1'h0;
    \8048 [240] = 1'h0;
    \8048 [241] = 1'h0;
    \8048 [242] = 1'h0;
    \8048 [243] = 1'h0;
    \8048 [244] = 1'h0;
    \8048 [245] = 1'h0;
    \8048 [246] = 1'h0;
    \8048 [247] = 1'h0;
    \8048 [248] = 1'h0;
    \8048 [249] = 1'h0;
    \8048 [250] = 1'h0;
    \8048 [251] = 1'h0;
    \8048 [252] = 1'h0;
    \8048 [253] = 1'h0;
    \8048 [254] = 1'h0;
    \8048 [255] = 1'h0;
    \8048 [256] = 1'h0;
    \8048 [257] = 1'h0;
    \8048 [258] = 1'h0;
    \8048 [259] = 1'h0;
    \8048 [260] = 1'h0;
    \8048 [261] = 1'h0;
    \8048 [262] = 1'h0;
    \8048 [263] = 1'h0;
    \8048 [264] = 1'h0;
    \8048 [265] = 1'h0;
    \8048 [266] = 1'h0;
    \8048 [267] = 1'h0;
    \8048 [268] = 1'h0;
    \8048 [269] = 1'h0;
    \8048 [270] = 1'h0;
    \8048 [271] = 1'h0;
    \8048 [272] = 1'h0;
    \8048 [273] = 1'h0;
    \8048 [274] = 1'h0;
    \8048 [275] = 1'h0;
    \8048 [276] = 1'h0;
    \8048 [277] = 1'h0;
    \8048 [278] = 1'h0;
    \8048 [279] = 1'h0;
    \8048 [280] = 1'h0;
    \8048 [281] = 1'h0;
    \8048 [282] = 1'h0;
    \8048 [283] = 1'h0;
    \8048 [284] = 1'h0;
    \8048 [285] = 1'h0;
    \8048 [286] = 1'h0;
    \8048 [287] = 1'h0;
    \8048 [288] = 1'h0;
    \8048 [289] = 1'h0;
    \8048 [290] = 1'h0;
    \8048 [291] = 1'h0;
    \8048 [292] = 1'h0;
    \8048 [293] = 1'h0;
    \8048 [294] = 1'h0;
    \8048 [295] = 1'h0;
    \8048 [296] = 1'h0;
    \8048 [297] = 1'h0;
    \8048 [298] = 1'h0;
    \8048 [299] = 1'h0;
    \8048 [300] = 1'h0;
    \8048 [301] = 1'h0;
    \8048 [302] = 1'h0;
    \8048 [303] = 1'h0;
    \8048 [304] = 1'h0;
    \8048 [305] = 1'h0;
    \8048 [306] = 1'h0;
    \8048 [307] = 1'h0;
    \8048 [308] = 1'h0;
    \8048 [309] = 1'h0;
    \8048 [310] = 1'h0;
    \8048 [311] = 1'h0;
    \8048 [312] = 1'h0;
    \8048 [313] = 1'h0;
    \8048 [314] = 1'h0;
    \8048 [315] = 1'h0;
    \8048 [316] = 1'h0;
    \8048 [317] = 1'h0;
    \8048 [318] = 1'h0;
    \8048 [319] = 1'h0;
    \8048 [320] = 1'h0;
    \8048 [321] = 1'h0;
    \8048 [322] = 1'h0;
    \8048 [323] = 1'h0;
    \8048 [324] = 1'h0;
    \8048 [325] = 1'h0;
    \8048 [326] = 1'h0;
    \8048 [327] = 1'h0;
    \8048 [328] = 1'h0;
    \8048 [329] = 1'h0;
    \8048 [330] = 1'h0;
    \8048 [331] = 1'h0;
    \8048 [332] = 1'h0;
    \8048 [333] = 1'h0;
    \8048 [334] = 1'h0;
    \8048 [335] = 1'h0;
    \8048 [336] = 1'h0;
    \8048 [337] = 1'h0;
    \8048 [338] = 1'h0;
    \8048 [339] = 1'h0;
    \8048 [340] = 1'h0;
    \8048 [341] = 1'h0;
    \8048 [342] = 1'h0;
    \8048 [343] = 1'h0;
    \8048 [344] = 1'h0;
    \8048 [345] = 1'h0;
    \8048 [346] = 1'h0;
    \8048 [347] = 1'h0;
    \8048 [348] = 1'h0;
    \8048 [349] = 1'h0;
    \8048 [350] = 1'h0;
    \8048 [351] = 1'h0;
    \8048 [352] = 1'h0;
    \8048 [353] = 1'h0;
    \8048 [354] = 1'h0;
    \8048 [355] = 1'h0;
    \8048 [356] = 1'h0;
    \8048 [357] = 1'h0;
    \8048 [358] = 1'h0;
    \8048 [359] = 1'h0;
    \8048 [360] = 1'h0;
    \8048 [361] = 1'h0;
    \8048 [362] = 1'h0;
    \8048 [363] = 1'h0;
    \8048 [364] = 1'h0;
    \8048 [365] = 1'h0;
    \8048 [366] = 1'h0;
    \8048 [367] = 1'h0;
    \8048 [368] = 1'h0;
    \8048 [369] = 1'h0;
    \8048 [370] = 1'h0;
    \8048 [371] = 1'h0;
    \8048 [372] = 1'h0;
    \8048 [373] = 1'h0;
    \8048 [374] = 1'h0;
    \8048 [375] = 1'h0;
    \8048 [376] = 1'h0;
    \8048 [377] = 1'h0;
    \8048 [378] = 1'h0;
    \8048 [379] = 1'h0;
    \8048 [380] = 1'h0;
    \8048 [381] = 1'h0;
    \8048 [382] = 1'h0;
    \8048 [383] = 1'h0;
    \8048 [384] = 1'h1;
    \8048 [385] = 1'h1;
    \8048 [386] = 1'h1;
    \8048 [387] = 1'h1;
    \8048 [388] = 1'h1;
    \8048 [389] = 1'h1;
    \8048 [390] = 1'h1;
    \8048 [391] = 1'h1;
    \8048 [392] = 1'h1;
    \8048 [393] = 1'h1;
    \8048 [394] = 1'h1;
    \8048 [395] = 1'h1;
    \8048 [396] = 1'h1;
    \8048 [397] = 1'h1;
    \8048 [398] = 1'h1;
    \8048 [399] = 1'h1;
    \8048 [400] = 1'h1;
    \8048 [401] = 1'h1;
    \8048 [402] = 1'h1;
    \8048 [403] = 1'h1;
    \8048 [404] = 1'h1;
    \8048 [405] = 1'h1;
    \8048 [406] = 1'h1;
    \8048 [407] = 1'h1;
    \8048 [408] = 1'h1;
    \8048 [409] = 1'h1;
    \8048 [410] = 1'h1;
    \8048 [411] = 1'h1;
    \8048 [412] = 1'h1;
    \8048 [413] = 1'h1;
    \8048 [414] = 1'h1;
    \8048 [415] = 1'h1;
    \8048 [416] = 1'h0;
    \8048 [417] = 1'h0;
    \8048 [418] = 1'h0;
    \8048 [419] = 1'h0;
    \8048 [420] = 1'h0;
    \8048 [421] = 1'h0;
    \8048 [422] = 1'h0;
    \8048 [423] = 1'h0;
    \8048 [424] = 1'h0;
    \8048 [425] = 1'h0;
    \8048 [426] = 1'h0;
    \8048 [427] = 1'h0;
    \8048 [428] = 1'h0;
    \8048 [429] = 1'h0;
    \8048 [430] = 1'h0;
    \8048 [431] = 1'h0;
    \8048 [432] = 1'h0;
    \8048 [433] = 1'h0;
    \8048 [434] = 1'h0;
    \8048 [435] = 1'h0;
    \8048 [436] = 1'h0;
    \8048 [437] = 1'h0;
    \8048 [438] = 1'h0;
    \8048 [439] = 1'h0;
    \8048 [440] = 1'h0;
    \8048 [441] = 1'h0;
    \8048 [442] = 1'h0;
    \8048 [443] = 1'h0;
    \8048 [444] = 1'h0;
    \8048 [445] = 1'h0;
    \8048 [446] = 1'h0;
    \8048 [447] = 1'h0;
    \8048 [448] = 1'h1;
    \8048 [449] = 1'h1;
    \8048 [450] = 1'h1;
    \8048 [451] = 1'h1;
    \8048 [452] = 1'h1;
    \8048 [453] = 1'h1;
    \8048 [454] = 1'h1;
    \8048 [455] = 1'h1;
    \8048 [456] = 1'h1;
    \8048 [457] = 1'h1;
    \8048 [458] = 1'h1;
    \8048 [459] = 1'h1;
    \8048 [460] = 1'h1;
    \8048 [461] = 1'h1;
    \8048 [462] = 1'h1;
    \8048 [463] = 1'h1;
    \8048 [464] = 1'h1;
    \8048 [465] = 1'h1;
    \8048 [466] = 1'h1;
    \8048 [467] = 1'h1;
    \8048 [468] = 1'h1;
    \8048 [469] = 1'h1;
    \8048 [470] = 1'h1;
    \8048 [471] = 1'h1;
    \8048 [472] = 1'h1;
    \8048 [473] = 1'h1;
    \8048 [474] = 1'h1;
    \8048 [475] = 1'h1;
    \8048 [476] = 1'h1;
    \8048 [477] = 1'h1;
    \8048 [478] = 1'h1;
    \8048 [479] = 1'h1;
    \8048 [480] = 1'h1;
    \8048 [481] = 1'h1;
    \8048 [482] = 1'h1;
    \8048 [483] = 1'h1;
    \8048 [484] = 1'h1;
    \8048 [485] = 1'h1;
    \8048 [486] = 1'h1;
    \8048 [487] = 1'h1;
    \8048 [488] = 1'h1;
    \8048 [489] = 1'h1;
    \8048 [490] = 1'h1;
    \8048 [491] = 1'h1;
    \8048 [492] = 1'h1;
    \8048 [493] = 1'h1;
    \8048 [494] = 1'h1;
    \8048 [495] = 1'h1;
    \8048 [496] = 1'h1;
    \8048 [497] = 1'h1;
    \8048 [498] = 1'h1;
    \8048 [499] = 1'h1;
    \8048 [500] = 1'h1;
    \8048 [501] = 1'h1;
    \8048 [502] = 1'h1;
    \8048 [503] = 1'h1;
    \8048 [504] = 1'h1;
    \8048 [505] = 1'h1;
    \8048 [506] = 1'h1;
    \8048 [507] = 1'h1;
    \8048 [508] = 1'h1;
    \8048 [509] = 1'h1;
    \8048 [510] = 1'h1;
    \8048 [511] = 1'h1;
    \8048 [512] = 1'h0;
    \8048 [513] = 1'h0;
    \8048 [514] = 1'h0;
    \8048 [515] = 1'h0;
    \8048 [516] = 1'h0;
    \8048 [517] = 1'h0;
    \8048 [518] = 1'h0;
    \8048 [519] = 1'h0;
    \8048 [520] = 1'h0;
    \8048 [521] = 1'h0;
    \8048 [522] = 1'h0;
    \8048 [523] = 1'h0;
    \8048 [524] = 1'h0;
    \8048 [525] = 1'h0;
    \8048 [526] = 1'h0;
    \8048 [527] = 1'h0;
    \8048 [528] = 1'h0;
    \8048 [529] = 1'h0;
    \8048 [530] = 1'h0;
    \8048 [531] = 1'h0;
    \8048 [532] = 1'h0;
    \8048 [533] = 1'h0;
    \8048 [534] = 1'h0;
    \8048 [535] = 1'h0;
    \8048 [536] = 1'h0;
    \8048 [537] = 1'h0;
    \8048 [538] = 1'h0;
    \8048 [539] = 1'h0;
    \8048 [540] = 1'h0;
    \8048 [541] = 1'h0;
    \8048 [542] = 1'h0;
    \8048 [543] = 1'h0;
    \8048 [544] = 1'h0;
    \8048 [545] = 1'h0;
    \8048 [546] = 1'h0;
    \8048 [547] = 1'h0;
    \8048 [548] = 1'h0;
    \8048 [549] = 1'h0;
    \8048 [550] = 1'h0;
    \8048 [551] = 1'h0;
    \8048 [552] = 1'h0;
    \8048 [553] = 1'h0;
    \8048 [554] = 1'h0;
    \8048 [555] = 1'h0;
    \8048 [556] = 1'h0;
    \8048 [557] = 1'h0;
    \8048 [558] = 1'h0;
    \8048 [559] = 1'h0;
    \8048 [560] = 1'h0;
    \8048 [561] = 1'h0;
    \8048 [562] = 1'h0;
    \8048 [563] = 1'h0;
    \8048 [564] = 1'h0;
    \8048 [565] = 1'h0;
    \8048 [566] = 1'h0;
    \8048 [567] = 1'h0;
    \8048 [568] = 1'h0;
    \8048 [569] = 1'h0;
    \8048 [570] = 1'h0;
    \8048 [571] = 1'h0;
    \8048 [572] = 1'h0;
    \8048 [573] = 1'h0;
    \8048 [574] = 1'h0;
    \8048 [575] = 1'h0;
    \8048 [576] = 1'h0;
    \8048 [577] = 1'h0;
    \8048 [578] = 1'h0;
    \8048 [579] = 1'h0;
    \8048 [580] = 1'h0;
    \8048 [581] = 1'h0;
    \8048 [582] = 1'h0;
    \8048 [583] = 1'h0;
    \8048 [584] = 1'h0;
    \8048 [585] = 1'h0;
    \8048 [586] = 1'h0;
    \8048 [587] = 1'h0;
    \8048 [588] = 1'h0;
    \8048 [589] = 1'h0;
    \8048 [590] = 1'h0;
    \8048 [591] = 1'h0;
    \8048 [592] = 1'h0;
    \8048 [593] = 1'h0;
    \8048 [594] = 1'h0;
    \8048 [595] = 1'h0;
    \8048 [596] = 1'h0;
    \8048 [597] = 1'h0;
    \8048 [598] = 1'h0;
    \8048 [599] = 1'h0;
    \8048 [600] = 1'h0;
    \8048 [601] = 1'h0;
    \8048 [602] = 1'h0;
    \8048 [603] = 1'h0;
    \8048 [604] = 1'h0;
    \8048 [605] = 1'h0;
    \8048 [606] = 1'h0;
    \8048 [607] = 1'h0;
    \8048 [608] = 1'h0;
    \8048 [609] = 1'h0;
    \8048 [610] = 1'h0;
    \8048 [611] = 1'h0;
    \8048 [612] = 1'h0;
    \8048 [613] = 1'h0;
    \8048 [614] = 1'h0;
    \8048 [615] = 1'h0;
    \8048 [616] = 1'h0;
    \8048 [617] = 1'h0;
    \8048 [618] = 1'h0;
    \8048 [619] = 1'h0;
    \8048 [620] = 1'h0;
    \8048 [621] = 1'h0;
    \8048 [622] = 1'h0;
    \8048 [623] = 1'h0;
    \8048 [624] = 1'h0;
    \8048 [625] = 1'h0;
    \8048 [626] = 1'h0;
    \8048 [627] = 1'h0;
    \8048 [628] = 1'h0;
    \8048 [629] = 1'h0;
    \8048 [630] = 1'h0;
    \8048 [631] = 1'h0;
    \8048 [632] = 1'h0;
    \8048 [633] = 1'h0;
    \8048 [634] = 1'h0;
    \8048 [635] = 1'h0;
    \8048 [636] = 1'h0;
    \8048 [637] = 1'h0;
    \8048 [638] = 1'h0;
    \8048 [639] = 1'h0;
    \8048 [640] = 1'h0;
    \8048 [641] = 1'h0;
    \8048 [642] = 1'h0;
    \8048 [643] = 1'h0;
    \8048 [644] = 1'h0;
    \8048 [645] = 1'h0;
    \8048 [646] = 1'h0;
    \8048 [647] = 1'h0;
    \8048 [648] = 1'h0;
    \8048 [649] = 1'h0;
    \8048 [650] = 1'h0;
    \8048 [651] = 1'h0;
    \8048 [652] = 1'h0;
    \8048 [653] = 1'h0;
    \8048 [654] = 1'h0;
    \8048 [655] = 1'h0;
    \8048 [656] = 1'h0;
    \8048 [657] = 1'h0;
    \8048 [658] = 1'h0;
    \8048 [659] = 1'h0;
    \8048 [660] = 1'h0;
    \8048 [661] = 1'h0;
    \8048 [662] = 1'h0;
    \8048 [663] = 1'h0;
    \8048 [664] = 1'h0;
    \8048 [665] = 1'h0;
    \8048 [666] = 1'h0;
    \8048 [667] = 1'h0;
    \8048 [668] = 1'h0;
    \8048 [669] = 1'h0;
    \8048 [670] = 1'h0;
    \8048 [671] = 1'h0;
    \8048 [672] = 1'h0;
    \8048 [673] = 1'h0;
    \8048 [674] = 1'h0;
    \8048 [675] = 1'h0;
    \8048 [676] = 1'h0;
    \8048 [677] = 1'h0;
    \8048 [678] = 1'h0;
    \8048 [679] = 1'h0;
    \8048 [680] = 1'h0;
    \8048 [681] = 1'h0;
    \8048 [682] = 1'h0;
    \8048 [683] = 1'h0;
    \8048 [684] = 1'h0;
    \8048 [685] = 1'h0;
    \8048 [686] = 1'h0;
    \8048 [687] = 1'h0;
    \8048 [688] = 1'h0;
    \8048 [689] = 1'h0;
    \8048 [690] = 1'h0;
    \8048 [691] = 1'h0;
    \8048 [692] = 1'h0;
    \8048 [693] = 1'h0;
    \8048 [694] = 1'h0;
    \8048 [695] = 1'h0;
    \8048 [696] = 1'h0;
    \8048 [697] = 1'h0;
    \8048 [698] = 1'h0;
    \8048 [699] = 1'h0;
    \8048 [700] = 1'h0;
    \8048 [701] = 1'h0;
    \8048 [702] = 1'h0;
    \8048 [703] = 1'h0;
    \8048 [704] = 1'h0;
    \8048 [705] = 1'h0;
    \8048 [706] = 1'h0;
    \8048 [707] = 1'h0;
    \8048 [708] = 1'h0;
    \8048 [709] = 1'h0;
    \8048 [710] = 1'h0;
    \8048 [711] = 1'h0;
    \8048 [712] = 1'h0;
    \8048 [713] = 1'h0;
    \8048 [714] = 1'h0;
    \8048 [715] = 1'h0;
    \8048 [716] = 1'h0;
    \8048 [717] = 1'h0;
    \8048 [718] = 1'h0;
    \8048 [719] = 1'h0;
    \8048 [720] = 1'h0;
    \8048 [721] = 1'h0;
    \8048 [722] = 1'h0;
    \8048 [723] = 1'h0;
    \8048 [724] = 1'h0;
    \8048 [725] = 1'h0;
    \8048 [726] = 1'h0;
    \8048 [727] = 1'h0;
    \8048 [728] = 1'h0;
    \8048 [729] = 1'h0;
    \8048 [730] = 1'h0;
    \8048 [731] = 1'h0;
    \8048 [732] = 1'h0;
    \8048 [733] = 1'h0;
    \8048 [734] = 1'h0;
    \8048 [735] = 1'h0;
    \8048 [736] = 1'h0;
    \8048 [737] = 1'h0;
    \8048 [738] = 1'h0;
    \8048 [739] = 1'h0;
    \8048 [740] = 1'h0;
    \8048 [741] = 1'h0;
    \8048 [742] = 1'h0;
    \8048 [743] = 1'h0;
    \8048 [744] = 1'h0;
    \8048 [745] = 1'h0;
    \8048 [746] = 1'h0;
    \8048 [747] = 1'h0;
    \8048 [748] = 1'h0;
    \8048 [749] = 1'h0;
    \8048 [750] = 1'h0;
    \8048 [751] = 1'h0;
    \8048 [752] = 1'h0;
    \8048 [753] = 1'h0;
    \8048 [754] = 1'h0;
    \8048 [755] = 1'h0;
    \8048 [756] = 1'h0;
    \8048 [757] = 1'h0;
    \8048 [758] = 1'h0;
    \8048 [759] = 1'h0;
    \8048 [760] = 1'h0;
    \8048 [761] = 1'h0;
    \8048 [762] = 1'h0;
    \8048 [763] = 1'h0;
    \8048 [764] = 1'h0;
    \8048 [765] = 1'h0;
    \8048 [766] = 1'h0;
    \8048 [767] = 1'h0;
    \8048 [768] = 1'h0;
    \8048 [769] = 1'h0;
    \8048 [770] = 1'h0;
    \8048 [771] = 1'h0;
    \8048 [772] = 1'h0;
    \8048 [773] = 1'h0;
    \8048 [774] = 1'h0;
    \8048 [775] = 1'h0;
    \8048 [776] = 1'h0;
    \8048 [777] = 1'h0;
    \8048 [778] = 1'h0;
    \8048 [779] = 1'h0;
    \8048 [780] = 1'h0;
    \8048 [781] = 1'h0;
    \8048 [782] = 1'h0;
    \8048 [783] = 1'h0;
    \8048 [784] = 1'h0;
    \8048 [785] = 1'h0;
    \8048 [786] = 1'h0;
    \8048 [787] = 1'h0;
    \8048 [788] = 1'h0;
    \8048 [789] = 1'h0;
    \8048 [790] = 1'h0;
    \8048 [791] = 1'h0;
    \8048 [792] = 1'h0;
    \8048 [793] = 1'h0;
    \8048 [794] = 1'h0;
    \8048 [795] = 1'h0;
    \8048 [796] = 1'h0;
    \8048 [797] = 1'h0;
    \8048 [798] = 1'h0;
    \8048 [799] = 1'h0;
    \8048 [800] = 1'h0;
    \8048 [801] = 1'h0;
    \8048 [802] = 1'h0;
    \8048 [803] = 1'h0;
    \8048 [804] = 1'h0;
    \8048 [805] = 1'h0;
    \8048 [806] = 1'h0;
    \8048 [807] = 1'h0;
    \8048 [808] = 1'h0;
    \8048 [809] = 1'h0;
    \8048 [810] = 1'h0;
    \8048 [811] = 1'h0;
    \8048 [812] = 1'h0;
    \8048 [813] = 1'h0;
    \8048 [814] = 1'h0;
    \8048 [815] = 1'h0;
    \8048 [816] = 1'h0;
    \8048 [817] = 1'h0;
    \8048 [818] = 1'h0;
    \8048 [819] = 1'h0;
    \8048 [820] = 1'h0;
    \8048 [821] = 1'h0;
    \8048 [822] = 1'h0;
    \8048 [823] = 1'h0;
    \8048 [824] = 1'h0;
    \8048 [825] = 1'h0;
    \8048 [826] = 1'h0;
    \8048 [827] = 1'h0;
    \8048 [828] = 1'h0;
    \8048 [829] = 1'h0;
    \8048 [830] = 1'h0;
    \8048 [831] = 1'h0;
    \8048 [832] = 1'h0;
    \8048 [833] = 1'h0;
    \8048 [834] = 1'h0;
    \8048 [835] = 1'h0;
    \8048 [836] = 1'h0;
    \8048 [837] = 1'h0;
    \8048 [838] = 1'h0;
    \8048 [839] = 1'h0;
    \8048 [840] = 1'h0;
    \8048 [841] = 1'h0;
    \8048 [842] = 1'h0;
    \8048 [843] = 1'h0;
    \8048 [844] = 1'h0;
    \8048 [845] = 1'h0;
    \8048 [846] = 1'h0;
    \8048 [847] = 1'h0;
    \8048 [848] = 1'h0;
    \8048 [849] = 1'h0;
    \8048 [850] = 1'h0;
    \8048 [851] = 1'h0;
    \8048 [852] = 1'h0;
    \8048 [853] = 1'h0;
    \8048 [854] = 1'h0;
    \8048 [855] = 1'h0;
    \8048 [856] = 1'h0;
    \8048 [857] = 1'h0;
    \8048 [858] = 1'h0;
    \8048 [859] = 1'h0;
    \8048 [860] = 1'h0;
    \8048 [861] = 1'h0;
    \8048 [862] = 1'h0;
    \8048 [863] = 1'h0;
    \8048 [864] = 1'h0;
    \8048 [865] = 1'h0;
    \8048 [866] = 1'h0;
    \8048 [867] = 1'h0;
    \8048 [868] = 1'h0;
    \8048 [869] = 1'h0;
    \8048 [870] = 1'h0;
    \8048 [871] = 1'h0;
    \8048 [872] = 1'h0;
    \8048 [873] = 1'h0;
    \8048 [874] = 1'h0;
    \8048 [875] = 1'h0;
    \8048 [876] = 1'h0;
    \8048 [877] = 1'h0;
    \8048 [878] = 1'h0;
    \8048 [879] = 1'h0;
    \8048 [880] = 1'h0;
    \8048 [881] = 1'h0;
    \8048 [882] = 1'h0;
    \8048 [883] = 1'h0;
    \8048 [884] = 1'h0;
    \8048 [885] = 1'h0;
    \8048 [886] = 1'h0;
    \8048 [887] = 1'h0;
    \8048 [888] = 1'h0;
    \8048 [889] = 1'h0;
    \8048 [890] = 1'h0;
    \8048 [891] = 1'h0;
    \8048 [892] = 1'h0;
    \8048 [893] = 1'h0;
    \8048 [894] = 1'h0;
    \8048 [895] = 1'h0;
    \8048 [896] = 1'h0;
    \8048 [897] = 1'h0;
    \8048 [898] = 1'h0;
    \8048 [899] = 1'h0;
    \8048 [900] = 1'h0;
    \8048 [901] = 1'h0;
    \8048 [902] = 1'h0;
    \8048 [903] = 1'h0;
    \8048 [904] = 1'h0;
    \8048 [905] = 1'h0;
    \8048 [906] = 1'h0;
    \8048 [907] = 1'h0;
    \8048 [908] = 1'h0;
    \8048 [909] = 1'h0;
    \8048 [910] = 1'h0;
    \8048 [911] = 1'h0;
    \8048 [912] = 1'h0;
    \8048 [913] = 1'h0;
    \8048 [914] = 1'h0;
    \8048 [915] = 1'h0;
    \8048 [916] = 1'h0;
    \8048 [917] = 1'h0;
    \8048 [918] = 1'h0;
    \8048 [919] = 1'h0;
    \8048 [920] = 1'h0;
    \8048 [921] = 1'h0;
    \8048 [922] = 1'h0;
    \8048 [923] = 1'h0;
    \8048 [924] = 1'h0;
    \8048 [925] = 1'h0;
    \8048 [926] = 1'h0;
    \8048 [927] = 1'h0;
    \8048 [928] = 1'h0;
    \8048 [929] = 1'h0;
    \8048 [930] = 1'h0;
    \8048 [931] = 1'h0;
    \8048 [932] = 1'h0;
    \8048 [933] = 1'h0;
    \8048 [934] = 1'h0;
    \8048 [935] = 1'h0;
    \8048 [936] = 1'h0;
    \8048 [937] = 1'h0;
    \8048 [938] = 1'h0;
    \8048 [939] = 1'h0;
    \8048 [940] = 1'h0;
    \8048 [941] = 1'h0;
    \8048 [942] = 1'h0;
    \8048 [943] = 1'h0;
    \8048 [944] = 1'h0;
    \8048 [945] = 1'h0;
    \8048 [946] = 1'h0;
    \8048 [947] = 1'h0;
    \8048 [948] = 1'h0;
    \8048 [949] = 1'h0;
    \8048 [950] = 1'h0;
    \8048 [951] = 1'h0;
    \8048 [952] = 1'h0;
    \8048 [953] = 1'h0;
    \8048 [954] = 1'h0;
    \8048 [955] = 1'h0;
    \8048 [956] = 1'h0;
    \8048 [957] = 1'h0;
    \8048 [958] = 1'h0;
    \8048 [959] = 1'h0;
    \8048 [960] = 1'h0;
    \8048 [961] = 1'h0;
    \8048 [962] = 1'h0;
    \8048 [963] = 1'h0;
    \8048 [964] = 1'h0;
    \8048 [965] = 1'h0;
    \8048 [966] = 1'h0;
    \8048 [967] = 1'h0;
    \8048 [968] = 1'h0;
    \8048 [969] = 1'h0;
    \8048 [970] = 1'h0;
    \8048 [971] = 1'h0;
    \8048 [972] = 1'h0;
    \8048 [973] = 1'h0;
    \8048 [974] = 1'h0;
    \8048 [975] = 1'h0;
    \8048 [976] = 1'h0;
    \8048 [977] = 1'h0;
    \8048 [978] = 1'h0;
    \8048 [979] = 1'h0;
    \8048 [980] = 1'h0;
    \8048 [981] = 1'h0;
    \8048 [982] = 1'h0;
    \8048 [983] = 1'h0;
    \8048 [984] = 1'h0;
    \8048 [985] = 1'h0;
    \8048 [986] = 1'h0;
    \8048 [987] = 1'h0;
    \8048 [988] = 1'h0;
    \8048 [989] = 1'h0;
    \8048 [990] = 1'h0;
    \8048 [991] = 1'h0;
    \8048 [992] = 1'h0;
    \8048 [993] = 1'h0;
    \8048 [994] = 1'h0;
    \8048 [995] = 1'h0;
    \8048 [996] = 1'h0;
    \8048 [997] = 1'h0;
    \8048 [998] = 1'h0;
    \8048 [999] = 1'h0;
    \8048 [1000] = 1'h0;
    \8048 [1001] = 1'h0;
    \8048 [1002] = 1'h0;
    \8048 [1003] = 1'h0;
    \8048 [1004] = 1'h0;
    \8048 [1005] = 1'h0;
    \8048 [1006] = 1'h0;
    \8048 [1007] = 1'h0;
    \8048 [1008] = 1'h0;
    \8048 [1009] = 1'h0;
    \8048 [1010] = 1'h0;
    \8048 [1011] = 1'h0;
    \8048 [1012] = 1'h0;
    \8048 [1013] = 1'h0;
    \8048 [1014] = 1'h0;
    \8048 [1015] = 1'h0;
    \8048 [1016] = 1'h0;
    \8048 [1017] = 1'h0;
    \8048 [1018] = 1'h0;
    \8048 [1019] = 1'h0;
    \8048 [1020] = 1'h0;
    \8048 [1021] = 1'h0;
    \8048 [1022] = 1'h0;
    \8048 [1023] = 1'h0;
    \8048 [1024] = 1'h0;
    \8048 [1025] = 1'h0;
    \8048 [1026] = 1'h0;
    \8048 [1027] = 1'h0;
    \8048 [1028] = 1'h0;
    \8048 [1029] = 1'h0;
    \8048 [1030] = 1'h0;
    \8048 [1031] = 1'h0;
    \8048 [1032] = 1'h0;
    \8048 [1033] = 1'h0;
    \8048 [1034] = 1'h0;
    \8048 [1035] = 1'h0;
    \8048 [1036] = 1'h0;
    \8048 [1037] = 1'h0;
    \8048 [1038] = 1'h0;
    \8048 [1039] = 1'h0;
    \8048 [1040] = 1'h0;
    \8048 [1041] = 1'h0;
    \8048 [1042] = 1'h0;
    \8048 [1043] = 1'h0;
    \8048 [1044] = 1'h0;
    \8048 [1045] = 1'h0;
    \8048 [1046] = 1'h0;
    \8048 [1047] = 1'h0;
    \8048 [1048] = 1'h0;
    \8048 [1049] = 1'h0;
    \8048 [1050] = 1'h0;
    \8048 [1051] = 1'h0;
    \8048 [1052] = 1'h0;
    \8048 [1053] = 1'h0;
    \8048 [1054] = 1'h0;
    \8048 [1055] = 1'h0;
    \8048 [1056] = 1'h0;
    \8048 [1057] = 1'h0;
    \8048 [1058] = 1'h0;
    \8048 [1059] = 1'h0;
    \8048 [1060] = 1'h0;
    \8048 [1061] = 1'h0;
    \8048 [1062] = 1'h0;
    \8048 [1063] = 1'h0;
    \8048 [1064] = 1'h0;
    \8048 [1065] = 1'h0;
    \8048 [1066] = 1'h0;
    \8048 [1067] = 1'h0;
    \8048 [1068] = 1'h0;
    \8048 [1069] = 1'h0;
    \8048 [1070] = 1'h0;
    \8048 [1071] = 1'h0;
    \8048 [1072] = 1'h0;
    \8048 [1073] = 1'h0;
    \8048 [1074] = 1'h0;
    \8048 [1075] = 1'h0;
    \8048 [1076] = 1'h0;
    \8048 [1077] = 1'h0;
    \8048 [1078] = 1'h0;
    \8048 [1079] = 1'h0;
    \8048 [1080] = 1'h0;
    \8048 [1081] = 1'h0;
    \8048 [1082] = 1'h0;
    \8048 [1083] = 1'h0;
    \8048 [1084] = 1'h0;
    \8048 [1085] = 1'h0;
    \8048 [1086] = 1'h0;
    \8048 [1087] = 1'h0;
    \8048 [1088] = 1'h0;
    \8048 [1089] = 1'h0;
    \8048 [1090] = 1'h0;
    \8048 [1091] = 1'h0;
    \8048 [1092] = 1'h0;
    \8048 [1093] = 1'h0;
    \8048 [1094] = 1'h0;
    \8048 [1095] = 1'h0;
    \8048 [1096] = 1'h0;
    \8048 [1097] = 1'h0;
    \8048 [1098] = 1'h0;
    \8048 [1099] = 1'h0;
    \8048 [1100] = 1'h0;
    \8048 [1101] = 1'h0;
    \8048 [1102] = 1'h0;
    \8048 [1103] = 1'h0;
    \8048 [1104] = 1'h0;
    \8048 [1105] = 1'h0;
    \8048 [1106] = 1'h0;
    \8048 [1107] = 1'h0;
    \8048 [1108] = 1'h0;
    \8048 [1109] = 1'h0;
    \8048 [1110] = 1'h0;
    \8048 [1111] = 1'h0;
    \8048 [1112] = 1'h0;
    \8048 [1113] = 1'h0;
    \8048 [1114] = 1'h0;
    \8048 [1115] = 1'h0;
    \8048 [1116] = 1'h0;
    \8048 [1117] = 1'h0;
    \8048 [1118] = 1'h0;
    \8048 [1119] = 1'h0;
    \8048 [1120] = 1'h0;
    \8048 [1121] = 1'h0;
    \8048 [1122] = 1'h0;
    \8048 [1123] = 1'h0;
    \8048 [1124] = 1'h0;
    \8048 [1125] = 1'h0;
    \8048 [1126] = 1'h0;
    \8048 [1127] = 1'h0;
    \8048 [1128] = 1'h0;
    \8048 [1129] = 1'h0;
    \8048 [1130] = 1'h0;
    \8048 [1131] = 1'h0;
    \8048 [1132] = 1'h0;
    \8048 [1133] = 1'h0;
    \8048 [1134] = 1'h0;
    \8048 [1135] = 1'h0;
    \8048 [1136] = 1'h0;
    \8048 [1137] = 1'h0;
    \8048 [1138] = 1'h0;
    \8048 [1139] = 1'h0;
    \8048 [1140] = 1'h0;
    \8048 [1141] = 1'h0;
    \8048 [1142] = 1'h0;
    \8048 [1143] = 1'h0;
    \8048 [1144] = 1'h0;
    \8048 [1145] = 1'h0;
    \8048 [1146] = 1'h0;
    \8048 [1147] = 1'h0;
    \8048 [1148] = 1'h0;
    \8048 [1149] = 1'h0;
    \8048 [1150] = 1'h0;
    \8048 [1151] = 1'h0;
    \8048 [1152] = 1'h0;
    \8048 [1153] = 1'h0;
    \8048 [1154] = 1'h0;
    \8048 [1155] = 1'h0;
    \8048 [1156] = 1'h0;
    \8048 [1157] = 1'h0;
    \8048 [1158] = 1'h0;
    \8048 [1159] = 1'h0;
    \8048 [1160] = 1'h0;
    \8048 [1161] = 1'h0;
    \8048 [1162] = 1'h0;
    \8048 [1163] = 1'h0;
    \8048 [1164] = 1'h0;
    \8048 [1165] = 1'h0;
    \8048 [1166] = 1'h0;
    \8048 [1167] = 1'h0;
    \8048 [1168] = 1'h0;
    \8048 [1169] = 1'h0;
    \8048 [1170] = 1'h0;
    \8048 [1171] = 1'h0;
    \8048 [1172] = 1'h0;
    \8048 [1173] = 1'h0;
    \8048 [1174] = 1'h0;
    \8048 [1175] = 1'h0;
    \8048 [1176] = 1'h0;
    \8048 [1177] = 1'h0;
    \8048 [1178] = 1'h0;
    \8048 [1179] = 1'h0;
    \8048 [1180] = 1'h0;
    \8048 [1181] = 1'h0;
    \8048 [1182] = 1'h0;
    \8048 [1183] = 1'h0;
    \8048 [1184] = 1'h0;
    \8048 [1185] = 1'h0;
    \8048 [1186] = 1'h0;
    \8048 [1187] = 1'h0;
    \8048 [1188] = 1'h0;
    \8048 [1189] = 1'h0;
    \8048 [1190] = 1'h0;
    \8048 [1191] = 1'h0;
    \8048 [1192] = 1'h0;
    \8048 [1193] = 1'h0;
    \8048 [1194] = 1'h0;
    \8048 [1195] = 1'h0;
    \8048 [1196] = 1'h0;
    \8048 [1197] = 1'h0;
    \8048 [1198] = 1'h0;
    \8048 [1199] = 1'h0;
    \8048 [1200] = 1'h0;
    \8048 [1201] = 1'h0;
    \8048 [1202] = 1'h0;
    \8048 [1203] = 1'h0;
    \8048 [1204] = 1'h0;
    \8048 [1205] = 1'h0;
    \8048 [1206] = 1'h0;
    \8048 [1207] = 1'h0;
    \8048 [1208] = 1'h0;
    \8048 [1209] = 1'h0;
    \8048 [1210] = 1'h0;
    \8048 [1211] = 1'h0;
    \8048 [1212] = 1'h0;
    \8048 [1213] = 1'h0;
    \8048 [1214] = 1'h0;
    \8048 [1215] = 1'h0;
    \8048 [1216] = 1'h0;
    \8048 [1217] = 1'h0;
    \8048 [1218] = 1'h0;
    \8048 [1219] = 1'h0;
    \8048 [1220] = 1'h0;
    \8048 [1221] = 1'h0;
    \8048 [1222] = 1'h0;
    \8048 [1223] = 1'h0;
    \8048 [1224] = 1'h0;
    \8048 [1225] = 1'h0;
    \8048 [1226] = 1'h0;
    \8048 [1227] = 1'h0;
    \8048 [1228] = 1'h0;
    \8048 [1229] = 1'h0;
    \8048 [1230] = 1'h0;
    \8048 [1231] = 1'h0;
    \8048 [1232] = 1'h0;
    \8048 [1233] = 1'h0;
    \8048 [1234] = 1'h0;
    \8048 [1235] = 1'h0;
    \8048 [1236] = 1'h0;
    \8048 [1237] = 1'h0;
    \8048 [1238] = 1'h0;
    \8048 [1239] = 1'h0;
    \8048 [1240] = 1'h0;
    \8048 [1241] = 1'h0;
    \8048 [1242] = 1'h0;
    \8048 [1243] = 1'h0;
    \8048 [1244] = 1'h0;
    \8048 [1245] = 1'h0;
    \8048 [1246] = 1'h0;
    \8048 [1247] = 1'h0;
    \8048 [1248] = 1'h0;
    \8048 [1249] = 1'h0;
    \8048 [1250] = 1'h0;
    \8048 [1251] = 1'h0;
    \8048 [1252] = 1'h0;
    \8048 [1253] = 1'h0;
    \8048 [1254] = 1'h0;
    \8048 [1255] = 1'h0;
    \8048 [1256] = 1'h0;
    \8048 [1257] = 1'h0;
    \8048 [1258] = 1'h0;
    \8048 [1259] = 1'h0;
    \8048 [1260] = 1'h0;
    \8048 [1261] = 1'h0;
    \8048 [1262] = 1'h0;
    \8048 [1263] = 1'h0;
    \8048 [1264] = 1'h0;
    \8048 [1265] = 1'h0;
    \8048 [1266] = 1'h0;
    \8048 [1267] = 1'h0;
    \8048 [1268] = 1'h0;
    \8048 [1269] = 1'h0;
    \8048 [1270] = 1'h0;
    \8048 [1271] = 1'h0;
    \8048 [1272] = 1'h0;
    \8048 [1273] = 1'h0;
    \8048 [1274] = 1'h0;
    \8048 [1275] = 1'h0;
    \8048 [1276] = 1'h0;
    \8048 [1277] = 1'h0;
    \8048 [1278] = 1'h0;
    \8048 [1279] = 1'h0;
    \8048 [1280] = 1'h0;
    \8048 [1281] = 1'h0;
    \8048 [1282] = 1'h0;
    \8048 [1283] = 1'h0;
    \8048 [1284] = 1'h0;
    \8048 [1285] = 1'h0;
    \8048 [1286] = 1'h0;
    \8048 [1287] = 1'h0;
    \8048 [1288] = 1'h0;
    \8048 [1289] = 1'h0;
    \8048 [1290] = 1'h0;
    \8048 [1291] = 1'h0;
    \8048 [1292] = 1'h0;
    \8048 [1293] = 1'h0;
    \8048 [1294] = 1'h0;
    \8048 [1295] = 1'h0;
    \8048 [1296] = 1'h0;
    \8048 [1297] = 1'h0;
    \8048 [1298] = 1'h0;
    \8048 [1299] = 1'h0;
    \8048 [1300] = 1'h0;
    \8048 [1301] = 1'h0;
    \8048 [1302] = 1'h0;
    \8048 [1303] = 1'h0;
    \8048 [1304] = 1'h0;
    \8048 [1305] = 1'h0;
    \8048 [1306] = 1'h0;
    \8048 [1307] = 1'h0;
    \8048 [1308] = 1'h0;
    \8048 [1309] = 1'h0;
    \8048 [1310] = 1'h0;
    \8048 [1311] = 1'h0;
    \8048 [1312] = 1'h0;
    \8048 [1313] = 1'h0;
    \8048 [1314] = 1'h0;
    \8048 [1315] = 1'h0;
    \8048 [1316] = 1'h0;
    \8048 [1317] = 1'h0;
    \8048 [1318] = 1'h0;
    \8048 [1319] = 1'h0;
    \8048 [1320] = 1'h0;
    \8048 [1321] = 1'h0;
    \8048 [1322] = 1'h0;
    \8048 [1323] = 1'h0;
    \8048 [1324] = 1'h0;
    \8048 [1325] = 1'h0;
    \8048 [1326] = 1'h0;
    \8048 [1327] = 1'h0;
    \8048 [1328] = 1'h0;
    \8048 [1329] = 1'h0;
    \8048 [1330] = 1'h0;
    \8048 [1331] = 1'h0;
    \8048 [1332] = 1'h0;
    \8048 [1333] = 1'h0;
    \8048 [1334] = 1'h0;
    \8048 [1335] = 1'h0;
    \8048 [1336] = 1'h0;
    \8048 [1337] = 1'h0;
    \8048 [1338] = 1'h0;
    \8048 [1339] = 1'h0;
    \8048 [1340] = 1'h0;
    \8048 [1341] = 1'h0;
    \8048 [1342] = 1'h0;
    \8048 [1343] = 1'h0;
    \8048 [1344] = 1'h0;
    \8048 [1345] = 1'h0;
    \8048 [1346] = 1'h0;
    \8048 [1347] = 1'h0;
    \8048 [1348] = 1'h0;
    \8048 [1349] = 1'h0;
    \8048 [1350] = 1'h0;
    \8048 [1351] = 1'h0;
    \8048 [1352] = 1'h0;
    \8048 [1353] = 1'h0;
    \8048 [1354] = 1'h0;
    \8048 [1355] = 1'h0;
    \8048 [1356] = 1'h0;
    \8048 [1357] = 1'h0;
    \8048 [1358] = 1'h0;
    \8048 [1359] = 1'h0;
    \8048 [1360] = 1'h0;
    \8048 [1361] = 1'h0;
    \8048 [1362] = 1'h0;
    \8048 [1363] = 1'h0;
    \8048 [1364] = 1'h0;
    \8048 [1365] = 1'h0;
    \8048 [1366] = 1'h0;
    \8048 [1367] = 1'h0;
    \8048 [1368] = 1'h0;
    \8048 [1369] = 1'h0;
    \8048 [1370] = 1'h0;
    \8048 [1371] = 1'h0;
    \8048 [1372] = 1'h0;
    \8048 [1373] = 1'h0;
    \8048 [1374] = 1'h0;
    \8048 [1375] = 1'h0;
    \8048 [1376] = 1'h0;
    \8048 [1377] = 1'h0;
    \8048 [1378] = 1'h0;
    \8048 [1379] = 1'h0;
    \8048 [1380] = 1'h0;
    \8048 [1381] = 1'h0;
    \8048 [1382] = 1'h0;
    \8048 [1383] = 1'h0;
    \8048 [1384] = 1'h0;
    \8048 [1385] = 1'h0;
    \8048 [1386] = 1'h0;
    \8048 [1387] = 1'h0;
    \8048 [1388] = 1'h0;
    \8048 [1389] = 1'h0;
    \8048 [1390] = 1'h0;
    \8048 [1391] = 1'h0;
    \8048 [1392] = 1'h0;
    \8048 [1393] = 1'h0;
    \8048 [1394] = 1'h0;
    \8048 [1395] = 1'h0;
    \8048 [1396] = 1'h0;
    \8048 [1397] = 1'h0;
    \8048 [1398] = 1'h0;
    \8048 [1399] = 1'h0;
    \8048 [1400] = 1'h0;
    \8048 [1401] = 1'h0;
    \8048 [1402] = 1'h0;
    \8048 [1403] = 1'h0;
    \8048 [1404] = 1'h0;
    \8048 [1405] = 1'h0;
    \8048 [1406] = 1'h0;
    \8048 [1407] = 1'h0;
    \8048 [1408] = 1'h0;
    \8048 [1409] = 1'h0;
    \8048 [1410] = 1'h0;
    \8048 [1411] = 1'h0;
    \8048 [1412] = 1'h0;
    \8048 [1413] = 1'h0;
    \8048 [1414] = 1'h0;
    \8048 [1415] = 1'h0;
    \8048 [1416] = 1'h0;
    \8048 [1417] = 1'h0;
    \8048 [1418] = 1'h0;
    \8048 [1419] = 1'h0;
    \8048 [1420] = 1'h0;
    \8048 [1421] = 1'h0;
    \8048 [1422] = 1'h0;
    \8048 [1423] = 1'h0;
    \8048 [1424] = 1'h0;
    \8048 [1425] = 1'h0;
    \8048 [1426] = 1'h0;
    \8048 [1427] = 1'h0;
    \8048 [1428] = 1'h0;
    \8048 [1429] = 1'h0;
    \8048 [1430] = 1'h0;
    \8048 [1431] = 1'h0;
    \8048 [1432] = 1'h0;
    \8048 [1433] = 1'h0;
    \8048 [1434] = 1'h0;
    \8048 [1435] = 1'h0;
    \8048 [1436] = 1'h0;
    \8048 [1437] = 1'h0;
    \8048 [1438] = 1'h0;
    \8048 [1439] = 1'h0;
    \8048 [1440] = 1'h0;
    \8048 [1441] = 1'h0;
    \8048 [1442] = 1'h0;
    \8048 [1443] = 1'h0;
    \8048 [1444] = 1'h0;
    \8048 [1445] = 1'h0;
    \8048 [1446] = 1'h0;
    \8048 [1447] = 1'h0;
    \8048 [1448] = 1'h0;
    \8048 [1449] = 1'h0;
    \8048 [1450] = 1'h0;
    \8048 [1451] = 1'h0;
    \8048 [1452] = 1'h0;
    \8048 [1453] = 1'h0;
    \8048 [1454] = 1'h0;
    \8048 [1455] = 1'h0;
    \8048 [1456] = 1'h0;
    \8048 [1457] = 1'h0;
    \8048 [1458] = 1'h0;
    \8048 [1459] = 1'h0;
    \8048 [1460] = 1'h0;
    \8048 [1461] = 1'h0;
    \8048 [1462] = 1'h0;
    \8048 [1463] = 1'h0;
    \8048 [1464] = 1'h0;
    \8048 [1465] = 1'h0;
    \8048 [1466] = 1'h0;
    \8048 [1467] = 1'h0;
    \8048 [1468] = 1'h0;
    \8048 [1469] = 1'h0;
    \8048 [1470] = 1'h0;
    \8048 [1471] = 1'h0;
    \8048 [1472] = 1'h0;
    \8048 [1473] = 1'h0;
    \8048 [1474] = 1'h0;
    \8048 [1475] = 1'h0;
    \8048 [1476] = 1'h0;
    \8048 [1477] = 1'h0;
    \8048 [1478] = 1'h0;
    \8048 [1479] = 1'h0;
    \8048 [1480] = 1'h0;
    \8048 [1481] = 1'h0;
    \8048 [1482] = 1'h0;
    \8048 [1483] = 1'h0;
    \8048 [1484] = 1'h0;
    \8048 [1485] = 1'h0;
    \8048 [1486] = 1'h0;
    \8048 [1487] = 1'h0;
    \8048 [1488] = 1'h0;
    \8048 [1489] = 1'h0;
    \8048 [1490] = 1'h0;
    \8048 [1491] = 1'h0;
    \8048 [1492] = 1'h0;
    \8048 [1493] = 1'h0;
    \8048 [1494] = 1'h0;
    \8048 [1495] = 1'h0;
    \8048 [1496] = 1'h0;
    \8048 [1497] = 1'h0;
    \8048 [1498] = 1'h0;
    \8048 [1499] = 1'h0;
    \8048 [1500] = 1'h0;
    \8048 [1501] = 1'h0;
    \8048 [1502] = 1'h0;
    \8048 [1503] = 1'h0;
    \8048 [1504] = 1'h0;
    \8048 [1505] = 1'h0;
    \8048 [1506] = 1'h0;
    \8048 [1507] = 1'h0;
    \8048 [1508] = 1'h0;
    \8048 [1509] = 1'h0;
    \8048 [1510] = 1'h0;
    \8048 [1511] = 1'h0;
    \8048 [1512] = 1'h0;
    \8048 [1513] = 1'h0;
    \8048 [1514] = 1'h0;
    \8048 [1515] = 1'h0;
    \8048 [1516] = 1'h0;
    \8048 [1517] = 1'h0;
    \8048 [1518] = 1'h0;
    \8048 [1519] = 1'h0;
    \8048 [1520] = 1'h0;
    \8048 [1521] = 1'h0;
    \8048 [1522] = 1'h0;
    \8048 [1523] = 1'h0;
    \8048 [1524] = 1'h0;
    \8048 [1525] = 1'h0;
    \8048 [1526] = 1'h0;
    \8048 [1527] = 1'h0;
    \8048 [1528] = 1'h0;
    \8048 [1529] = 1'h0;
    \8048 [1530] = 1'h0;
    \8048 [1531] = 1'h0;
    \8048 [1532] = 1'h0;
    \8048 [1533] = 1'h0;
    \8048 [1534] = 1'h0;
    \8048 [1535] = 1'h0;
    \8048 [1536] = 1'h0;
    \8048 [1537] = 1'h0;
    \8048 [1538] = 1'h0;
    \8048 [1539] = 1'h0;
    \8048 [1540] = 1'h0;
    \8048 [1541] = 1'h0;
    \8048 [1542] = 1'h0;
    \8048 [1543] = 1'h0;
    \8048 [1544] = 1'h0;
    \8048 [1545] = 1'h0;
    \8048 [1546] = 1'h0;
    \8048 [1547] = 1'h0;
    \8048 [1548] = 1'h0;
    \8048 [1549] = 1'h0;
    \8048 [1550] = 1'h0;
    \8048 [1551] = 1'h0;
    \8048 [1552] = 1'h0;
    \8048 [1553] = 1'h0;
    \8048 [1554] = 1'h0;
    \8048 [1555] = 1'h0;
    \8048 [1556] = 1'h0;
    \8048 [1557] = 1'h0;
    \8048 [1558] = 1'h0;
    \8048 [1559] = 1'h0;
    \8048 [1560] = 1'h0;
    \8048 [1561] = 1'h0;
    \8048 [1562] = 1'h0;
    \8048 [1563] = 1'h0;
    \8048 [1564] = 1'h0;
    \8048 [1565] = 1'h0;
    \8048 [1566] = 1'h0;
    \8048 [1567] = 1'h0;
    \8048 [1568] = 1'h0;
    \8048 [1569] = 1'h0;
    \8048 [1570] = 1'h0;
    \8048 [1571] = 1'h0;
    \8048 [1572] = 1'h0;
    \8048 [1573] = 1'h0;
    \8048 [1574] = 1'h0;
    \8048 [1575] = 1'h0;
    \8048 [1576] = 1'h0;
    \8048 [1577] = 1'h0;
    \8048 [1578] = 1'h0;
    \8048 [1579] = 1'h0;
    \8048 [1580] = 1'h0;
    \8048 [1581] = 1'h0;
    \8048 [1582] = 1'h0;
    \8048 [1583] = 1'h0;
    \8048 [1584] = 1'h0;
    \8048 [1585] = 1'h0;
    \8048 [1586] = 1'h0;
    \8048 [1587] = 1'h0;
    \8048 [1588] = 1'h0;
    \8048 [1589] = 1'h0;
    \8048 [1590] = 1'h0;
    \8048 [1591] = 1'h0;
    \8048 [1592] = 1'h0;
    \8048 [1593] = 1'h0;
    \8048 [1594] = 1'h0;
    \8048 [1595] = 1'h0;
    \8048 [1596] = 1'h0;
    \8048 [1597] = 1'h0;
    \8048 [1598] = 1'h0;
    \8048 [1599] = 1'h0;
    \8048 [1600] = 1'h0;
    \8048 [1601] = 1'h0;
    \8048 [1602] = 1'h0;
    \8048 [1603] = 1'h0;
    \8048 [1604] = 1'h0;
    \8048 [1605] = 1'h0;
    \8048 [1606] = 1'h0;
    \8048 [1607] = 1'h0;
    \8048 [1608] = 1'h0;
    \8048 [1609] = 1'h0;
    \8048 [1610] = 1'h0;
    \8048 [1611] = 1'h0;
    \8048 [1612] = 1'h0;
    \8048 [1613] = 1'h0;
    \8048 [1614] = 1'h0;
    \8048 [1615] = 1'h0;
    \8048 [1616] = 1'h0;
    \8048 [1617] = 1'h0;
    \8048 [1618] = 1'h0;
    \8048 [1619] = 1'h0;
    \8048 [1620] = 1'h0;
    \8048 [1621] = 1'h0;
    \8048 [1622] = 1'h0;
    \8048 [1623] = 1'h0;
    \8048 [1624] = 1'h0;
    \8048 [1625] = 1'h0;
    \8048 [1626] = 1'h0;
    \8048 [1627] = 1'h0;
    \8048 [1628] = 1'h0;
    \8048 [1629] = 1'h0;
    \8048 [1630] = 1'h0;
    \8048 [1631] = 1'h0;
    \8048 [1632] = 1'h0;
    \8048 [1633] = 1'h0;
    \8048 [1634] = 1'h0;
    \8048 [1635] = 1'h0;
    \8048 [1636] = 1'h0;
    \8048 [1637] = 1'h0;
    \8048 [1638] = 1'h0;
    \8048 [1639] = 1'h0;
    \8048 [1640] = 1'h0;
    \8048 [1641] = 1'h0;
    \8048 [1642] = 1'h0;
    \8048 [1643] = 1'h0;
    \8048 [1644] = 1'h0;
    \8048 [1645] = 1'h0;
    \8048 [1646] = 1'h0;
    \8048 [1647] = 1'h0;
    \8048 [1648] = 1'h0;
    \8048 [1649] = 1'h0;
    \8048 [1650] = 1'h0;
    \8048 [1651] = 1'h0;
    \8048 [1652] = 1'h0;
    \8048 [1653] = 1'h0;
    \8048 [1654] = 1'h0;
    \8048 [1655] = 1'h0;
    \8048 [1656] = 1'h0;
    \8048 [1657] = 1'h0;
    \8048 [1658] = 1'h0;
    \8048 [1659] = 1'h0;
    \8048 [1660] = 1'h0;
    \8048 [1661] = 1'h0;
    \8048 [1662] = 1'h0;
    \8048 [1663] = 1'h0;
    \8048 [1664] = 1'h0;
    \8048 [1665] = 1'h0;
    \8048 [1666] = 1'h0;
    \8048 [1667] = 1'h0;
    \8048 [1668] = 1'h0;
    \8048 [1669] = 1'h0;
    \8048 [1670] = 1'h0;
    \8048 [1671] = 1'h0;
    \8048 [1672] = 1'h0;
    \8048 [1673] = 1'h0;
    \8048 [1674] = 1'h0;
    \8048 [1675] = 1'h0;
    \8048 [1676] = 1'h0;
    \8048 [1677] = 1'h0;
    \8048 [1678] = 1'h0;
    \8048 [1679] = 1'h0;
    \8048 [1680] = 1'h0;
    \8048 [1681] = 1'h0;
    \8048 [1682] = 1'h0;
    \8048 [1683] = 1'h0;
    \8048 [1684] = 1'h0;
    \8048 [1685] = 1'h0;
    \8048 [1686] = 1'h0;
    \8048 [1687] = 1'h0;
    \8048 [1688] = 1'h0;
    \8048 [1689] = 1'h0;
    \8048 [1690] = 1'h0;
    \8048 [1691] = 1'h0;
    \8048 [1692] = 1'h0;
    \8048 [1693] = 1'h0;
    \8048 [1694] = 1'h0;
    \8048 [1695] = 1'h0;
    \8048 [1696] = 1'h0;
    \8048 [1697] = 1'h0;
    \8048 [1698] = 1'h0;
    \8048 [1699] = 1'h0;
    \8048 [1700] = 1'h0;
    \8048 [1701] = 1'h0;
    \8048 [1702] = 1'h0;
    \8048 [1703] = 1'h0;
    \8048 [1704] = 1'h0;
    \8048 [1705] = 1'h0;
    \8048 [1706] = 1'h0;
    \8048 [1707] = 1'h0;
    \8048 [1708] = 1'h0;
    \8048 [1709] = 1'h0;
    \8048 [1710] = 1'h0;
    \8048 [1711] = 1'h0;
    \8048 [1712] = 1'h0;
    \8048 [1713] = 1'h0;
    \8048 [1714] = 1'h0;
    \8048 [1715] = 1'h0;
    \8048 [1716] = 1'h0;
    \8048 [1717] = 1'h0;
    \8048 [1718] = 1'h0;
    \8048 [1719] = 1'h0;
    \8048 [1720] = 1'h0;
    \8048 [1721] = 1'h0;
    \8048 [1722] = 1'h0;
    \8048 [1723] = 1'h0;
    \8048 [1724] = 1'h0;
    \8048 [1725] = 1'h0;
    \8048 [1726] = 1'h0;
    \8048 [1727] = 1'h0;
    \8048 [1728] = 1'h0;
    \8048 [1729] = 1'h0;
    \8048 [1730] = 1'h0;
    \8048 [1731] = 1'h0;
    \8048 [1732] = 1'h0;
    \8048 [1733] = 1'h0;
    \8048 [1734] = 1'h0;
    \8048 [1735] = 1'h0;
    \8048 [1736] = 1'h0;
    \8048 [1737] = 1'h0;
    \8048 [1738] = 1'h0;
    \8048 [1739] = 1'h0;
    \8048 [1740] = 1'h0;
    \8048 [1741] = 1'h0;
    \8048 [1742] = 1'h0;
    \8048 [1743] = 1'h0;
    \8048 [1744] = 1'h0;
    \8048 [1745] = 1'h0;
    \8048 [1746] = 1'h0;
    \8048 [1747] = 1'h0;
    \8048 [1748] = 1'h0;
    \8048 [1749] = 1'h0;
    \8048 [1750] = 1'h0;
    \8048 [1751] = 1'h0;
    \8048 [1752] = 1'h0;
    \8048 [1753] = 1'h0;
    \8048 [1754] = 1'h0;
    \8048 [1755] = 1'h0;
    \8048 [1756] = 1'h0;
    \8048 [1757] = 1'h0;
    \8048 [1758] = 1'h0;
    \8048 [1759] = 1'h0;
    \8048 [1760] = 1'h0;
    \8048 [1761] = 1'h0;
    \8048 [1762] = 1'h0;
    \8048 [1763] = 1'h0;
    \8048 [1764] = 1'h0;
    \8048 [1765] = 1'h0;
    \8048 [1766] = 1'h0;
    \8048 [1767] = 1'h0;
    \8048 [1768] = 1'h0;
    \8048 [1769] = 1'h0;
    \8048 [1770] = 1'h0;
    \8048 [1771] = 1'h0;
    \8048 [1772] = 1'h0;
    \8048 [1773] = 1'h0;
    \8048 [1774] = 1'h0;
    \8048 [1775] = 1'h0;
    \8048 [1776] = 1'h0;
    \8048 [1777] = 1'h0;
    \8048 [1778] = 1'h0;
    \8048 [1779] = 1'h0;
    \8048 [1780] = 1'h0;
    \8048 [1781] = 1'h0;
    \8048 [1782] = 1'h0;
    \8048 [1783] = 1'h0;
    \8048 [1784] = 1'h0;
    \8048 [1785] = 1'h0;
    \8048 [1786] = 1'h0;
    \8048 [1787] = 1'h0;
    \8048 [1788] = 1'h0;
    \8048 [1789] = 1'h0;
    \8048 [1790] = 1'h0;
    \8048 [1791] = 1'h0;
    \8048 [1792] = 1'h0;
    \8048 [1793] = 1'h0;
    \8048 [1794] = 1'h0;
    \8048 [1795] = 1'h0;
    \8048 [1796] = 1'h0;
    \8048 [1797] = 1'h0;
    \8048 [1798] = 1'h0;
    \8048 [1799] = 1'h0;
    \8048 [1800] = 1'h0;
    \8048 [1801] = 1'h0;
    \8048 [1802] = 1'h0;
    \8048 [1803] = 1'h0;
    \8048 [1804] = 1'h0;
    \8048 [1805] = 1'h0;
    \8048 [1806] = 1'h0;
    \8048 [1807] = 1'h0;
    \8048 [1808] = 1'h0;
    \8048 [1809] = 1'h0;
    \8048 [1810] = 1'h0;
    \8048 [1811] = 1'h0;
    \8048 [1812] = 1'h0;
    \8048 [1813] = 1'h0;
    \8048 [1814] = 1'h0;
    \8048 [1815] = 1'h0;
    \8048 [1816] = 1'h0;
    \8048 [1817] = 1'h0;
    \8048 [1818] = 1'h0;
    \8048 [1819] = 1'h0;
    \8048 [1820] = 1'h0;
    \8048 [1821] = 1'h0;
    \8048 [1822] = 1'h0;
    \8048 [1823] = 1'h0;
    \8048 [1824] = 1'h0;
    \8048 [1825] = 1'h0;
    \8048 [1826] = 1'h0;
    \8048 [1827] = 1'h0;
    \8048 [1828] = 1'h0;
    \8048 [1829] = 1'h0;
    \8048 [1830] = 1'h0;
    \8048 [1831] = 1'h0;
    \8048 [1832] = 1'h0;
    \8048 [1833] = 1'h0;
    \8048 [1834] = 1'h0;
    \8048 [1835] = 1'h0;
    \8048 [1836] = 1'h0;
    \8048 [1837] = 1'h0;
    \8048 [1838] = 1'h0;
    \8048 [1839] = 1'h0;
    \8048 [1840] = 1'h0;
    \8048 [1841] = 1'h0;
    \8048 [1842] = 1'h0;
    \8048 [1843] = 1'h0;
    \8048 [1844] = 1'h0;
    \8048 [1845] = 1'h0;
    \8048 [1846] = 1'h0;
    \8048 [1847] = 1'h0;
    \8048 [1848] = 1'h0;
    \8048 [1849] = 1'h0;
    \8048 [1850] = 1'h0;
    \8048 [1851] = 1'h0;
    \8048 [1852] = 1'h0;
    \8048 [1853] = 1'h0;
    \8048 [1854] = 1'h0;
    \8048 [1855] = 1'h0;
    \8048 [1856] = 1'h0;
    \8048 [1857] = 1'h0;
    \8048 [1858] = 1'h0;
    \8048 [1859] = 1'h0;
    \8048 [1860] = 1'h0;
    \8048 [1861] = 1'h0;
    \8048 [1862] = 1'h0;
    \8048 [1863] = 1'h0;
    \8048 [1864] = 1'h0;
    \8048 [1865] = 1'h0;
    \8048 [1866] = 1'h0;
    \8048 [1867] = 1'h0;
    \8048 [1868] = 1'h0;
    \8048 [1869] = 1'h0;
    \8048 [1870] = 1'h0;
    \8048 [1871] = 1'h0;
    \8048 [1872] = 1'h0;
    \8048 [1873] = 1'h0;
    \8048 [1874] = 1'h0;
    \8048 [1875] = 1'h0;
    \8048 [1876] = 1'h0;
    \8048 [1877] = 1'h0;
    \8048 [1878] = 1'h0;
    \8048 [1879] = 1'h0;
    \8048 [1880] = 1'h0;
    \8048 [1881] = 1'h0;
    \8048 [1882] = 1'h0;
    \8048 [1883] = 1'h0;
    \8048 [1884] = 1'h0;
    \8048 [1885] = 1'h0;
    \8048 [1886] = 1'h0;
    \8048 [1887] = 1'h0;
    \8048 [1888] = 1'h0;
    \8048 [1889] = 1'h0;
    \8048 [1890] = 1'h0;
    \8048 [1891] = 1'h0;
    \8048 [1892] = 1'h0;
    \8048 [1893] = 1'h0;
    \8048 [1894] = 1'h0;
    \8048 [1895] = 1'h0;
    \8048 [1896] = 1'h0;
    \8048 [1897] = 1'h0;
    \8048 [1898] = 1'h0;
    \8048 [1899] = 1'h0;
    \8048 [1900] = 1'h0;
    \8048 [1901] = 1'h0;
    \8048 [1902] = 1'h0;
    \8048 [1903] = 1'h0;
    \8048 [1904] = 1'h0;
    \8048 [1905] = 1'h0;
    \8048 [1906] = 1'h0;
    \8048 [1907] = 1'h0;
    \8048 [1908] = 1'h0;
    \8048 [1909] = 1'h0;
    \8048 [1910] = 1'h0;
    \8048 [1911] = 1'h0;
    \8048 [1912] = 1'h0;
    \8048 [1913] = 1'h0;
    \8048 [1914] = 1'h0;
    \8048 [1915] = 1'h0;
    \8048 [1916] = 1'h0;
    \8048 [1917] = 1'h0;
    \8048 [1918] = 1'h0;
    \8048 [1919] = 1'h0;
    \8048 [1920] = 1'h0;
    \8048 [1921] = 1'h0;
    \8048 [1922] = 1'h0;
    \8048 [1923] = 1'h0;
    \8048 [1924] = 1'h0;
    \8048 [1925] = 1'h0;
    \8048 [1926] = 1'h0;
    \8048 [1927] = 1'h0;
    \8048 [1928] = 1'h0;
    \8048 [1929] = 1'h0;
    \8048 [1930] = 1'h0;
    \8048 [1931] = 1'h0;
    \8048 [1932] = 1'h0;
    \8048 [1933] = 1'h0;
    \8048 [1934] = 1'h0;
    \8048 [1935] = 1'h0;
    \8048 [1936] = 1'h0;
    \8048 [1937] = 1'h0;
    \8048 [1938] = 1'h0;
    \8048 [1939] = 1'h0;
    \8048 [1940] = 1'h0;
    \8048 [1941] = 1'h0;
    \8048 [1942] = 1'h0;
    \8048 [1943] = 1'h0;
    \8048 [1944] = 1'h0;
    \8048 [1945] = 1'h0;
    \8048 [1946] = 1'h0;
    \8048 [1947] = 1'h0;
    \8048 [1948] = 1'h0;
    \8048 [1949] = 1'h0;
    \8048 [1950] = 1'h0;
    \8048 [1951] = 1'h0;
    \8048 [1952] = 1'h0;
    \8048 [1953] = 1'h0;
    \8048 [1954] = 1'h0;
    \8048 [1955] = 1'h0;
    \8048 [1956] = 1'h0;
    \8048 [1957] = 1'h0;
    \8048 [1958] = 1'h0;
    \8048 [1959] = 1'h0;
    \8048 [1960] = 1'h0;
    \8048 [1961] = 1'h0;
    \8048 [1962] = 1'h0;
    \8048 [1963] = 1'h0;
    \8048 [1964] = 1'h0;
    \8048 [1965] = 1'h0;
    \8048 [1966] = 1'h0;
    \8048 [1967] = 1'h0;
    \8048 [1968] = 1'h0;
    \8048 [1969] = 1'h0;
    \8048 [1970] = 1'h0;
    \8048 [1971] = 1'h0;
    \8048 [1972] = 1'h0;
    \8048 [1973] = 1'h0;
    \8048 [1974] = 1'h0;
    \8048 [1975] = 1'h0;
    \8048 [1976] = 1'h0;
    \8048 [1977] = 1'h0;
    \8048 [1978] = 1'h0;
    \8048 [1979] = 1'h0;
    \8048 [1980] = 1'h0;
    \8048 [1981] = 1'h0;
    \8048 [1982] = 1'h0;
    \8048 [1983] = 1'h0;
    \8048 [1984] = 1'h0;
    \8048 [1985] = 1'h0;
    \8048 [1986] = 1'h0;
    \8048 [1987] = 1'h0;
    \8048 [1988] = 1'h0;
    \8048 [1989] = 1'h0;
    \8048 [1990] = 1'h0;
    \8048 [1991] = 1'h0;
    \8048 [1992] = 1'h0;
    \8048 [1993] = 1'h0;
    \8048 [1994] = 1'h0;
    \8048 [1995] = 1'h0;
    \8048 [1996] = 1'h0;
    \8048 [1997] = 1'h0;
    \8048 [1998] = 1'h0;
    \8048 [1999] = 1'h0;
    \8048 [2000] = 1'h0;
    \8048 [2001] = 1'h0;
    \8048 [2002] = 1'h0;
    \8048 [2003] = 1'h0;
    \8048 [2004] = 1'h0;
    \8048 [2005] = 1'h0;
    \8048 [2006] = 1'h0;
    \8048 [2007] = 1'h0;
    \8048 [2008] = 1'h0;
    \8048 [2009] = 1'h0;
    \8048 [2010] = 1'h0;
    \8048 [2011] = 1'h0;
    \8048 [2012] = 1'h0;
    \8048 [2013] = 1'h0;
    \8048 [2014] = 1'h0;
    \8048 [2015] = 1'h0;
    \8048 [2016] = 1'h0;
    \8048 [2017] = 1'h0;
    \8048 [2018] = 1'h0;
    \8048 [2019] = 1'h0;
    \8048 [2020] = 1'h0;
    \8048 [2021] = 1'h0;
    \8048 [2022] = 1'h0;
    \8048 [2023] = 1'h0;
    \8048 [2024] = 1'h0;
    \8048 [2025] = 1'h0;
    \8048 [2026] = 1'h0;
    \8048 [2027] = 1'h0;
    \8048 [2028] = 1'h0;
    \8048 [2029] = 1'h0;
    \8048 [2030] = 1'h0;
    \8048 [2031] = 1'h0;
    \8048 [2032] = 1'h0;
    \8048 [2033] = 1'h0;
    \8048 [2034] = 1'h0;
    \8048 [2035] = 1'h0;
    \8048 [2036] = 1'h0;
    \8048 [2037] = 1'h0;
    \8048 [2038] = 1'h0;
    \8048 [2039] = 1'h0;
    \8048 [2040] = 1'h0;
    \8048 [2041] = 1'h0;
    \8048 [2042] = 1'h0;
    \8048 [2043] = 1'h0;
    \8048 [2044] = 1'h0;
    \8048 [2045] = 1'h0;
    \8048 [2046] = 1'h0;
    \8048 [2047] = 1'h0;
  end
  assign _191_ = \8048 [_033_];
  reg [43:0] \8050  [63:0];
  initial begin
    \8050 [0] = 44'h00000000000;
    \8050 [1] = 44'h00000000000;
    \8050 [2] = 44'h00000000000;
    \8050 [3] = 44'h00000000000;
    \8050 [4] = 44'h00000000000;
    \8050 [5] = 44'h00000000000;
    \8050 [6] = 44'h00000000000;
    \8050 [7] = 44'h00000000000;
    \8050 [8] = 44'h00000000000;
    \8050 [9] = 44'h00000000000;
    \8050 [10] = 44'h00000000000;
    \8050 [11] = 44'h00000000000;
    \8050 [12] = 44'h020000a1349;
    \8050 [13] = 44'h00000000000;
    \8050 [14] = 44'h000000a1351;
    \8050 [15] = 44'h020000a1351;
    \8050 [16] = 44'h00000000000;
    \8050 [17] = 44'h00000000000;
    \8050 [18] = 44'h00000000000;
    \8050 [19] = 44'h00000000000;
    \8050 [20] = 44'h00000000000;
    \8050 [21] = 44'h00000000000;
    \8050 [22] = 44'h00000000000;
    \8050 [23] = 44'h00000000000;
    \8050 [24] = 44'h00000000000;
    \8050 [25] = 44'h00000000000;
    \8050 [26] = 44'h00000000000;
    \8050 [27] = 44'h00000000000;
    \8050 [28] = 44'h00000000000;
    \8050 [29] = 44'h00000000000;
    \8050 [30] = 44'h00000000000;
    \8050 [31] = 44'h00000000000;
    \8050 [32] = 44'h00000000000;
    \8050 [33] = 44'h00000000000;
    \8050 [34] = 44'h00000000000;
    \8050 [35] = 44'h00000000000;
    \8050 [36] = 44'h00000000000;
    \8050 [37] = 44'h00000000000;
    \8050 [38] = 44'h00000000000;
    \8050 [39] = 44'h00000000000;
    \8050 [40] = 44'h00000000000;
    \8050 [41] = 44'h00000000000;
    \8050 [42] = 44'h00000000000;
    \8050 [43] = 44'h00000000000;
    \8050 [44] = 44'h00000000000;
    \8050 [45] = 44'h00000000000;
    \8050 [46] = 44'h00000000000;
    \8050 [47] = 44'h00000000000;
    \8050 [48] = 44'h00000000000;
    \8050 [49] = 44'h00000000000;
    \8050 [50] = 44'h00000000000;
    \8050 [51] = 44'h00000000000;
    \8050 [52] = 44'h00000000000;
    \8050 [53] = 44'h00000000000;
    \8050 [54] = 44'h00000000000;
    \8050 [55] = 44'h00000000000;
    \8050 [56] = 44'h00000000000;
    \8050 [57] = 44'h00000000000;
    \8050 [58] = 44'h00000000000;
    \8050 [59] = 44'h00000000000;
    \8050 [60] = 44'h00000000000;
    \8050 [61] = 44'h00000000000;
    \8050 [62] = 44'h00000000000;
    \8050 [63] = 44'h00000000000;
  end
  assign _193_ = \8050 [_035_];
  reg [43:0] \8052  [1023:0];
  initial begin
    \8052 [0] = 44'h00000000000;
    \8052 [1] = 44'h00000000000;
    \8052 [2] = 44'h00000000000;
    \8052 [3] = 44'h00000000000;
    \8052 [4] = 44'h00000000000;
    \8052 [5] = 44'h00000000000;
    \8052 [6] = 44'h00000000000;
    \8052 [7] = 44'h00000000000;
    \8052 [8] = 44'h00000000000;
    \8052 [9] = 44'h000000014a2;
    \8052 [10] = 44'h00080011502;
    \8052 [11] = 44'h00000000000;
    \8052 [12] = 44'h00000000000;
    \8052 [13] = 44'h00000000000;
    \8052 [14] = 44'h00000000000;
    \8052 [15] = 44'h00000000000;
    \8052 [16] = 44'h000004814e9;
    \8052 [17] = 44'h00000000000;
    \8052 [18] = 44'h00000000000;
    \8052 [19] = 44'h00000000000;
    \8052 [20] = 44'h0b0000812a9;
    \8052 [21] = 44'h00000000000;
    \8052 [22] = 44'h0a0000812a9;
    \8052 [23] = 44'h00000000000;
    \8052 [24] = 44'h00000000000;
    \8052 [25] = 44'h00000000000;
    \8052 [26] = 44'h00000000000;
    \8052 [27] = 44'h00000000000;
    \8052 [28] = 44'h00000000000;
    \8052 [29] = 44'h00000000000;
    \8052 [30] = 44'h00000000000;
    \8052 [31] = 44'h00000000000;
    \8052 [32] = 44'h00000000000;
    \8052 [33] = 44'h00000000000;
    \8052 [34] = 44'h00000000000;
    \8052 [35] = 44'h00000000000;
    \8052 [36] = 44'h00000000000;
    \8052 [37] = 44'h080601100b9;
    \8052 [38] = 44'h00000000000;
    \8052 [39] = 44'h00000000000;
    \8052 [40] = 44'h00060041506;
    \8052 [41] = 44'h200000000d9;
    \8052 [42] = 44'h00020011502;
    \8052 [43] = 44'h00000000000;
    \8052 [44] = 44'h00000000000;
    \8052 [45] = 44'h00000000000;
    \8052 [46] = 44'h00000000000;
    \8052 [47] = 44'h00000000000;
    \8052 [48] = 44'h000004814e9;
    \8052 [49] = 44'h00000000000;
    \8052 [50] = 44'h00000000000;
    \8052 [51] = 44'h00000000000;
    \8052 [52] = 44'h090000812a9;
    \8052 [53] = 44'h00000000000;
    \8052 [54] = 44'h080000812a9;
    \8052 [55] = 44'h00000000000;
    \8052 [56] = 44'h00000000000;
    \8052 [57] = 44'h00000000000;
    \8052 [58] = 44'h00000000000;
    \8052 [59] = 44'h00000000000;
    \8052 [60] = 44'h00000000000;
    \8052 [61] = 44'h00000000000;
    \8052 [62] = 44'h00000000000;
    \8052 [63] = 44'h00000000000;
    \8052 [64] = 44'h00000000000;
    \8052 [65] = 44'h00000000000;
    \8052 [66] = 44'h00000000000;
    \8052 [67] = 44'h00000000000;
    \8052 [68] = 44'h00000000000;
    \8052 [69] = 44'h080201100b9;
    \8052 [70] = 44'h00000000000;
    \8052 [71] = 44'h00000000000;
    \8052 [72] = 44'h00000000000;
    \8052 [73] = 44'h00000000000;
    \8052 [74] = 44'h00040011502;
    \8052 [75] = 44'h00000000000;
    \8052 [76] = 44'h00000000000;
    \8052 [77] = 44'h00000000000;
    \8052 [78] = 44'h00000000000;
    \8052 [79] = 44'h00000000000;
    \8052 [80] = 44'h000004814e9;
    \8052 [81] = 44'h00000000000;
    \8052 [82] = 44'h00000000000;
    \8052 [83] = 44'h00000000000;
    \8052 [84] = 44'h0b0000812b1;
    \8052 [85] = 44'h00000000000;
    \8052 [86] = 44'h0a0000812b1;
    \8052 [87] = 44'h00000000000;
    \8052 [88] = 44'h00000000000;
    \8052 [89] = 44'h00000000000;
    \8052 [90] = 44'h00000000000;
    \8052 [91] = 44'h00000000000;
    \8052 [92] = 44'h00000000000;
    \8052 [93] = 44'h00000000000;
    \8052 [94] = 44'h00000000000;
    \8052 [95] = 44'h00000000000;
    \8052 [96] = 44'h00000000000;
    \8052 [97] = 44'h00000000000;
    \8052 [98] = 44'h00000000000;
    \8052 [99] = 44'h00000000000;
    \8052 [100] = 44'h00000000000;
    \8052 [101] = 44'h080401100b9;
    \8052 [102] = 44'h00000000000;
    \8052 [103] = 44'h00000000000;
    \8052 [104] = 44'h00000000000;
    \8052 [105] = 44'h00140011502;
    \8052 [106] = 44'h00060011502;
    \8052 [107] = 44'h00000000000;
    \8052 [108] = 44'h00000000000;
    \8052 [109] = 44'h00000000000;
    \8052 [110] = 44'h00000000000;
    \8052 [111] = 44'h00000000000;
    \8052 [112] = 44'h000004814e9;
    \8052 [113] = 44'h00000000000;
    \8052 [114] = 44'h00000000000;
    \8052 [115] = 44'h00000000000;
    \8052 [116] = 44'h090000812b1;
    \8052 [117] = 44'h00000000000;
    \8052 [118] = 44'h080000812b1;
    \8052 [119] = 44'h00000000000;
    \8052 [120] = 44'h00000000000;
    \8052 [121] = 44'h00000000000;
    \8052 [122] = 44'h00000000000;
    \8052 [123] = 44'h00000000000;
    \8052 [124] = 44'h00000000000;
    \8052 [125] = 44'h00000000000;
    \8052 [126] = 44'h00000000000;
    \8052 [127] = 44'h00000000000;
    \8052 [128] = 44'h00000000000;
    \8052 [129] = 44'h00000000000;
    \8052 [130] = 44'h00000000000;
    \8052 [131] = 44'h00000000000;
    \8052 [132] = 44'h0800011c0c1;
    \8052 [133] = 44'h0800011c0c1;
    \8052 [134] = 44'h00000000000;
    \8052 [135] = 44'h00000000000;
    \8052 [136] = 44'h000602014fe;
    \8052 [137] = 44'h00000000000;
    \8052 [138] = 44'h000800814fa;
    \8052 [139] = 44'h00000000000;
    \8052 [140] = 44'h00000000000;
    \8052 [141] = 44'h00000000000;
    \8052 [142] = 44'h00000000000;
    \8052 [143] = 44'h00000000000;
    \8052 [144] = 44'h000004814e9;
    \8052 [145] = 44'h00000000000;
    \8052 [146] = 44'h00000000000;
    \8052 [147] = 44'h00000000000;
    \8052 [148] = 44'h00000000000;
    \8052 [149] = 44'h00000000000;
    \8052 [150] = 44'h00000000000;
    \8052 [151] = 44'h00000000000;
    \8052 [152] = 44'h00000000000;
    \8052 [153] = 44'h00000000000;
    \8052 [154] = 44'h00000000000;
    \8052 [155] = 44'h00000000000;
    \8052 [156] = 44'h00000000000;
    \8052 [157] = 44'h00000000000;
    \8052 [158] = 44'h00000000000;
    \8052 [159] = 44'h00000000000;
    \8052 [160] = 44'h00000000000;
    \8052 [161] = 44'h00000000000;
    \8052 [162] = 44'h00000000000;
    \8052 [163] = 44'h00000000000;
    \8052 [164] = 44'h00000000000;
    \8052 [165] = 44'h00000000000;
    \8052 [166] = 44'h00000000000;
    \8052 [167] = 44'h00000000000;
    \8052 [168] = 44'h002602014fe;
    \8052 [169] = 44'h20000000009;
    \8052 [170] = 44'h000200814fa;
    \8052 [171] = 44'h00000000000;
    \8052 [172] = 44'h00000000000;
    \8052 [173] = 44'h00000000000;
    \8052 [174] = 44'h00000000000;
    \8052 [175] = 44'h00000000000;
    \8052 [176] = 44'h000004814e9;
    \8052 [177] = 44'h00000000000;
    \8052 [178] = 44'h00000000000;
    \8052 [179] = 44'h00000000000;
    \8052 [180] = 44'h00000000000;
    \8052 [181] = 44'h00000000000;
    \8052 [182] = 44'h00000000000;
    \8052 [183] = 44'h00000000000;
    \8052 [184] = 44'h00000000000;
    \8052 [185] = 44'h00000000000;
    \8052 [186] = 44'h00000000000;
    \8052 [187] = 44'h00000000000;
    \8052 [188] = 44'h00000000000;
    \8052 [189] = 44'h00000000000;
    \8052 [190] = 44'h00000000000;
    \8052 [191] = 44'h00000000000;
    \8052 [192] = 44'h00000000000;
    \8052 [193] = 44'h00000000000;
    \8052 [194] = 44'h00000000000;
    \8052 [195] = 44'h00000000000;
    \8052 [196] = 44'h0a01011c1b1;
    \8052 [197] = 44'h0a01011c1b1;
    \8052 [198] = 44'h00000000000;
    \8052 [199] = 44'h0b01011d1b1;
    \8052 [200] = 44'h00000000000;
    \8052 [201] = 44'h00000000009;
    \8052 [202] = 44'h000400814fa;
    \8052 [203] = 44'h00000000000;
    \8052 [204] = 44'h00000000000;
    \8052 [205] = 44'h00000000000;
    \8052 [206] = 44'h00000000000;
    \8052 [207] = 44'h00000000000;
    \8052 [208] = 44'h000004814e9;
    \8052 [209] = 44'h00000000000;
    \8052 [210] = 44'h00000000000;
    \8052 [211] = 44'h00000000000;
    \8052 [212] = 44'h00000000000;
    \8052 [213] = 44'h00000000000;
    \8052 [214] = 44'h00000000000;
    \8052 [215] = 44'h00000000000;
    \8052 [216] = 44'h00000000000;
    \8052 [217] = 44'h00000000000;
    \8052 [218] = 44'h00000000000;
    \8052 [219] = 44'h00000000000;
    \8052 [220] = 44'h00000000000;
    \8052 [221] = 44'h00000000000;
    \8052 [222] = 44'h00000000000;
    \8052 [223] = 44'h00000000000;
    \8052 [224] = 44'h00000000000;
    \8052 [225] = 44'h00000000000;
    \8052 [226] = 44'h00000000000;
    \8052 [227] = 44'h00000000000;
    \8052 [228] = 44'h00000000000;
    \8052 [229] = 44'h0a0101111b1;
    \8052 [230] = 44'h00000000000;
    \8052 [231] = 44'h0b0101111b1;
    \8052 [232] = 44'h00000000000;
    \8052 [233] = 44'h001400814fa;
    \8052 [234] = 44'h000600814fa;
    \8052 [235] = 44'h00000000000;
    \8052 [236] = 44'h00000000000;
    \8052 [237] = 44'h00000000000;
    \8052 [238] = 44'h00000000000;
    \8052 [239] = 44'h00000000000;
    \8052 [240] = 44'h000004814e9;
    \8052 [241] = 44'h00000000000;
    \8052 [242] = 44'h00000000000;
    \8052 [243] = 44'h00000000000;
    \8052 [244] = 44'h03000081329;
    \8052 [245] = 44'h08000081211;
    \8052 [246] = 44'h02000081329;
    \8052 [247] = 44'h00000000000;
    \8052 [248] = 44'h00000000000;
    \8052 [249] = 44'h00000000000;
    \8052 [250] = 44'h00000000000;
    \8052 [251] = 44'h00000000000;
    \8052 [252] = 44'h00000000000;
    \8052 [253] = 44'h00000000000;
    \8052 [254] = 44'h00000000000;
    \8052 [255] = 44'h00000000000;
    \8052 [256] = 44'h00000000000;
    \8052 [257] = 44'h00000000000;
    \8052 [258] = 44'h00000000000;
    \8052 [259] = 44'h00000000000;
    \8052 [260] = 44'h00000000000;
    \8052 [261] = 44'h00000000000;
    \8052 [262] = 44'h00000000000;
    \8052 [263] = 44'h00000000000;
    \8052 [264] = 44'h00480141506;
    \8052 [265] = 44'h00000000000;
    \8052 [266] = 44'h00000000000;
    \8052 [267] = 44'h00000000000;
    \8052 [268] = 44'h00000080079;
    \8052 [269] = 44'h00000000009;
    \8052 [270] = 44'h00000000000;
    \8052 [271] = 44'h00000000000;
    \8052 [272] = 44'h000004814e9;
    \8052 [273] = 44'h00000000000;
    \8052 [274] = 44'h00000000000;
    \8052 [275] = 44'h00000000000;
    \8052 [276] = 44'h0b000081349;
    \8052 [277] = 44'h0801408b211;
    \8052 [278] = 44'h0a000081349;
    \8052 [279] = 44'h0801508b211;
    \8052 [280] = 44'h00000000000;
    \8052 [281] = 44'h00000000000;
    \8052 [282] = 44'h00000000000;
    \8052 [283] = 44'h00000000000;
    \8052 [284] = 44'h00000000000;
    \8052 [285] = 44'h00000000000;
    \8052 [286] = 44'h00000000000;
    \8052 [287] = 44'h00000000000;
    \8052 [288] = 44'h00000000000;
    \8052 [289] = 44'h00000000000;
    \8052 [290] = 44'h00000000000;
    \8052 [291] = 44'h00000000000;
    \8052 [292] = 44'h00000000000;
    \8052 [293] = 44'h00000000000;
    \8052 [294] = 44'h00000000000;
    \8052 [295] = 44'h00000000000;
    \8052 [296] = 44'h00080041506;
    \8052 [297] = 44'h04840011502;
    \8052 [298] = 44'h00000000000;
    \8052 [299] = 44'h00000000000;
    \8052 [300] = 44'h00000000000;
    \8052 [301] = 44'h00000000009;
    \8052 [302] = 44'h00000000000;
    \8052 [303] = 44'h00000000000;
    \8052 [304] = 44'h000004814e9;
    \8052 [305] = 44'h00000000000;
    \8052 [306] = 44'h00000000000;
    \8052 [307] = 44'h00000000000;
    \8052 [308] = 44'h00000000000;
    \8052 [309] = 44'h08014080211;
    \8052 [310] = 44'h00000000000;
    \8052 [311] = 44'h08015080211;
    \8052 [312] = 44'h00000000000;
    \8052 [313] = 44'h00000000000;
    \8052 [314] = 44'h00000000000;
    \8052 [315] = 44'h00000000000;
    \8052 [316] = 44'h00000000000;
    \8052 [317] = 44'h00000000000;
    \8052 [318] = 44'h00000000000;
    \8052 [319] = 44'h00000000000;
    \8052 [320] = 44'h00000000000;
    \8052 [321] = 44'h00000000000;
    \8052 [322] = 44'h00000000000;
    \8052 [323] = 44'h00000000000;
    \8052 [324] = 44'h00000000000;
    \8052 [325] = 44'h00000000000;
    \8052 [326] = 44'h00000000000;
    \8052 [327] = 44'h00000000000;
    \8052 [328] = 44'h01460141506;
    \8052 [329] = 44'h04820011502;
    \8052 [330] = 44'h00000000000;
    \8052 [331] = 44'h00000000000;
    \8052 [332] = 44'h00000000000;
    \8052 [333] = 44'h00000000009;
    \8052 [334] = 44'h00000000000;
    \8052 [335] = 44'h00000000000;
    \8052 [336] = 44'h000004814e9;
    \8052 [337] = 44'h00000000000;
    \8052 [338] = 44'h00000000000;
    \8052 [339] = 44'h00000000000;
    \8052 [340] = 44'h00000000000;
    \8052 [341] = 44'h00000000000;
    \8052 [342] = 44'h00000000000;
    \8052 [343] = 44'h00000000000;
    \8052 [344] = 44'h00000000000;
    \8052 [345] = 44'h00000000000;
    \8052 [346] = 44'h00000000000;
    \8052 [347] = 44'h00000000000;
    \8052 [348] = 44'h00000000000;
    \8052 [349] = 44'h00000000000;
    \8052 [350] = 44'h00000000000;
    \8052 [351] = 44'h00000000000;
    \8052 [352] = 44'h00000000000;
    \8052 [353] = 44'h00000000000;
    \8052 [354] = 44'h00000000000;
    \8052 [355] = 44'h00000000000;
    \8052 [356] = 44'h00000000000;
    \8052 [357] = 44'h00000000000;
    \8052 [358] = 44'h00000000000;
    \8052 [359] = 44'h00000000000;
    \8052 [360] = 44'h01060041506;
    \8052 [361] = 44'h00160011502;
    \8052 [362] = 44'h00000000000;
    \8052 [363] = 44'h00180011502;
    \8052 [364] = 44'h00000000000;
    \8052 [365] = 44'h00000000009;
    \8052 [366] = 44'h00000000000;
    \8052 [367] = 44'h00000000000;
    \8052 [368] = 44'h000004814e9;
    \8052 [369] = 44'h00000000000;
    \8052 [370] = 44'h00000000000;
    \8052 [371] = 44'h00000000000;
    \8052 [372] = 44'h00000000000;
    \8052 [373] = 44'h08014081211;
    \8052 [374] = 44'h00000000000;
    \8052 [375] = 44'h08015081211;
    \8052 [376] = 44'h00000000000;
    \8052 [377] = 44'h00000000000;
    \8052 [378] = 44'h00000000000;
    \8052 [379] = 44'h00000000000;
    \8052 [380] = 44'h00000000000;
    \8052 [381] = 44'h00000000000;
    \8052 [382] = 44'h00000000000;
    \8052 [383] = 44'h00000000000;
    \8052 [384] = 44'h00000000000;
    \8052 [385] = 44'h00000000000;
    \8052 [386] = 44'h00000000000;
    \8052 [387] = 44'h00000000000;
    \8052 [388] = 44'h00000000000;
    \8052 [389] = 44'h00000000000;
    \8052 [390] = 44'h00000000000;
    \8052 [391] = 44'h00000000000;
    \8052 [392] = 44'hc04802014fe;
    \8052 [393] = 44'h00000000000;
    \8052 [394] = 44'h00000000000;
    \8052 [395] = 44'h00000000000;
    \8052 [396] = 44'h00000000000;
    \8052 [397] = 44'h00000000009;
    \8052 [398] = 44'h00000000000;
    \8052 [399] = 44'h00000000000;
    \8052 [400] = 44'h000004814e9;
    \8052 [401] = 44'h00000000000;
    \8052 [402] = 44'h00000000000;
    \8052 [403] = 44'h00000000000;
    \8052 [404] = 44'h00000000000;
    \8052 [405] = 44'h00000000000;
    \8052 [406] = 44'h00000000000;
    \8052 [407] = 44'h0800d080211;
    \8052 [408] = 44'h00000000000;
    \8052 [409] = 44'h00000000000;
    \8052 [410] = 44'h00000000000;
    \8052 [411] = 44'h00000000000;
    \8052 [412] = 44'h00000000000;
    \8052 [413] = 44'h00000000000;
    \8052 [414] = 44'h00000000000;
    \8052 [415] = 44'h00000000000;
    \8052 [416] = 44'h00000000000;
    \8052 [417] = 44'h00000000000;
    \8052 [418] = 44'h00000000000;
    \8052 [419] = 44'h00000000000;
    \8052 [420] = 44'h00000000000;
    \8052 [421] = 44'h00000000000;
    \8052 [422] = 44'h00000000000;
    \8052 [423] = 44'h00000000000;
    \8052 [424] = 44'h000802014fe;
    \8052 [425] = 44'h20000000009;
    \8052 [426] = 44'h00000000000;
    \8052 [427] = 44'h00000000000;
    \8052 [428] = 44'h00000000000;
    \8052 [429] = 44'h00000000009;
    \8052 [430] = 44'h00000000000;
    \8052 [431] = 44'h00000000000;
    \8052 [432] = 44'h000004814e9;
    \8052 [433] = 44'h00000000000;
    \8052 [434] = 44'h00000000000;
    \8052 [435] = 44'h00000000000;
    \8052 [436] = 44'h0b000081359;
    \8052 [437] = 44'h00000000000;
    \8052 [438] = 44'h0a000081351;
    \8052 [439] = 44'h00000000000;
    \8052 [440] = 44'h00000000000;
    \8052 [441] = 44'h00000000000;
    \8052 [442] = 44'h00000000000;
    \8052 [443] = 44'h00000000000;
    \8052 [444] = 44'h00000000000;
    \8052 [445] = 44'h00000000000;
    \8052 [446] = 44'h00000000000;
    \8052 [447] = 44'h00000800109;
    \8052 [448] = 44'h00000000000;
    \8052 [449] = 44'h00000000000;
    \8052 [450] = 44'h00000000000;
    \8052 [451] = 44'h00000000000;
    \8052 [452] = 44'h00000000000;
    \8052 [453] = 44'h08000110069;
    \8052 [454] = 44'h00000000000;
    \8052 [455] = 44'h00000000000;
    \8052 [456] = 44'hc14602014fe;
    \8052 [457] = 44'h20000000009;
    \8052 [458] = 44'h00000000000;
    \8052 [459] = 44'h00000000000;
    \8052 [460] = 44'h00000000000;
    \8052 [461] = 44'h00000000009;
    \8052 [462] = 44'h00000000000;
    \8052 [463] = 44'h00000000000;
    \8052 [464] = 44'h000004814e9;
    \8052 [465] = 44'h00000000000;
    \8052 [466] = 44'h00000000000;
    \8052 [467] = 44'h00000000000;
    \8052 [468] = 44'h00000000000;
    \8052 [469] = 44'h00000000000;
    \8052 [470] = 44'h00000000000;
    \8052 [471] = 44'h0800d081211;
    \8052 [472] = 44'h00000000000;
    \8052 [473] = 44'h00000000000;
    \8052 [474] = 44'h00000000000;
    \8052 [475] = 44'h00000000000;
    \8052 [476] = 44'h00000000000;
    \8052 [477] = 44'h00000000000;
    \8052 [478] = 44'h00000000000;
    \8052 [479] = 44'h00000000000;
    \8052 [480] = 44'h00000000000;
    \8052 [481] = 44'h00000000000;
    \8052 [482] = 44'h00000000000;
    \8052 [483] = 44'h00000000000;
    \8052 [484] = 44'h080001111b1;
    \8052 [485] = 44'h09000110069;
    \8052 [486] = 44'h00000000000;
    \8052 [487] = 44'h090001111b1;
    \8052 [488] = 44'h010602014fe;
    \8052 [489] = 44'h001600814fa;
    \8052 [490] = 44'h00000000000;
    \8052 [491] = 44'h001800814fa;
    \8052 [492] = 44'h00000000000;
    \8052 [493] = 44'h00000000009;
    \8052 [494] = 44'h00000000000;
    \8052 [495] = 44'h00000000000;
    \8052 [496] = 44'h000004814e9;
    \8052 [497] = 44'h00000000000;
    \8052 [498] = 44'h00000000000;
    \8052 [499] = 44'h00000000000;
    \8052 [500] = 44'h09000081359;
    \8052 [501] = 44'h08010081211;
    \8052 [502] = 44'h08000081351;
    \8052 [503] = 44'h0801d081211;
    \8052 [504] = 44'h00000000000;
    \8052 [505] = 44'h00000000000;
    \8052 [506] = 44'h00000000000;
    \8052 [507] = 44'h00000000000;
    \8052 [508] = 44'h00000000000;
    \8052 [509] = 44'h00000000000;
    \8052 [510] = 44'h00000000000;
    \8052 [511] = 44'h00000000000;
    \8052 [512] = 44'h00000000000;
    \8052 [513] = 44'h00000000000;
    \8052 [514] = 44'h00000000000;
    \8052 [515] = 44'h00000111051;
    \8052 [516] = 44'h00000000000;
    \8052 [517] = 44'h00080110169;
    \8052 [518] = 44'h00000000000;
    \8052 [519] = 44'h00000000000;
    \8052 [520] = 44'h00000000000;
    \8052 [521] = 44'h00000000000;
    \8052 [522] = 44'h00000000000;
    \8052 [523] = 44'h00000000000;
    \8052 [524] = 44'h00000000000;
    \8052 [525] = 44'h000000001c2;
    \8052 [526] = 44'h00000000000;
    \8052 [527] = 44'h00000000000;
    \8052 [528] = 44'h000004814e9;
    \8052 [529] = 44'h00000000000;
    \8052 [530] = 44'h00000000000;
    \8052 [531] = 44'h00000000000;
    \8052 [532] = 44'h0b0000812a9;
    \8052 [533] = 44'h00000000000;
    \8052 [534] = 44'h0a0000812a9;
    \8052 [535] = 44'h00000000000;
    \8052 [536] = 44'h00000000000;
    \8052 [537] = 44'h00000000000;
    \8052 [538] = 44'h00000000000;
    \8052 [539] = 44'h00000000000;
    \8052 [540] = 44'h00000000000;
    \8052 [541] = 44'h00000000000;
    \8052 [542] = 44'h00000000000;
    \8052 [543] = 44'h00000000000;
    \8052 [544] = 44'h00000000000;
    \8052 [545] = 44'h00000000000;
    \8052 [546] = 44'h00000000000;
    \8052 [547] = 44'h08002111019;
    \8052 [548] = 44'h00000000000;
    \8052 [549] = 44'h00000000000;
    \8052 [550] = 44'h00000000000;
    \8052 [551] = 44'h00000000000;
    \8052 [552] = 44'h00000000000;
    \8052 [553] = 44'h00000000000;
    \8052 [554] = 44'h00000000000;
    \8052 [555] = 44'h00000000000;
    \8052 [556] = 44'h00000190141;
    \8052 [557] = 44'h00000000000;
    \8052 [558] = 44'h00000000000;
    \8052 [559] = 44'h00000000000;
    \8052 [560] = 44'h000004814e9;
    \8052 [561] = 44'h00000000000;
    \8052 [562] = 44'h00000000000;
    \8052 [563] = 44'h00000000000;
    \8052 [564] = 44'h090000812a9;
    \8052 [565] = 44'h00000000000;
    \8052 [566] = 44'h080000812a9;
    \8052 [567] = 44'h00000000000;
    \8052 [568] = 44'h00000000000;
    \8052 [569] = 44'h00000000000;
    \8052 [570] = 44'h00000000000;
    \8052 [571] = 44'h00000000000;
    \8052 [572] = 44'h00000000000;
    \8052 [573] = 44'h00000000000;
    \8052 [574] = 44'h00000000000;
    \8052 [575] = 44'h00000000000;
    \8052 [576] = 44'h00000000000;
    \8052 [577] = 44'h00000000000;
    \8052 [578] = 44'h00000000000;
    \8052 [579] = 44'h08000111161;
    \8052 [580] = 44'h00000000000;
    \8052 [581] = 44'h00000000000;
    \8052 [582] = 44'h00000000000;
    \8052 [583] = 44'h00000000000;
    \8052 [584] = 44'h00440111502;
    \8052 [585] = 44'h00000000000;
    \8052 [586] = 44'h00000000000;
    \8052 [587] = 44'h00000000000;
    \8052 [588] = 44'h00000000000;
    \8052 [589] = 44'h00000000000;
    \8052 [590] = 44'h00000000000;
    \8052 [591] = 44'h00000000000;
    \8052 [592] = 44'h000004814e9;
    \8052 [593] = 44'h00000000000;
    \8052 [594] = 44'h00000000000;
    \8052 [595] = 44'h00000000000;
    \8052 [596] = 44'h0b0000812b1;
    \8052 [597] = 44'h00000000000;
    \8052 [598] = 44'h0a0000812b1;
    \8052 [599] = 44'h00000000000;
    \8052 [600] = 44'h00000000000;
    \8052 [601] = 44'h00000000000;
    \8052 [602] = 44'h00000000000;
    \8052 [603] = 44'h00000000000;
    \8052 [604] = 44'h00000000000;
    \8052 [605] = 44'h00000000000;
    \8052 [606] = 44'h00000000000;
    \8052 [607] = 44'h00000000000;
    \8052 [608] = 44'h00000000000;
    \8052 [609] = 44'h00000000000;
    \8052 [610] = 44'h00000000000;
    \8052 [611] = 44'h08001111161;
    \8052 [612] = 44'h00000000000;
    \8052 [613] = 44'h00000000000;
    \8052 [614] = 44'h00000000000;
    \8052 [615] = 44'h00000000000;
    \8052 [616] = 44'h00040011502;
    \8052 [617] = 44'h00000000000;
    \8052 [618] = 44'h00000000000;
    \8052 [619] = 44'h00000000000;
    \8052 [620] = 44'h00000000000;
    \8052 [621] = 44'h00000000000;
    \8052 [622] = 44'h00000000000;
    \8052 [623] = 44'h00000000000;
    \8052 [624] = 44'h000004814e9;
    \8052 [625] = 44'h00000000000;
    \8052 [626] = 44'h00000000000;
    \8052 [627] = 44'h00000000000;
    \8052 [628] = 44'h090000812b1;
    \8052 [629] = 44'h00000000000;
    \8052 [630] = 44'h080000812b1;
    \8052 [631] = 44'h00000000000;
    \8052 [632] = 44'h00000000000;
    \8052 [633] = 44'h00000000000;
    \8052 [634] = 44'h00000000000;
    \8052 [635] = 44'h00000000000;
    \8052 [636] = 44'h00000000000;
    \8052 [637] = 44'h00000000000;
    \8052 [638] = 44'h00000000000;
    \8052 [639] = 44'h00000000000;
    \8052 [640] = 44'h00000000000;
    \8052 [641] = 44'h00000000000;
    \8052 [642] = 44'h00000000000;
    \8052 [643] = 44'h00000000000;
    \8052 [644] = 44'h00000000000;
    \8052 [645] = 44'h00060110169;
    \8052 [646] = 44'h00000000000;
    \8052 [647] = 44'h00000000000;
    \8052 [648] = 44'hc06400814fa;
    \8052 [649] = 44'h00000000009;
    \8052 [650] = 44'hc06600814fa;
    \8052 [651] = 44'h00000000000;
    \8052 [652] = 44'h00000000000;
    \8052 [653] = 44'h00000000000;
    \8052 [654] = 44'h00000000000;
    \8052 [655] = 44'h00000000000;
    \8052 [656] = 44'h000004814e9;
    \8052 [657] = 44'h00000000000;
    \8052 [658] = 44'h00000000000;
    \8052 [659] = 44'h00000000000;
    \8052 [660] = 44'h00000000000;
    \8052 [661] = 44'h00000000000;
    \8052 [662] = 44'h00000000000;
    \8052 [663] = 44'h00000000000;
    \8052 [664] = 44'h00000000000;
    \8052 [665] = 44'h00000000000;
    \8052 [666] = 44'h00000000000;
    \8052 [667] = 44'h00000000000;
    \8052 [668] = 44'h00000000000;
    \8052 [669] = 44'h00000000000;
    \8052 [670] = 44'h00000000000;
    \8052 [671] = 44'h00000000000;
    \8052 [672] = 44'h00000000000;
    \8052 [673] = 44'h00000000000;
    \8052 [674] = 44'h00000000000;
    \8052 [675] = 44'h00000000000;
    \8052 [676] = 44'h00000000000;
    \8052 [677] = 44'h00000000000;
    \8052 [678] = 44'h00000000000;
    \8052 [679] = 44'h00000000000;
    \8052 [680] = 44'h002400814fa;
    \8052 [681] = 44'h00000000009;
    \8052 [682] = 44'h002600814fa;
    \8052 [683] = 44'h00000000000;
    \8052 [684] = 44'h00000090721;
    \8052 [685] = 44'h00000000000;
    \8052 [686] = 44'h00000000000;
    \8052 [687] = 44'h00000000000;
    \8052 [688] = 44'h000004814e9;
    \8052 [689] = 44'h00000000000;
    \8052 [690] = 44'h00000000000;
    \8052 [691] = 44'h00000000000;
    \8052 [692] = 44'h00000000000;
    \8052 [693] = 44'h00000000000;
    \8052 [694] = 44'h00000000000;
    \8052 [695] = 44'h00000000000;
    \8052 [696] = 44'h00000000000;
    \8052 [697] = 44'h00000000000;
    \8052 [698] = 44'h00000000000;
    \8052 [699] = 44'h00000000000;
    \8052 [700] = 44'h00000000000;
    \8052 [701] = 44'h00000000000;
    \8052 [702] = 44'h00000000000;
    \8052 [703] = 44'h00000000000;
    \8052 [704] = 44'h00000000000;
    \8052 [705] = 44'h00000000000;
    \8052 [706] = 44'h00000000000;
    \8052 [707] = 44'h080001111d1;
    \8052 [708] = 44'h00000000000;
    \8052 [709] = 44'h000001101d9;
    \8052 [710] = 44'h00000000000;
    \8052 [711] = 44'h00000000000;
    \8052 [712] = 44'hc04400814fa;
    \8052 [713] = 44'h00000000000;
    \8052 [714] = 44'h00000000000;
    \8052 [715] = 44'h00000000000;
    \8052 [716] = 44'h00000000000;
    \8052 [717] = 44'h000000111c2;
    \8052 [718] = 44'h00000000000;
    \8052 [719] = 44'h00000000000;
    \8052 [720] = 44'h000004814e9;
    \8052 [721] = 44'h00000000000;
    \8052 [722] = 44'h00000000000;
    \8052 [723] = 44'h00000000000;
    \8052 [724] = 44'h00000000000;
    \8052 [725] = 44'h00000000000;
    \8052 [726] = 44'h00000000000;
    \8052 [727] = 44'h00000000000;
    \8052 [728] = 44'h00000000000;
    \8052 [729] = 44'h00000000000;
    \8052 [730] = 44'h00000000000;
    \8052 [731] = 44'h00000000000;
    \8052 [732] = 44'h00000000000;
    \8052 [733] = 44'h00000000000;
    \8052 [734] = 44'h00000000000;
    \8052 [735] = 44'h00000000000;
    \8052 [736] = 44'h00000000000;
    \8052 [737] = 44'h00000000000;
    \8052 [738] = 44'h00000000000;
    \8052 [739] = 44'h080021111d1;
    \8052 [740] = 44'h00000000000;
    \8052 [741] = 44'h000011101d9;
    \8052 [742] = 44'h00000000000;
    \8052 [743] = 44'h00000000000;
    \8052 [744] = 44'h000400814fa;
    \8052 [745] = 44'h20000000091;
    \8052 [746] = 44'h00000000000;
    \8052 [747] = 44'h808800814fa;
    \8052 [748] = 44'h00000000000;
    \8052 [749] = 44'h000000111c2;
    \8052 [750] = 44'h00000000000;
    \8052 [751] = 44'h00000000000;
    \8052 [752] = 44'h000004814e9;
    \8052 [753] = 44'h00000000000;
    \8052 [754] = 44'h00000000000;
    \8052 [755] = 44'h00000000000;
    \8052 [756] = 44'h01000081329;
    \8052 [757] = 44'h08000081211;
    \8052 [758] = 44'h00000081329;
    \8052 [759] = 44'h00000000000;
    \8052 [760] = 44'h00000000000;
    \8052 [761] = 44'h00000000000;
    \8052 [762] = 44'h00000000000;
    \8052 [763] = 44'h00000000000;
    \8052 [764] = 44'h00000000000;
    \8052 [765] = 44'h00000000000;
    \8052 [766] = 44'h00000000000;
    \8052 [767] = 44'h00000000000;
    \8052 [768] = 44'h00000000000;
    \8052 [769] = 44'h00000000000;
    \8052 [770] = 44'h00000000000;
    \8052 [771] = 44'h00000111041;
    \8052 [772] = 44'h00000000000;
    \8052 [773] = 44'h00000000000;
    \8052 [774] = 44'h00000000000;
    \8052 [775] = 44'h00000000000;
    \8052 [776] = 44'h00420111502;
    \8052 [777] = 44'h20000000099;
    \8052 [778] = 44'h00000000000;
    \8052 [779] = 44'h00000000000;
    \8052 [780] = 44'h00000000000;
    \8052 [781] = 44'h00000000000;
    \8052 [782] = 44'h00000000000;
    \8052 [783] = 44'h00000000000;
    \8052 [784] = 44'h000004814e9;
    \8052 [785] = 44'h00000000000;
    \8052 [786] = 44'h00000000000;
    \8052 [787] = 44'h00000000000;
    \8052 [788] = 44'h0b000081349;
    \8052 [789] = 44'h0801408b211;
    \8052 [790] = 44'h0a000081349;
    \8052 [791] = 44'h0801508b211;
    \8052 [792] = 44'h00000000000;
    \8052 [793] = 44'h00000000000;
    \8052 [794] = 44'h00000000000;
    \8052 [795] = 44'h00000000000;
    \8052 [796] = 44'h00000000000;
    \8052 [797] = 44'h00000000000;
    \8052 [798] = 44'h00000000000;
    \8052 [799] = 44'h00000801259;
    \8052 [800] = 44'h00000000000;
    \8052 [801] = 44'h00000000000;
    \8052 [802] = 44'h00000000000;
    \8052 [803] = 44'h00000000000;
    \8052 [804] = 44'h00000000000;
    \8052 [805] = 44'h00000000000;
    \8052 [806] = 44'h00000000000;
    \8052 [807] = 44'h00000000000;
    \8052 [808] = 44'h00020011502;
    \8052 [809] = 44'h04880011502;
    \8052 [810] = 44'h00000000000;
    \8052 [811] = 44'h00000000000;
    \8052 [812] = 44'h00000000000;
    \8052 [813] = 44'h00000000000;
    \8052 [814] = 44'h00000000000;
    \8052 [815] = 44'h00000000000;
    \8052 [816] = 44'h000004814e9;
    \8052 [817] = 44'h00000000000;
    \8052 [818] = 44'h00000000000;
    \8052 [819] = 44'h00000000000;
    \8052 [820] = 44'h00000000000;
    \8052 [821] = 44'h08014080211;
    \8052 [822] = 44'h00000000000;
    \8052 [823] = 44'h08015080211;
    \8052 [824] = 44'h00000000000;
    \8052 [825] = 44'h00000000000;
    \8052 [826] = 44'h00000000000;
    \8052 [827] = 44'h00000000000;
    \8052 [828] = 44'h00000000000;
    \8052 [829] = 44'h00000000000;
    \8052 [830] = 44'h00000000000;
    \8052 [831] = 44'h00000801261;
    \8052 [832] = 44'h00000000000;
    \8052 [833] = 44'h00000000000;
    \8052 [834] = 44'h00000000000;
    \8052 [835] = 44'h00000000000;
    \8052 [836] = 44'h00000000000;
    \8052 [837] = 44'h00080110171;
    \8052 [838] = 44'h00000000000;
    \8052 [839] = 44'h00000000000;
    \8052 [840] = 44'h00460111502;
    \8052 [841] = 44'h44880011502;
    \8052 [842] = 44'h00480111502;
    \8052 [843] = 44'h00000000000;
    \8052 [844] = 44'h00000000000;
    \8052 [845] = 44'h20000010139;
    \8052 [846] = 44'h00000000000;
    \8052 [847] = 44'h00000000000;
    \8052 [848] = 44'h000004814e9;
    \8052 [849] = 44'h00000000000;
    \8052 [850] = 44'h00000000000;
    \8052 [851] = 44'h00000000000;
    \8052 [852] = 44'h00000000000;
    \8052 [853] = 44'h08018081211;
    \8052 [854] = 44'h00000000000;
    \8052 [855] = 44'h00000000000;
    \8052 [856] = 44'h00000000000;
    \8052 [857] = 44'h00000000000;
    \8052 [858] = 44'h00000000000;
    \8052 [859] = 44'h00000000000;
    \8052 [860] = 44'h00000000000;
    \8052 [861] = 44'h00000000000;
    \8052 [862] = 44'h00000000000;
    \8052 [863] = 44'h00000000000;
    \8052 [864] = 44'h00000000000;
    \8052 [865] = 44'h00000000000;
    \8052 [866] = 44'h00000000000;
    \8052 [867] = 44'h00000000000;
    \8052 [868] = 44'h00000000000;
    \8052 [869] = 44'h00060110171;
    \8052 [870] = 44'h00000000000;
    \8052 [871] = 44'h00000000000;
    \8052 [872] = 44'h00060011502;
    \8052 [873] = 44'h04860011502;
    \8052 [874] = 44'h00080011502;
    \8052 [875] = 44'h00000000000;
    \8052 [876] = 44'h00000000000;
    \8052 [877] = 44'h21000010139;
    \8052 [878] = 44'h00000000000;
    \8052 [879] = 44'h00000810131;
    \8052 [880] = 44'h000004814e9;
    \8052 [881] = 44'h00000000000;
    \8052 [882] = 44'h00000000000;
    \8052 [883] = 44'h00000000000;
    \8052 [884] = 44'h00000000000;
    \8052 [885] = 44'h08014081211;
    \8052 [886] = 44'h00000000000;
    \8052 [887] = 44'h08015081211;
    \8052 [888] = 44'h00000000000;
    \8052 [889] = 44'h00000000000;
    \8052 [890] = 44'h00000000000;
    \8052 [891] = 44'h00000000000;
    \8052 [892] = 44'h00000000000;
    \8052 [893] = 44'h00000000000;
    \8052 [894] = 44'h00000000000;
    \8052 [895] = 44'h000004801a1;
    \8052 [896] = 44'h00000000000;
    \8052 [897] = 44'h00000000000;
    \8052 [898] = 44'h00000000000;
    \8052 [899] = 44'h08002111161;
    \8052 [900] = 44'h00000000000;
    \8052 [901] = 44'h00020110169;
    \8052 [902] = 44'h00000000000;
    \8052 [903] = 44'h00000000000;
    \8052 [904] = 44'hc04200814fa;
    \8052 [905] = 44'h00000000000;
    \8052 [906] = 44'h00000000000;
    \8052 [907] = 44'h008400814fa;
    \8052 [908] = 44'h00000000000;
    \8052 [909] = 44'h00000000000;
    \8052 [910] = 44'h00000000000;
    \8052 [911] = 44'h00000000000;
    \8052 [912] = 44'h000004814e9;
    \8052 [913] = 44'h00000000000;
    \8052 [914] = 44'h00000000000;
    \8052 [915] = 44'h00000000000;
    \8052 [916] = 44'h00000000000;
    \8052 [917] = 44'h00000000000;
    \8052 [918] = 44'h00000000000;
    \8052 [919] = 44'h0800d080211;
    \8052 [920] = 44'h00000000000;
    \8052 [921] = 44'h00000000000;
    \8052 [922] = 44'h00000000000;
    \8052 [923] = 44'h00000000000;
    \8052 [924] = 44'h00000000000;
    \8052 [925] = 44'h00000000000;
    \8052 [926] = 44'h00000000000;
    \8052 [927] = 44'h00000000000;
    \8052 [928] = 44'h00000000000;
    \8052 [929] = 44'h00000000000;
    \8052 [930] = 44'h00000000000;
    \8052 [931] = 44'h00000000000;
    \8052 [932] = 44'h00000000000;
    \8052 [933] = 44'h00000000000;
    \8052 [934] = 44'h00000000000;
    \8052 [935] = 44'h00000000000;
    \8052 [936] = 44'h000200814fa;
    \8052 [937] = 44'h20000000081;
    \8052 [938] = 44'h00000000000;
    \8052 [939] = 44'h008800814fa;
    \8052 [940] = 44'h20000080119;
    \8052 [941] = 44'h00000000000;
    \8052 [942] = 44'h00000000000;
    \8052 [943] = 44'h00000000000;
    \8052 [944] = 44'h000004814e9;
    \8052 [945] = 44'h00000000000;
    \8052 [946] = 44'h00000000000;
    \8052 [947] = 44'h00000000000;
    \8052 [948] = 44'h0b000081359;
    \8052 [949] = 44'h000000813e1;
    \8052 [950] = 44'h0a000081351;
    \8052 [951] = 44'h00000000000;
    \8052 [952] = 44'h00000000000;
    \8052 [953] = 44'h00000000000;
    \8052 [954] = 44'h00000000000;
    \8052 [955] = 44'h000000013c9;
    \8052 [956] = 44'h00000000000;
    \8052 [957] = 44'h00000000000;
    \8052 [958] = 44'h00000000000;
    \8052 [959] = 44'h00000000000;
    \8052 [960] = 44'h00000000000;
    \8052 [961] = 44'h00000000000;
    \8052 [962] = 44'h00000000000;
    \8052 [963] = 44'h08001111019;
    \8052 [964] = 44'h00000000000;
    \8052 [965] = 44'h08000110069;
    \8052 [966] = 44'h00000000000;
    \8052 [967] = 44'h00000000000;
    \8052 [968] = 44'hc04600814fa;
    \8052 [969] = 44'h20000000089;
    \8052 [970] = 44'hc04800814fa;
    \8052 [971] = 44'h008200814fa;
    \8052 [972] = 44'h00000000000;
    \8052 [973] = 44'h00000000000;
    \8052 [974] = 44'h00000000000;
    \8052 [975] = 44'h00000000000;
    \8052 [976] = 44'h000004814e9;
    \8052 [977] = 44'h00000000000;
    \8052 [978] = 44'h00000000000;
    \8052 [979] = 44'h00000000000;
    \8052 [980] = 44'h00000000000;
    \8052 [981] = 44'h00000000000;
    \8052 [982] = 44'h00000000000;
    \8052 [983] = 44'h0800d081211;
    \8052 [984] = 44'h00000000000;
    \8052 [985] = 44'h00000000000;
    \8052 [986] = 44'h00000000000;
    \8052 [987] = 44'h00000000000;
    \8052 [988] = 44'h00000000000;
    \8052 [989] = 44'h00000000000;
    \8052 [990] = 44'h00000000000;
    \8052 [991] = 44'h0000d801249;
    \8052 [992] = 44'h00000000000;
    \8052 [993] = 44'h20000000009;
    \8052 [994] = 44'h00000000000;
    \8052 [995] = 44'h08000111019;
    \8052 [996] = 44'h080001111a9;
    \8052 [997] = 44'h09000110069;
    \8052 [998] = 44'h00000000000;
    \8052 [999] = 44'h090001111a9;
    \8052 [1000] = 44'h000600814fa;
    \8052 [1001] = 44'h200000000e1;
    \8052 [1002] = 44'h000800814fa;
    \8052 [1003] = 44'h008600814fa;
    \8052 [1004] = 44'h00000480111;
    \8052 [1005] = 44'h00000000000;
    \8052 [1006] = 44'h00000000000;
    \8052 [1007] = 44'h00000000000;
    \8052 [1008] = 44'h000004814e9;
    \8052 [1009] = 44'h00000000000;
    \8052 [1010] = 44'h00000000000;
    \8052 [1011] = 44'h00000000000;
    \8052 [1012] = 44'h09000081359;
    \8052 [1013] = 44'h08010081211;
    \8052 [1014] = 44'h08000081351;
    \8052 [1015] = 44'h0801d081211;
    \8052 [1016] = 44'h00000000000;
    \8052 [1017] = 44'h00000000000;
    \8052 [1018] = 44'h00000000000;
    \8052 [1019] = 44'h010000013c9;
    \8052 [1020] = 44'h00000000000;
    \8052 [1021] = 44'h00000000000;
    \8052 [1022] = 44'h00000000000;
    \8052 [1023] = 44'h0200d801249;
  end
  assign _195_ = \8052 [_037_];
  reg [0:0] \8054  [1023:0];
  initial begin
    \8054 [0] = 1'h0;
    \8054 [1] = 1'h0;
    \8054 [2] = 1'h0;
    \8054 [3] = 1'h0;
    \8054 [4] = 1'h0;
    \8054 [5] = 1'h0;
    \8054 [6] = 1'h0;
    \8054 [7] = 1'h0;
    \8054 [8] = 1'h0;
    \8054 [9] = 1'h0;
    \8054 [10] = 1'h0;
    \8054 [11] = 1'h0;
    \8054 [12] = 1'h0;
    \8054 [13] = 1'h0;
    \8054 [14] = 1'h0;
    \8054 [15] = 1'h0;
    \8054 [16] = 1'h0;
    \8054 [17] = 1'h0;
    \8054 [18] = 1'h0;
    \8054 [19] = 1'h0;
    \8054 [20] = 1'h0;
    \8054 [21] = 1'h0;
    \8054 [22] = 1'h0;
    \8054 [23] = 1'h0;
    \8054 [24] = 1'h0;
    \8054 [25] = 1'h0;
    \8054 [26] = 1'h0;
    \8054 [27] = 1'h0;
    \8054 [28] = 1'h0;
    \8054 [29] = 1'h0;
    \8054 [30] = 1'h0;
    \8054 [31] = 1'h0;
    \8054 [32] = 1'h0;
    \8054 [33] = 1'h0;
    \8054 [34] = 1'h0;
    \8054 [35] = 1'h0;
    \8054 [36] = 1'h0;
    \8054 [37] = 1'h0;
    \8054 [38] = 1'h0;
    \8054 [39] = 1'h0;
    \8054 [40] = 1'h0;
    \8054 [41] = 1'h0;
    \8054 [42] = 1'h0;
    \8054 [43] = 1'h0;
    \8054 [44] = 1'h0;
    \8054 [45] = 1'h0;
    \8054 [46] = 1'h0;
    \8054 [47] = 1'h0;
    \8054 [48] = 1'h0;
    \8054 [49] = 1'h0;
    \8054 [50] = 1'h0;
    \8054 [51] = 1'h0;
    \8054 [52] = 1'h0;
    \8054 [53] = 1'h0;
    \8054 [54] = 1'h0;
    \8054 [55] = 1'h0;
    \8054 [56] = 1'h0;
    \8054 [57] = 1'h0;
    \8054 [58] = 1'h0;
    \8054 [59] = 1'h0;
    \8054 [60] = 1'h0;
    \8054 [61] = 1'h0;
    \8054 [62] = 1'h0;
    \8054 [63] = 1'h0;
    \8054 [64] = 1'h0;
    \8054 [65] = 1'h0;
    \8054 [66] = 1'h0;
    \8054 [67] = 1'h0;
    \8054 [68] = 1'h0;
    \8054 [69] = 1'h0;
    \8054 [70] = 1'h0;
    \8054 [71] = 1'h0;
    \8054 [72] = 1'h0;
    \8054 [73] = 1'h0;
    \8054 [74] = 1'h0;
    \8054 [75] = 1'h0;
    \8054 [76] = 1'h0;
    \8054 [77] = 1'h0;
    \8054 [78] = 1'h0;
    \8054 [79] = 1'h0;
    \8054 [80] = 1'h0;
    \8054 [81] = 1'h0;
    \8054 [82] = 1'h0;
    \8054 [83] = 1'h0;
    \8054 [84] = 1'h0;
    \8054 [85] = 1'h0;
    \8054 [86] = 1'h0;
    \8054 [87] = 1'h0;
    \8054 [88] = 1'h0;
    \8054 [89] = 1'h0;
    \8054 [90] = 1'h0;
    \8054 [91] = 1'h0;
    \8054 [92] = 1'h0;
    \8054 [93] = 1'h0;
    \8054 [94] = 1'h0;
    \8054 [95] = 1'h0;
    \8054 [96] = 1'h0;
    \8054 [97] = 1'h0;
    \8054 [98] = 1'h0;
    \8054 [99] = 1'h0;
    \8054 [100] = 1'h0;
    \8054 [101] = 1'h0;
    \8054 [102] = 1'h0;
    \8054 [103] = 1'h0;
    \8054 [104] = 1'h0;
    \8054 [105] = 1'h0;
    \8054 [106] = 1'h0;
    \8054 [107] = 1'h0;
    \8054 [108] = 1'h0;
    \8054 [109] = 1'h0;
    \8054 [110] = 1'h0;
    \8054 [111] = 1'h0;
    \8054 [112] = 1'h0;
    \8054 [113] = 1'h0;
    \8054 [114] = 1'h0;
    \8054 [115] = 1'h0;
    \8054 [116] = 1'h0;
    \8054 [117] = 1'h0;
    \8054 [118] = 1'h0;
    \8054 [119] = 1'h0;
    \8054 [120] = 1'h0;
    \8054 [121] = 1'h0;
    \8054 [122] = 1'h0;
    \8054 [123] = 1'h0;
    \8054 [124] = 1'h0;
    \8054 [125] = 1'h0;
    \8054 [126] = 1'h0;
    \8054 [127] = 1'h0;
    \8054 [128] = 1'h0;
    \8054 [129] = 1'h0;
    \8054 [130] = 1'h0;
    \8054 [131] = 1'h0;
    \8054 [132] = 1'h0;
    \8054 [133] = 1'h0;
    \8054 [134] = 1'h0;
    \8054 [135] = 1'h0;
    \8054 [136] = 1'h0;
    \8054 [137] = 1'h0;
    \8054 [138] = 1'h0;
    \8054 [139] = 1'h0;
    \8054 [140] = 1'h0;
    \8054 [141] = 1'h0;
    \8054 [142] = 1'h0;
    \8054 [143] = 1'h0;
    \8054 [144] = 1'h0;
    \8054 [145] = 1'h0;
    \8054 [146] = 1'h0;
    \8054 [147] = 1'h0;
    \8054 [148] = 1'h0;
    \8054 [149] = 1'h0;
    \8054 [150] = 1'h0;
    \8054 [151] = 1'h0;
    \8054 [152] = 1'h0;
    \8054 [153] = 1'h0;
    \8054 [154] = 1'h0;
    \8054 [155] = 1'h0;
    \8054 [156] = 1'h0;
    \8054 [157] = 1'h0;
    \8054 [158] = 1'h0;
    \8054 [159] = 1'h0;
    \8054 [160] = 1'h0;
    \8054 [161] = 1'h0;
    \8054 [162] = 1'h0;
    \8054 [163] = 1'h0;
    \8054 [164] = 1'h0;
    \8054 [165] = 1'h0;
    \8054 [166] = 1'h0;
    \8054 [167] = 1'h0;
    \8054 [168] = 1'h0;
    \8054 [169] = 1'h0;
    \8054 [170] = 1'h0;
    \8054 [171] = 1'h0;
    \8054 [172] = 1'h0;
    \8054 [173] = 1'h0;
    \8054 [174] = 1'h0;
    \8054 [175] = 1'h0;
    \8054 [176] = 1'h0;
    \8054 [177] = 1'h0;
    \8054 [178] = 1'h0;
    \8054 [179] = 1'h0;
    \8054 [180] = 1'h0;
    \8054 [181] = 1'h0;
    \8054 [182] = 1'h0;
    \8054 [183] = 1'h0;
    \8054 [184] = 1'h0;
    \8054 [185] = 1'h0;
    \8054 [186] = 1'h0;
    \8054 [187] = 1'h0;
    \8054 [188] = 1'h0;
    \8054 [189] = 1'h0;
    \8054 [190] = 1'h0;
    \8054 [191] = 1'h0;
    \8054 [192] = 1'h0;
    \8054 [193] = 1'h0;
    \8054 [194] = 1'h0;
    \8054 [195] = 1'h0;
    \8054 [196] = 1'h0;
    \8054 [197] = 1'h0;
    \8054 [198] = 1'h0;
    \8054 [199] = 1'h0;
    \8054 [200] = 1'h0;
    \8054 [201] = 1'h0;
    \8054 [202] = 1'h0;
    \8054 [203] = 1'h0;
    \8054 [204] = 1'h0;
    \8054 [205] = 1'h0;
    \8054 [206] = 1'h0;
    \8054 [207] = 1'h0;
    \8054 [208] = 1'h0;
    \8054 [209] = 1'h0;
    \8054 [210] = 1'h0;
    \8054 [211] = 1'h0;
    \8054 [212] = 1'h0;
    \8054 [213] = 1'h0;
    \8054 [214] = 1'h0;
    \8054 [215] = 1'h0;
    \8054 [216] = 1'h0;
    \8054 [217] = 1'h0;
    \8054 [218] = 1'h0;
    \8054 [219] = 1'h0;
    \8054 [220] = 1'h0;
    \8054 [221] = 1'h0;
    \8054 [222] = 1'h0;
    \8054 [223] = 1'h0;
    \8054 [224] = 1'h0;
    \8054 [225] = 1'h0;
    \8054 [226] = 1'h0;
    \8054 [227] = 1'h0;
    \8054 [228] = 1'h0;
    \8054 [229] = 1'h0;
    \8054 [230] = 1'h0;
    \8054 [231] = 1'h0;
    \8054 [232] = 1'h0;
    \8054 [233] = 1'h0;
    \8054 [234] = 1'h0;
    \8054 [235] = 1'h0;
    \8054 [236] = 1'h0;
    \8054 [237] = 1'h0;
    \8054 [238] = 1'h0;
    \8054 [239] = 1'h0;
    \8054 [240] = 1'h0;
    \8054 [241] = 1'h0;
    \8054 [242] = 1'h0;
    \8054 [243] = 1'h0;
    \8054 [244] = 1'h0;
    \8054 [245] = 1'h0;
    \8054 [246] = 1'h0;
    \8054 [247] = 1'h0;
    \8054 [248] = 1'h0;
    \8054 [249] = 1'h0;
    \8054 [250] = 1'h0;
    \8054 [251] = 1'h0;
    \8054 [252] = 1'h0;
    \8054 [253] = 1'h0;
    \8054 [254] = 1'h0;
    \8054 [255] = 1'h0;
    \8054 [256] = 1'h0;
    \8054 [257] = 1'h0;
    \8054 [258] = 1'h0;
    \8054 [259] = 1'h0;
    \8054 [260] = 1'h0;
    \8054 [261] = 1'h0;
    \8054 [262] = 1'h0;
    \8054 [263] = 1'h0;
    \8054 [264] = 1'h0;
    \8054 [265] = 1'h0;
    \8054 [266] = 1'h0;
    \8054 [267] = 1'h0;
    \8054 [268] = 1'h0;
    \8054 [269] = 1'h0;
    \8054 [270] = 1'h0;
    \8054 [271] = 1'h0;
    \8054 [272] = 1'h0;
    \8054 [273] = 1'h0;
    \8054 [274] = 1'h0;
    \8054 [275] = 1'h0;
    \8054 [276] = 1'h0;
    \8054 [277] = 1'h0;
    \8054 [278] = 1'h0;
    \8054 [279] = 1'h0;
    \8054 [280] = 1'h0;
    \8054 [281] = 1'h0;
    \8054 [282] = 1'h0;
    \8054 [283] = 1'h0;
    \8054 [284] = 1'h0;
    \8054 [285] = 1'h0;
    \8054 [286] = 1'h0;
    \8054 [287] = 1'h0;
    \8054 [288] = 1'h0;
    \8054 [289] = 1'h0;
    \8054 [290] = 1'h0;
    \8054 [291] = 1'h0;
    \8054 [292] = 1'h0;
    \8054 [293] = 1'h0;
    \8054 [294] = 1'h0;
    \8054 [295] = 1'h0;
    \8054 [296] = 1'h0;
    \8054 [297] = 1'h0;
    \8054 [298] = 1'h0;
    \8054 [299] = 1'h0;
    \8054 [300] = 1'h0;
    \8054 [301] = 1'h0;
    \8054 [302] = 1'h0;
    \8054 [303] = 1'h0;
    \8054 [304] = 1'h0;
    \8054 [305] = 1'h0;
    \8054 [306] = 1'h0;
    \8054 [307] = 1'h0;
    \8054 [308] = 1'h0;
    \8054 [309] = 1'h0;
    \8054 [310] = 1'h0;
    \8054 [311] = 1'h0;
    \8054 [312] = 1'h0;
    \8054 [313] = 1'h0;
    \8054 [314] = 1'h0;
    \8054 [315] = 1'h1;
    \8054 [316] = 1'h0;
    \8054 [317] = 1'h0;
    \8054 [318] = 1'h0;
    \8054 [319] = 1'h0;
    \8054 [320] = 1'h0;
    \8054 [321] = 1'h0;
    \8054 [322] = 1'h0;
    \8054 [323] = 1'h0;
    \8054 [324] = 1'h0;
    \8054 [325] = 1'h0;
    \8054 [326] = 1'h0;
    \8054 [327] = 1'h0;
    \8054 [328] = 1'h0;
    \8054 [329] = 1'h0;
    \8054 [330] = 1'h0;
    \8054 [331] = 1'h0;
    \8054 [332] = 1'h0;
    \8054 [333] = 1'h0;
    \8054 [334] = 1'h0;
    \8054 [335] = 1'h0;
    \8054 [336] = 1'h0;
    \8054 [337] = 1'h0;
    \8054 [338] = 1'h0;
    \8054 [339] = 1'h0;
    \8054 [340] = 1'h0;
    \8054 [341] = 1'h0;
    \8054 [342] = 1'h0;
    \8054 [343] = 1'h0;
    \8054 [344] = 1'h0;
    \8054 [345] = 1'h0;
    \8054 [346] = 1'h0;
    \8054 [347] = 1'h0;
    \8054 [348] = 1'h0;
    \8054 [349] = 1'h0;
    \8054 [350] = 1'h0;
    \8054 [351] = 1'h0;
    \8054 [352] = 1'h0;
    \8054 [353] = 1'h0;
    \8054 [354] = 1'h0;
    \8054 [355] = 1'h0;
    \8054 [356] = 1'h0;
    \8054 [357] = 1'h0;
    \8054 [358] = 1'h0;
    \8054 [359] = 1'h0;
    \8054 [360] = 1'h0;
    \8054 [361] = 1'h0;
    \8054 [362] = 1'h0;
    \8054 [363] = 1'h0;
    \8054 [364] = 1'h0;
    \8054 [365] = 1'h0;
    \8054 [366] = 1'h0;
    \8054 [367] = 1'h0;
    \8054 [368] = 1'h0;
    \8054 [369] = 1'h0;
    \8054 [370] = 1'h0;
    \8054 [371] = 1'h0;
    \8054 [372] = 1'h0;
    \8054 [373] = 1'h0;
    \8054 [374] = 1'h0;
    \8054 [375] = 1'h0;
    \8054 [376] = 1'h0;
    \8054 [377] = 1'h0;
    \8054 [378] = 1'h0;
    \8054 [379] = 1'h0;
    \8054 [380] = 1'h0;
    \8054 [381] = 1'h0;
    \8054 [382] = 1'h0;
    \8054 [383] = 1'h0;
    \8054 [384] = 1'h0;
    \8054 [385] = 1'h0;
    \8054 [386] = 1'h0;
    \8054 [387] = 1'h0;
    \8054 [388] = 1'h0;
    \8054 [389] = 1'h0;
    \8054 [390] = 1'h0;
    \8054 [391] = 1'h0;
    \8054 [392] = 1'h0;
    \8054 [393] = 1'h0;
    \8054 [394] = 1'h0;
    \8054 [395] = 1'h0;
    \8054 [396] = 1'h0;
    \8054 [397] = 1'h0;
    \8054 [398] = 1'h0;
    \8054 [399] = 1'h0;
    \8054 [400] = 1'h0;
    \8054 [401] = 1'h0;
    \8054 [402] = 1'h0;
    \8054 [403] = 1'h0;
    \8054 [404] = 1'h0;
    \8054 [405] = 1'h0;
    \8054 [406] = 1'h0;
    \8054 [407] = 1'h0;
    \8054 [408] = 1'h0;
    \8054 [409] = 1'h0;
    \8054 [410] = 1'h0;
    \8054 [411] = 1'h0;
    \8054 [412] = 1'h0;
    \8054 [413] = 1'h0;
    \8054 [414] = 1'h0;
    \8054 [415] = 1'h0;
    \8054 [416] = 1'h0;
    \8054 [417] = 1'h0;
    \8054 [418] = 1'h0;
    \8054 [419] = 1'h0;
    \8054 [420] = 1'h0;
    \8054 [421] = 1'h0;
    \8054 [422] = 1'h0;
    \8054 [423] = 1'h0;
    \8054 [424] = 1'h0;
    \8054 [425] = 1'h0;
    \8054 [426] = 1'h0;
    \8054 [427] = 1'h0;
    \8054 [428] = 1'h0;
    \8054 [429] = 1'h0;
    \8054 [430] = 1'h0;
    \8054 [431] = 1'h0;
    \8054 [432] = 1'h0;
    \8054 [433] = 1'h0;
    \8054 [434] = 1'h0;
    \8054 [435] = 1'h0;
    \8054 [436] = 1'h0;
    \8054 [437] = 1'h0;
    \8054 [438] = 1'h0;
    \8054 [439] = 1'h0;
    \8054 [440] = 1'h0;
    \8054 [441] = 1'h0;
    \8054 [442] = 1'h0;
    \8054 [443] = 1'h0;
    \8054 [444] = 1'h0;
    \8054 [445] = 1'h0;
    \8054 [446] = 1'h0;
    \8054 [447] = 1'h1;
    \8054 [448] = 1'h0;
    \8054 [449] = 1'h0;
    \8054 [450] = 1'h0;
    \8054 [451] = 1'h0;
    \8054 [452] = 1'h0;
    \8054 [453] = 1'h0;
    \8054 [454] = 1'h0;
    \8054 [455] = 1'h0;
    \8054 [456] = 1'h0;
    \8054 [457] = 1'h0;
    \8054 [458] = 1'h0;
    \8054 [459] = 1'h0;
    \8054 [460] = 1'h0;
    \8054 [461] = 1'h0;
    \8054 [462] = 1'h0;
    \8054 [463] = 1'h0;
    \8054 [464] = 1'h0;
    \8054 [465] = 1'h0;
    \8054 [466] = 1'h0;
    \8054 [467] = 1'h0;
    \8054 [468] = 1'h0;
    \8054 [469] = 1'h0;
    \8054 [470] = 1'h0;
    \8054 [471] = 1'h0;
    \8054 [472] = 1'h0;
    \8054 [473] = 1'h0;
    \8054 [474] = 1'h0;
    \8054 [475] = 1'h0;
    \8054 [476] = 1'h0;
    \8054 [477] = 1'h0;
    \8054 [478] = 1'h0;
    \8054 [479] = 1'h0;
    \8054 [480] = 1'h0;
    \8054 [481] = 1'h0;
    \8054 [482] = 1'h0;
    \8054 [483] = 1'h0;
    \8054 [484] = 1'h0;
    \8054 [485] = 1'h0;
    \8054 [486] = 1'h0;
    \8054 [487] = 1'h0;
    \8054 [488] = 1'h0;
    \8054 [489] = 1'h0;
    \8054 [490] = 1'h0;
    \8054 [491] = 1'h0;
    \8054 [492] = 1'h0;
    \8054 [493] = 1'h0;
    \8054 [494] = 1'h1;
    \8054 [495] = 1'h1;
    \8054 [496] = 1'h0;
    \8054 [497] = 1'h0;
    \8054 [498] = 1'h0;
    \8054 [499] = 1'h0;
    \8054 [500] = 1'h0;
    \8054 [501] = 1'h0;
    \8054 [502] = 1'h0;
    \8054 [503] = 1'h0;
    \8054 [504] = 1'h0;
    \8054 [505] = 1'h0;
    \8054 [506] = 1'h0;
    \8054 [507] = 1'h0;
    \8054 [508] = 1'h0;
    \8054 [509] = 1'h0;
    \8054 [510] = 1'h0;
    \8054 [511] = 1'h1;
    \8054 [512] = 1'h0;
    \8054 [513] = 1'h0;
    \8054 [514] = 1'h0;
    \8054 [515] = 1'h0;
    \8054 [516] = 1'h0;
    \8054 [517] = 1'h0;
    \8054 [518] = 1'h0;
    \8054 [519] = 1'h0;
    \8054 [520] = 1'h0;
    \8054 [521] = 1'h0;
    \8054 [522] = 1'h0;
    \8054 [523] = 1'h0;
    \8054 [524] = 1'h0;
    \8054 [525] = 1'h0;
    \8054 [526] = 1'h0;
    \8054 [527] = 1'h0;
    \8054 [528] = 1'h0;
    \8054 [529] = 1'h0;
    \8054 [530] = 1'h0;
    \8054 [531] = 1'h0;
    \8054 [532] = 1'h0;
    \8054 [533] = 1'h0;
    \8054 [534] = 1'h0;
    \8054 [535] = 1'h0;
    \8054 [536] = 1'h0;
    \8054 [537] = 1'h0;
    \8054 [538] = 1'h0;
    \8054 [539] = 1'h0;
    \8054 [540] = 1'h0;
    \8054 [541] = 1'h0;
    \8054 [542] = 1'h0;
    \8054 [543] = 1'h0;
    \8054 [544] = 1'h0;
    \8054 [545] = 1'h0;
    \8054 [546] = 1'h0;
    \8054 [547] = 1'h0;
    \8054 [548] = 1'h0;
    \8054 [549] = 1'h0;
    \8054 [550] = 1'h0;
    \8054 [551] = 1'h0;
    \8054 [552] = 1'h0;
    \8054 [553] = 1'h0;
    \8054 [554] = 1'h0;
    \8054 [555] = 1'h0;
    \8054 [556] = 1'h0;
    \8054 [557] = 1'h0;
    \8054 [558] = 1'h0;
    \8054 [559] = 1'h0;
    \8054 [560] = 1'h0;
    \8054 [561] = 1'h0;
    \8054 [562] = 1'h0;
    \8054 [563] = 1'h0;
    \8054 [564] = 1'h0;
    \8054 [565] = 1'h0;
    \8054 [566] = 1'h0;
    \8054 [567] = 1'h0;
    \8054 [568] = 1'h0;
    \8054 [569] = 1'h0;
    \8054 [570] = 1'h0;
    \8054 [571] = 1'h0;
    \8054 [572] = 1'h0;
    \8054 [573] = 1'h0;
    \8054 [574] = 1'h0;
    \8054 [575] = 1'h0;
    \8054 [576] = 1'h0;
    \8054 [577] = 1'h0;
    \8054 [578] = 1'h0;
    \8054 [579] = 1'h0;
    \8054 [580] = 1'h0;
    \8054 [581] = 1'h0;
    \8054 [582] = 1'h0;
    \8054 [583] = 1'h0;
    \8054 [584] = 1'h0;
    \8054 [585] = 1'h0;
    \8054 [586] = 1'h0;
    \8054 [587] = 1'h0;
    \8054 [588] = 1'h0;
    \8054 [589] = 1'h0;
    \8054 [590] = 1'h0;
    \8054 [591] = 1'h0;
    \8054 [592] = 1'h0;
    \8054 [593] = 1'h0;
    \8054 [594] = 1'h0;
    \8054 [595] = 1'h0;
    \8054 [596] = 1'h0;
    \8054 [597] = 1'h0;
    \8054 [598] = 1'h0;
    \8054 [599] = 1'h0;
    \8054 [600] = 1'h0;
    \8054 [601] = 1'h0;
    \8054 [602] = 1'h0;
    \8054 [603] = 1'h0;
    \8054 [604] = 1'h0;
    \8054 [605] = 1'h0;
    \8054 [606] = 1'h0;
    \8054 [607] = 1'h0;
    \8054 [608] = 1'h0;
    \8054 [609] = 1'h0;
    \8054 [610] = 1'h0;
    \8054 [611] = 1'h0;
    \8054 [612] = 1'h0;
    \8054 [613] = 1'h0;
    \8054 [614] = 1'h0;
    \8054 [615] = 1'h0;
    \8054 [616] = 1'h0;
    \8054 [617] = 1'h0;
    \8054 [618] = 1'h0;
    \8054 [619] = 1'h0;
    \8054 [620] = 1'h0;
    \8054 [621] = 1'h0;
    \8054 [622] = 1'h0;
    \8054 [623] = 1'h0;
    \8054 [624] = 1'h0;
    \8054 [625] = 1'h0;
    \8054 [626] = 1'h0;
    \8054 [627] = 1'h0;
    \8054 [628] = 1'h0;
    \8054 [629] = 1'h0;
    \8054 [630] = 1'h0;
    \8054 [631] = 1'h0;
    \8054 [632] = 1'h0;
    \8054 [633] = 1'h0;
    \8054 [634] = 1'h0;
    \8054 [635] = 1'h0;
    \8054 [636] = 1'h0;
    \8054 [637] = 1'h0;
    \8054 [638] = 1'h0;
    \8054 [639] = 1'h0;
    \8054 [640] = 1'h0;
    \8054 [641] = 1'h0;
    \8054 [642] = 1'h0;
    \8054 [643] = 1'h0;
    \8054 [644] = 1'h0;
    \8054 [645] = 1'h0;
    \8054 [646] = 1'h0;
    \8054 [647] = 1'h0;
    \8054 [648] = 1'h0;
    \8054 [649] = 1'h0;
    \8054 [650] = 1'h0;
    \8054 [651] = 1'h0;
    \8054 [652] = 1'h0;
    \8054 [653] = 1'h0;
    \8054 [654] = 1'h0;
    \8054 [655] = 1'h0;
    \8054 [656] = 1'h0;
    \8054 [657] = 1'h0;
    \8054 [658] = 1'h0;
    \8054 [659] = 1'h0;
    \8054 [660] = 1'h0;
    \8054 [661] = 1'h0;
    \8054 [662] = 1'h0;
    \8054 [663] = 1'h0;
    \8054 [664] = 1'h0;
    \8054 [665] = 1'h0;
    \8054 [666] = 1'h0;
    \8054 [667] = 1'h0;
    \8054 [668] = 1'h0;
    \8054 [669] = 1'h0;
    \8054 [670] = 1'h0;
    \8054 [671] = 1'h0;
    \8054 [672] = 1'h0;
    \8054 [673] = 1'h0;
    \8054 [674] = 1'h0;
    \8054 [675] = 1'h0;
    \8054 [676] = 1'h0;
    \8054 [677] = 1'h0;
    \8054 [678] = 1'h0;
    \8054 [679] = 1'h0;
    \8054 [680] = 1'h0;
    \8054 [681] = 1'h0;
    \8054 [682] = 1'h0;
    \8054 [683] = 1'h0;
    \8054 [684] = 1'h0;
    \8054 [685] = 1'h0;
    \8054 [686] = 1'h0;
    \8054 [687] = 1'h0;
    \8054 [688] = 1'h0;
    \8054 [689] = 1'h0;
    \8054 [690] = 1'h0;
    \8054 [691] = 1'h0;
    \8054 [692] = 1'h0;
    \8054 [693] = 1'h0;
    \8054 [694] = 1'h0;
    \8054 [695] = 1'h0;
    \8054 [696] = 1'h0;
    \8054 [697] = 1'h0;
    \8054 [698] = 1'h0;
    \8054 [699] = 1'h0;
    \8054 [700] = 1'h0;
    \8054 [701] = 1'h0;
    \8054 [702] = 1'h0;
    \8054 [703] = 1'h0;
    \8054 [704] = 1'h0;
    \8054 [705] = 1'h0;
    \8054 [706] = 1'h0;
    \8054 [707] = 1'h0;
    \8054 [708] = 1'h0;
    \8054 [709] = 1'h0;
    \8054 [710] = 1'h0;
    \8054 [711] = 1'h0;
    \8054 [712] = 1'h0;
    \8054 [713] = 1'h0;
    \8054 [714] = 1'h0;
    \8054 [715] = 1'h0;
    \8054 [716] = 1'h0;
    \8054 [717] = 1'h0;
    \8054 [718] = 1'h0;
    \8054 [719] = 1'h0;
    \8054 [720] = 1'h0;
    \8054 [721] = 1'h0;
    \8054 [722] = 1'h0;
    \8054 [723] = 1'h0;
    \8054 [724] = 1'h0;
    \8054 [725] = 1'h0;
    \8054 [726] = 1'h0;
    \8054 [727] = 1'h0;
    \8054 [728] = 1'h0;
    \8054 [729] = 1'h0;
    \8054 [730] = 1'h0;
    \8054 [731] = 1'h0;
    \8054 [732] = 1'h0;
    \8054 [733] = 1'h0;
    \8054 [734] = 1'h0;
    \8054 [735] = 1'h0;
    \8054 [736] = 1'h0;
    \8054 [737] = 1'h0;
    \8054 [738] = 1'h0;
    \8054 [739] = 1'h0;
    \8054 [740] = 1'h0;
    \8054 [741] = 1'h0;
    \8054 [742] = 1'h0;
    \8054 [743] = 1'h0;
    \8054 [744] = 1'h0;
    \8054 [745] = 1'h0;
    \8054 [746] = 1'h0;
    \8054 [747] = 1'h0;
    \8054 [748] = 1'h0;
    \8054 [749] = 1'h0;
    \8054 [750] = 1'h0;
    \8054 [751] = 1'h0;
    \8054 [752] = 1'h0;
    \8054 [753] = 1'h0;
    \8054 [754] = 1'h0;
    \8054 [755] = 1'h0;
    \8054 [756] = 1'h0;
    \8054 [757] = 1'h0;
    \8054 [758] = 1'h0;
    \8054 [759] = 1'h0;
    \8054 [760] = 1'h0;
    \8054 [761] = 1'h0;
    \8054 [762] = 1'h0;
    \8054 [763] = 1'h0;
    \8054 [764] = 1'h0;
    \8054 [765] = 1'h0;
    \8054 [766] = 1'h0;
    \8054 [767] = 1'h0;
    \8054 [768] = 1'h0;
    \8054 [769] = 1'h0;
    \8054 [770] = 1'h0;
    \8054 [771] = 1'h0;
    \8054 [772] = 1'h0;
    \8054 [773] = 1'h0;
    \8054 [774] = 1'h0;
    \8054 [775] = 1'h0;
    \8054 [776] = 1'h0;
    \8054 [777] = 1'h0;
    \8054 [778] = 1'h0;
    \8054 [779] = 1'h0;
    \8054 [780] = 1'h0;
    \8054 [781] = 1'h0;
    \8054 [782] = 1'h0;
    \8054 [783] = 1'h0;
    \8054 [784] = 1'h0;
    \8054 [785] = 1'h0;
    \8054 [786] = 1'h0;
    \8054 [787] = 1'h0;
    \8054 [788] = 1'h0;
    \8054 [789] = 1'h0;
    \8054 [790] = 1'h0;
    \8054 [791] = 1'h0;
    \8054 [792] = 1'h0;
    \8054 [793] = 1'h0;
    \8054 [794] = 1'h0;
    \8054 [795] = 1'h0;
    \8054 [796] = 1'h0;
    \8054 [797] = 1'h0;
    \8054 [798] = 1'h0;
    \8054 [799] = 1'h0;
    \8054 [800] = 1'h0;
    \8054 [801] = 1'h0;
    \8054 [802] = 1'h0;
    \8054 [803] = 1'h0;
    \8054 [804] = 1'h0;
    \8054 [805] = 1'h0;
    \8054 [806] = 1'h0;
    \8054 [807] = 1'h0;
    \8054 [808] = 1'h0;
    \8054 [809] = 1'h0;
    \8054 [810] = 1'h0;
    \8054 [811] = 1'h0;
    \8054 [812] = 1'h0;
    \8054 [813] = 1'h0;
    \8054 [814] = 1'h0;
    \8054 [815] = 1'h0;
    \8054 [816] = 1'h0;
    \8054 [817] = 1'h0;
    \8054 [818] = 1'h0;
    \8054 [819] = 1'h0;
    \8054 [820] = 1'h0;
    \8054 [821] = 1'h0;
    \8054 [822] = 1'h0;
    \8054 [823] = 1'h0;
    \8054 [824] = 1'h0;
    \8054 [825] = 1'h0;
    \8054 [826] = 1'h0;
    \8054 [827] = 1'h0;
    \8054 [828] = 1'h0;
    \8054 [829] = 1'h0;
    \8054 [830] = 1'h0;
    \8054 [831] = 1'h0;
    \8054 [832] = 1'h0;
    \8054 [833] = 1'h0;
    \8054 [834] = 1'h0;
    \8054 [835] = 1'h0;
    \8054 [836] = 1'h0;
    \8054 [837] = 1'h0;
    \8054 [838] = 1'h0;
    \8054 [839] = 1'h0;
    \8054 [840] = 1'h0;
    \8054 [841] = 1'h0;
    \8054 [842] = 1'h0;
    \8054 [843] = 1'h0;
    \8054 [844] = 1'h0;
    \8054 [845] = 1'h0;
    \8054 [846] = 1'h0;
    \8054 [847] = 1'h0;
    \8054 [848] = 1'h0;
    \8054 [849] = 1'h0;
    \8054 [850] = 1'h0;
    \8054 [851] = 1'h0;
    \8054 [852] = 1'h0;
    \8054 [853] = 1'h0;
    \8054 [854] = 1'h0;
    \8054 [855] = 1'h0;
    \8054 [856] = 1'h0;
    \8054 [857] = 1'h0;
    \8054 [858] = 1'h0;
    \8054 [859] = 1'h0;
    \8054 [860] = 1'h0;
    \8054 [861] = 1'h0;
    \8054 [862] = 1'h0;
    \8054 [863] = 1'h0;
    \8054 [864] = 1'h0;
    \8054 [865] = 1'h0;
    \8054 [866] = 1'h0;
    \8054 [867] = 1'h0;
    \8054 [868] = 1'h0;
    \8054 [869] = 1'h0;
    \8054 [870] = 1'h0;
    \8054 [871] = 1'h0;
    \8054 [872] = 1'h0;
    \8054 [873] = 1'h0;
    \8054 [874] = 1'h0;
    \8054 [875] = 1'h0;
    \8054 [876] = 1'h0;
    \8054 [877] = 1'h0;
    \8054 [878] = 1'h0;
    \8054 [879] = 1'h0;
    \8054 [880] = 1'h0;
    \8054 [881] = 1'h0;
    \8054 [882] = 1'h0;
    \8054 [883] = 1'h0;
    \8054 [884] = 1'h0;
    \8054 [885] = 1'h0;
    \8054 [886] = 1'h0;
    \8054 [887] = 1'h0;
    \8054 [888] = 1'h0;
    \8054 [889] = 1'h0;
    \8054 [890] = 1'h0;
    \8054 [891] = 1'h0;
    \8054 [892] = 1'h0;
    \8054 [893] = 1'h0;
    \8054 [894] = 1'h0;
    \8054 [895] = 1'h0;
    \8054 [896] = 1'h0;
    \8054 [897] = 1'h0;
    \8054 [898] = 1'h0;
    \8054 [899] = 1'h0;
    \8054 [900] = 1'h0;
    \8054 [901] = 1'h0;
    \8054 [902] = 1'h0;
    \8054 [903] = 1'h0;
    \8054 [904] = 1'h0;
    \8054 [905] = 1'h0;
    \8054 [906] = 1'h0;
    \8054 [907] = 1'h0;
    \8054 [908] = 1'h0;
    \8054 [909] = 1'h0;
    \8054 [910] = 1'h0;
    \8054 [911] = 1'h0;
    \8054 [912] = 1'h0;
    \8054 [913] = 1'h0;
    \8054 [914] = 1'h0;
    \8054 [915] = 1'h0;
    \8054 [916] = 1'h0;
    \8054 [917] = 1'h0;
    \8054 [918] = 1'h0;
    \8054 [919] = 1'h0;
    \8054 [920] = 1'h0;
    \8054 [921] = 1'h0;
    \8054 [922] = 1'h0;
    \8054 [923] = 1'h0;
    \8054 [924] = 1'h0;
    \8054 [925] = 1'h0;
    \8054 [926] = 1'h0;
    \8054 [927] = 1'h0;
    \8054 [928] = 1'h1;
    \8054 [929] = 1'h1;
    \8054 [930] = 1'h1;
    \8054 [931] = 1'h1;
    \8054 [932] = 1'h1;
    \8054 [933] = 1'h1;
    \8054 [934] = 1'h1;
    \8054 [935] = 1'h1;
    \8054 [936] = 1'h1;
    \8054 [937] = 1'h1;
    \8054 [938] = 1'h1;
    \8054 [939] = 1'h1;
    \8054 [940] = 1'h1;
    \8054 [941] = 1'h1;
    \8054 [942] = 1'h1;
    \8054 [943] = 1'h1;
    \8054 [944] = 1'h1;
    \8054 [945] = 1'h1;
    \8054 [946] = 1'h1;
    \8054 [947] = 1'h1;
    \8054 [948] = 1'h1;
    \8054 [949] = 1'h1;
    \8054 [950] = 1'h1;
    \8054 [951] = 1'h1;
    \8054 [952] = 1'h1;
    \8054 [953] = 1'h1;
    \8054 [954] = 1'h1;
    \8054 [955] = 1'h1;
    \8054 [956] = 1'h1;
    \8054 [957] = 1'h1;
    \8054 [958] = 1'h1;
    \8054 [959] = 1'h1;
    \8054 [960] = 1'h0;
    \8054 [961] = 1'h0;
    \8054 [962] = 1'h0;
    \8054 [963] = 1'h0;
    \8054 [964] = 1'h0;
    \8054 [965] = 1'h0;
    \8054 [966] = 1'h0;
    \8054 [967] = 1'h0;
    \8054 [968] = 1'h0;
    \8054 [969] = 1'h0;
    \8054 [970] = 1'h0;
    \8054 [971] = 1'h0;
    \8054 [972] = 1'h0;
    \8054 [973] = 1'h0;
    \8054 [974] = 1'h0;
    \8054 [975] = 1'h0;
    \8054 [976] = 1'h0;
    \8054 [977] = 1'h1;
    \8054 [978] = 1'h1;
    \8054 [979] = 1'h0;
    \8054 [980] = 1'h0;
    \8054 [981] = 1'h0;
    \8054 [982] = 1'h1;
    \8054 [983] = 1'h1;
    \8054 [984] = 1'h1;
    \8054 [985] = 1'h1;
    \8054 [986] = 1'h0;
    \8054 [987] = 1'h1;
    \8054 [988] = 1'h0;
    \8054 [989] = 1'h0;
    \8054 [990] = 1'h1;
    \8054 [991] = 1'h0;
    \8054 [992] = 1'h0;
    \8054 [993] = 1'h0;
    \8054 [994] = 1'h0;
    \8054 [995] = 1'h0;
    \8054 [996] = 1'h0;
    \8054 [997] = 1'h0;
    \8054 [998] = 1'h0;
    \8054 [999] = 1'h0;
    \8054 [1000] = 1'h0;
    \8054 [1001] = 1'h0;
    \8054 [1002] = 1'h0;
    \8054 [1003] = 1'h0;
    \8054 [1004] = 1'h0;
    \8054 [1005] = 1'h0;
    \8054 [1006] = 1'h0;
    \8054 [1007] = 1'h0;
    \8054 [1008] = 1'h0;
    \8054 [1009] = 1'h0;
    \8054 [1010] = 1'h0;
    \8054 [1011] = 1'h0;
    \8054 [1012] = 1'h0;
    \8054 [1013] = 1'h0;
    \8054 [1014] = 1'h0;
    \8054 [1015] = 1'h0;
    \8054 [1016] = 1'h0;
    \8054 [1017] = 1'h0;
    \8054 [1018] = 1'h0;
    \8054 [1019] = 1'h0;
    \8054 [1020] = 1'h0;
    \8054 [1021] = 1'h0;
    \8054 [1022] = 1'h0;
    \8054 [1023] = 1'h1;
  end
  assign _197_ = \8054 [_111_];
  reg [43:0] \8056  [7:0];
  initial begin
    \8056 [0] = 44'h200000000f1;
    \8056 [1] = 44'h00000000000;
    \8056 [2] = 44'h0000000e779;
    \8056 [3] = 44'h1000058e639;
    \8056 [4] = 44'h00000000000;
    \8056 [5] = 44'h00000000000;
    \8056 [6] = 44'h00000088811;
    \8056 [7] = 44'h00000c00071;
  end
  assign _199_ = \8056 [_113_];
  reg [43:0] \8058  [15:0];
  initial begin
    \8058 [0] = 44'h00000000000;
    \8058 [1] = 44'h00000000000;
    \8058 [2] = 44'h00000000000;
    \8058 [3] = 44'h00000000000;
    \8058 [4] = 44'h00000000000;
    \8058 [5] = 44'h00000000000;
    \8058 [6] = 44'h08000111191;
    \8058 [7] = 44'h08000111189;
    \8058 [8] = 44'h0800011c381;
    \8058 [9] = 44'h0800011c381;
    \8058 [10] = 44'h0800011c181;
    \8058 [11] = 44'h0800011c181;
    \8058 [12] = 44'h0800011c191;
    \8058 [13] = 44'h0800011c191;
    \8058 [14] = 44'h0800011c189;
    \8058 [15] = 44'h0800011c189;
  end
  assign _201_ = \8058 [_133_];
  reg [43:0] \8060  [3:0];
  initial begin
    \8060 [0] = 44'h00000000000;
    \8060 [1] = 44'h002600894fa;
    \8060 [2] = 44'hc04800894fa;
    \8060 [3] = 44'h000800894fa;
  end
  assign _203_ = \8060 [_138_];
  reg [43:0] \8062  [31:0];
  initial begin
    \8062 [0] = 44'h0900023facf;
    \8062 [1] = 44'h0900023facf;
    \8062 [2] = 44'h0900023facf;
    \8062 [3] = 44'h0900023facf;
    \8062 [4] = 44'h00000000000;
    \8062 [5] = 44'h0900020f0cf;
    \8062 [6] = 44'h09000230acf;
    \8062 [7] = 44'h0900020f0cf;
    \8062 [8] = 44'h00000000000;
    \8062 [9] = 44'h0900020f0cf;
    \8062 [10] = 44'h0900020facf;
    \8062 [11] = 44'h0900020facf;
    \8062 [12] = 44'h00000000000;
    \8062 [13] = 44'h0900020facf;
    \8062 [14] = 44'h00000000000;
    \8062 [15] = 44'h00000000000;
    \8062 [16] = 44'h00000000000;
    \8062 [17] = 44'h0900020f0d7;
    \8062 [18] = 44'h00000000000;
    \8062 [19] = 44'h00000000000;
    \8062 [20] = 44'h00000000000;
    \8062 [21] = 44'h00000000000;
    \8062 [22] = 44'h00000000000;
    \8062 [23] = 44'h00000000000;
    \8062 [24] = 44'h00000000000;
    \8062 [25] = 44'h00000000000;
    \8062 [26] = 44'h00000000000;
    \8062 [27] = 44'h00000000000;
    \8062 [28] = 44'h00000000000;
    \8062 [29] = 44'h00000000000;
    \8062 [30] = 44'h00000000000;
    \8062 [31] = 44'h00000000000;
  end
  assign _205_ = \8062 [_140_];
  reg [43:0] \8064  [3:0];
  initial begin
    \8064 [0] = 44'h00000000000;
    \8064 [1] = 44'h40080019502;
    \8064 [2] = 44'h00480119502;
    \8064 [3] = 44'h00080019502;
  end
  assign _207_ = \8064 [_148_];
  reg [43:0] \8066  [511:0];
  initial begin
    \8066 [0] = 44'h00000000000;
    \8066 [1] = 44'h00000000000;
    \8066 [2] = 44'h0800020f0cf;
    \8066 [3] = 44'h00000000000;
    \8066 [4] = 44'h00000000000;
    \8066 [5] = 44'h00000000000;
    \8066 [6] = 44'h0800020f0cf;
    \8066 [7] = 44'h00000000000;
    \8066 [8] = 44'h00000000000;
    \8066 [9] = 44'h00000000000;
    \8066 [10] = 44'h00000000000;
    \8066 [11] = 44'h00000000000;
    \8066 [12] = 44'h00000000000;
    \8066 [13] = 44'h00000000000;
    \8066 [14] = 44'h00000000000;
    \8066 [15] = 44'h00000000000;
    \8066 [16] = 44'h00000000000;
    \8066 [17] = 44'h00000000000;
    \8066 [18] = 44'h00000000000;
    \8066 [19] = 44'h00000000000;
    \8066 [20] = 44'h00000000000;
    \8066 [21] = 44'h00000000000;
    \8066 [22] = 44'h00000000000;
    \8066 [23] = 44'h00000000000;
    \8066 [24] = 44'h00000000000;
    \8066 [25] = 44'h00000000000;
    \8066 [26] = 44'h00000000000;
    \8066 [27] = 44'h0800020f0cf;
    \8066 [28] = 44'h00000000000;
    \8066 [29] = 44'h00000000000;
    \8066 [30] = 44'h00000000000;
    \8066 [31] = 44'h0800020f0cf;
    \8066 [32] = 44'h00000000000;
    \8066 [33] = 44'h0800020f0d7;
    \8066 [34] = 44'h0800020f0cf;
    \8066 [35] = 44'h00000000000;
    \8066 [36] = 44'h00000000000;
    \8066 [37] = 44'h0800020f0d7;
    \8066 [38] = 44'h0800020f0cf;
    \8066 [39] = 44'h00000000000;
    \8066 [40] = 44'h00000000000;
    \8066 [41] = 44'h00000000000;
    \8066 [42] = 44'h00000000000;
    \8066 [43] = 44'h00000000000;
    \8066 [44] = 44'h00000000000;
    \8066 [45] = 44'h00000000000;
    \8066 [46] = 44'h00000000000;
    \8066 [47] = 44'h00000000000;
    \8066 [48] = 44'h00000000000;
    \8066 [49] = 44'h00000000000;
    \8066 [50] = 44'h00000000000;
    \8066 [51] = 44'h00000000000;
    \8066 [52] = 44'h00000000000;
    \8066 [53] = 44'h00000000000;
    \8066 [54] = 44'h00000000000;
    \8066 [55] = 44'h00000000000;
    \8066 [56] = 44'h00000000000;
    \8066 [57] = 44'h00000000000;
    \8066 [58] = 44'h00000000000;
    \8066 [59] = 44'h0800020f0cf;
    \8066 [60] = 44'h00000000000;
    \8066 [61] = 44'h00000000000;
    \8066 [62] = 44'h00000000000;
    \8066 [63] = 44'h0800020f0cf;
    \8066 [64] = 44'h00000000000;
    \8066 [65] = 44'h00000000000;
    \8066 [66] = 44'h00000000000;
    \8066 [67] = 44'h00000000000;
    \8066 [68] = 44'h00000000000;
    \8066 [69] = 44'h00000000000;
    \8066 [70] = 44'h00000000000;
    \8066 [71] = 44'h00000000000;
    \8066 [72] = 44'h00000000000;
    \8066 [73] = 44'h00000000000;
    \8066 [74] = 44'h00000000000;
    \8066 [75] = 44'h00000000000;
    \8066 [76] = 44'h00000000000;
    \8066 [77] = 44'h00000000000;
    \8066 [78] = 44'h00000000000;
    \8066 [79] = 44'h00000000000;
    \8066 [80] = 44'h00000000000;
    \8066 [81] = 44'h00000000000;
    \8066 [82] = 44'h00000000000;
    \8066 [83] = 44'h00000000000;
    \8066 [84] = 44'h00000000000;
    \8066 [85] = 44'h00000000000;
    \8066 [86] = 44'h00000000000;
    \8066 [87] = 44'h00000000000;
    \8066 [88] = 44'h00000000000;
    \8066 [89] = 44'h00000000000;
    \8066 [90] = 44'h00000000000;
    \8066 [91] = 44'h00000000000;
    \8066 [92] = 44'h00000000000;
    \8066 [93] = 44'h00000000000;
    \8066 [94] = 44'h00000000000;
    \8066 [95] = 44'h00000000000;
    \8066 [96] = 44'h00000000000;
    \8066 [97] = 44'h00000000000;
    \8066 [98] = 44'h00000000000;
    \8066 [99] = 44'h00000000000;
    \8066 [100] = 44'h00000000000;
    \8066 [101] = 44'h00000000000;
    \8066 [102] = 44'h00000000000;
    \8066 [103] = 44'h00000000000;
    \8066 [104] = 44'h00000000000;
    \8066 [105] = 44'h00000000000;
    \8066 [106] = 44'h00000000000;
    \8066 [107] = 44'h00000000000;
    \8066 [108] = 44'h00000000000;
    \8066 [109] = 44'h00000000000;
    \8066 [110] = 44'h00000000000;
    \8066 [111] = 44'h00000000000;
    \8066 [112] = 44'h00000000000;
    \8066 [113] = 44'h00000000000;
    \8066 [114] = 44'h00000000000;
    \8066 [115] = 44'h00000000000;
    \8066 [116] = 44'h00000000000;
    \8066 [117] = 44'h00000000000;
    \8066 [118] = 44'h00000000000;
    \8066 [119] = 44'h00000000000;
    \8066 [120] = 44'h00000000000;
    \8066 [121] = 44'h00000000000;
    \8066 [122] = 44'h00000000000;
    \8066 [123] = 44'h00000000000;
    \8066 [124] = 44'h00000000000;
    \8066 [125] = 44'h00000000000;
    \8066 [126] = 44'h00000000000;
    \8066 [127] = 44'h0900020f0cf;
    \8066 [128] = 44'h00000000000;
    \8066 [129] = 44'h00000000000;
    \8066 [130] = 44'h00000000000;
    \8066 [131] = 44'h00000000000;
    \8066 [132] = 44'h00000000000;
    \8066 [133] = 44'h00000000000;
    \8066 [134] = 44'h00000000000;
    \8066 [135] = 44'h00000000000;
    \8066 [136] = 44'h00000000000;
    \8066 [137] = 44'h00000000000;
    \8066 [138] = 44'h00000000000;
    \8066 [139] = 44'h00000000000;
    \8066 [140] = 44'h00000000000;
    \8066 [141] = 44'h00000000000;
    \8066 [142] = 44'h00000000000;
    \8066 [143] = 44'h00000000000;
    \8066 [144] = 44'h00000000000;
    \8066 [145] = 44'h00000000000;
    \8066 [146] = 44'h00000000000;
    \8066 [147] = 44'h00000000000;
    \8066 [148] = 44'h00000000000;
    \8066 [149] = 44'h00000000000;
    \8066 [150] = 44'h00000000000;
    \8066 [151] = 44'h00000000000;
    \8066 [152] = 44'h00000000000;
    \8066 [153] = 44'h00000000000;
    \8066 [154] = 44'h00000000000;
    \8066 [155] = 44'h00000000000;
    \8066 [156] = 44'h00000000000;
    \8066 [157] = 44'h00000000000;
    \8066 [158] = 44'h00000000000;
    \8066 [159] = 44'h00000000000;
    \8066 [160] = 44'h00000000000;
    \8066 [161] = 44'h00000000000;
    \8066 [162] = 44'h00000000000;
    \8066 [163] = 44'h00000000000;
    \8066 [164] = 44'h00000000000;
    \8066 [165] = 44'h00000000000;
    \8066 [166] = 44'h00000000000;
    \8066 [167] = 44'h00000000000;
    \8066 [168] = 44'h00000000000;
    \8066 [169] = 44'h00000000000;
    \8066 [170] = 44'h00000000000;
    \8066 [171] = 44'h00000000000;
    \8066 [172] = 44'h00000000000;
    \8066 [173] = 44'h00000000000;
    \8066 [174] = 44'h00000000000;
    \8066 [175] = 44'h00000000000;
    \8066 [176] = 44'h00000000000;
    \8066 [177] = 44'h00000000000;
    \8066 [178] = 44'h00000000000;
    \8066 [179] = 44'h00000000000;
    \8066 [180] = 44'h00000000000;
    \8066 [181] = 44'h00000000000;
    \8066 [182] = 44'h00000000000;
    \8066 [183] = 44'h00000000000;
    \8066 [184] = 44'h00000000000;
    \8066 [185] = 44'h00000000000;
    \8066 [186] = 44'h00000000000;
    \8066 [187] = 44'h00000000000;
    \8066 [188] = 44'h00000000000;
    \8066 [189] = 44'h00000000000;
    \8066 [190] = 44'h00000000000;
    \8066 [191] = 44'h00000000000;
    \8066 [192] = 44'h00000000000;
    \8066 [193] = 44'h00000000000;
    \8066 [194] = 44'h00000000000;
    \8066 [195] = 44'h00000000000;
    \8066 [196] = 44'h00000000000;
    \8066 [197] = 44'h00000000000;
    \8066 [198] = 44'h00000000000;
    \8066 [199] = 44'h00000000000;
    \8066 [200] = 44'h00000000000;
    \8066 [201] = 44'h00000000000;
    \8066 [202] = 44'h00000000000;
    \8066 [203] = 44'h00000000000;
    \8066 [204] = 44'h00000000000;
    \8066 [205] = 44'h00000000000;
    \8066 [206] = 44'h00000000000;
    \8066 [207] = 44'h00000000000;
    \8066 [208] = 44'h00000000000;
    \8066 [209] = 44'h00000000000;
    \8066 [210] = 44'h00000000000;
    \8066 [211] = 44'h00000000000;
    \8066 [212] = 44'h00000000000;
    \8066 [213] = 44'h00000000000;
    \8066 [214] = 44'h00000000000;
    \8066 [215] = 44'h00000000000;
    \8066 [216] = 44'h00000000000;
    \8066 [217] = 44'h00000000000;
    \8066 [218] = 44'h00000000000;
    \8066 [219] = 44'h00000000000;
    \8066 [220] = 44'h00000000000;
    \8066 [221] = 44'h00000000000;
    \8066 [222] = 44'h00000000000;
    \8066 [223] = 44'h00000000000;
    \8066 [224] = 44'h00000000000;
    \8066 [225] = 44'h00000000000;
    \8066 [226] = 44'h00000000000;
    \8066 [227] = 44'h00000000000;
    \8066 [228] = 44'h00000000000;
    \8066 [229] = 44'h00000000000;
    \8066 [230] = 44'h00000000000;
    \8066 [231] = 44'h00000000000;
    \8066 [232] = 44'h00000000000;
    \8066 [233] = 44'h00000000000;
    \8066 [234] = 44'h00000000000;
    \8066 [235] = 44'h00000000000;
    \8066 [236] = 44'h00000000000;
    \8066 [237] = 44'h00000000000;
    \8066 [238] = 44'h00000000000;
    \8066 [239] = 44'h00000000000;
    \8066 [240] = 44'h0800020f0cf;
    \8066 [241] = 44'h0800020f0cf;
    \8066 [242] = 44'h0800020f0cf;
    \8066 [243] = 44'h0800020f0cf;
    \8066 [244] = 44'h00000000000;
    \8066 [245] = 44'h00000000000;
    \8066 [246] = 44'h00000000000;
    \8066 [247] = 44'h0800020f0cf;
    \8066 [248] = 44'h00000000000;
    \8066 [249] = 44'h00000000000;
    \8066 [250] = 44'h00000000000;
    \8066 [251] = 44'h0800020f0cf;
    \8066 [252] = 44'h00000000000;
    \8066 [253] = 44'h0800020f0cf;
    \8066 [254] = 44'h0800020f0cf;
    \8066 [255] = 44'h0800020facf;
    \8066 [256] = 44'h00000000000;
    \8066 [257] = 44'h00000000000;
    \8066 [258] = 44'h00000000000;
    \8066 [259] = 44'h00000000000;
    \8066 [260] = 44'h00000000000;
    \8066 [261] = 44'h00000000000;
    \8066 [262] = 44'h00000000000;
    \8066 [263] = 44'h00000000000;
    \8066 [264] = 44'h00000000000;
    \8066 [265] = 44'h0800000f0d7;
    \8066 [266] = 44'h00000000000;
    \8066 [267] = 44'h00000000000;
    \8066 [268] = 44'h00000000000;
    \8066 [269] = 44'h0800020f0d7;
    \8066 [270] = 44'h00000000000;
    \8066 [271] = 44'h00000000000;
    \8066 [272] = 44'h00000000000;
    \8066 [273] = 44'h00000000000;
    \8066 [274] = 44'h00000000000;
    \8066 [275] = 44'h00000000000;
    \8066 [276] = 44'h00000000000;
    \8066 [277] = 44'h00000000000;
    \8066 [278] = 44'h00000000000;
    \8066 [279] = 44'h00000000000;
    \8066 [280] = 44'h00000000000;
    \8066 [281] = 44'h00000000000;
    \8066 [282] = 44'h00000000000;
    \8066 [283] = 44'h00000000000;
    \8066 [284] = 44'h00000000000;
    \8066 [285] = 44'h00000000000;
    \8066 [286] = 44'h00000000000;
    \8066 [287] = 44'h00000000000;
    \8066 [288] = 44'h00000000000;
    \8066 [289] = 44'h0000020fad7;
    \8066 [290] = 44'h00000000000;
    \8066 [291] = 44'h00000000000;
    \8066 [292] = 44'h00000000000;
    \8066 [293] = 44'h0000020fad7;
    \8066 [294] = 44'h00000000000;
    \8066 [295] = 44'h00000000000;
    \8066 [296] = 44'h00000000000;
    \8066 [297] = 44'h00000000000;
    \8066 [298] = 44'h00000000000;
    \8066 [299] = 44'h00000000000;
    \8066 [300] = 44'h00000000000;
    \8066 [301] = 44'h00000000000;
    \8066 [302] = 44'h00000000000;
    \8066 [303] = 44'h00000000000;
    \8066 [304] = 44'h00000000000;
    \8066 [305] = 44'h00000000000;
    \8066 [306] = 44'h00000000000;
    \8066 [307] = 44'h00000000000;
    \8066 [308] = 44'h00000000000;
    \8066 [309] = 44'h00000000000;
    \8066 [310] = 44'h00000000000;
    \8066 [311] = 44'h00000000000;
    \8066 [312] = 44'h00000000000;
    \8066 [313] = 44'h00000000000;
    \8066 [314] = 44'h00000000000;
    \8066 [315] = 44'h080000000cf;
    \8066 [316] = 44'h00000000000;
    \8066 [317] = 44'h080000000cf;
    \8066 [318] = 44'h080000000cf;
    \8066 [319] = 44'h00000000000;
    \8066 [320] = 44'h00000000000;
    \8066 [321] = 44'h00000000000;
    \8066 [322] = 44'h00000000000;
    \8066 [323] = 44'h00000000000;
    \8066 [324] = 44'h00000000000;
    \8066 [325] = 44'h00000000000;
    \8066 [326] = 44'h00000000000;
    \8066 [327] = 44'h00000000000;
    \8066 [328] = 44'h00000000000;
    \8066 [329] = 44'h00000000000;
    \8066 [330] = 44'h00000000000;
    \8066 [331] = 44'h00000000000;
    \8066 [332] = 44'h00000000000;
    \8066 [333] = 44'h00000000000;
    \8066 [334] = 44'h00000000000;
    \8066 [335] = 44'h00000000000;
    \8066 [336] = 44'h00000000000;
    \8066 [337] = 44'h00000000000;
    \8066 [338] = 44'h00000000000;
    \8066 [339] = 44'h00000000000;
    \8066 [340] = 44'h00000000000;
    \8066 [341] = 44'h00000000000;
    \8066 [342] = 44'h00000000000;
    \8066 [343] = 44'h00000000000;
    \8066 [344] = 44'h00000000000;
    \8066 [345] = 44'h00000000000;
    \8066 [346] = 44'h00000000000;
    \8066 [347] = 44'h00000000000;
    \8066 [348] = 44'h00000000000;
    \8066 [349] = 44'h00000000000;
    \8066 [350] = 44'h00000000000;
    \8066 [351] = 44'h00000000000;
    \8066 [352] = 44'h00000000000;
    \8066 [353] = 44'h00000000000;
    \8066 [354] = 44'h00000000000;
    \8066 [355] = 44'h00000000000;
    \8066 [356] = 44'h00000000000;
    \8066 [357] = 44'h00000000000;
    \8066 [358] = 44'h00000000000;
    \8066 [359] = 44'h00000000000;
    \8066 [360] = 44'h00000000000;
    \8066 [361] = 44'h00000000000;
    \8066 [362] = 44'h00000000000;
    \8066 [363] = 44'h00000000000;
    \8066 [364] = 44'h00000000000;
    \8066 [365] = 44'h00000000000;
    \8066 [366] = 44'h00000000000;
    \8066 [367] = 44'h00000000000;
    \8066 [368] = 44'h00000000000;
    \8066 [369] = 44'h00000000000;
    \8066 [370] = 44'h00000000000;
    \8066 [371] = 44'h00000000000;
    \8066 [372] = 44'h00000000000;
    \8066 [373] = 44'h00000000000;
    \8066 [374] = 44'h00000000000;
    \8066 [375] = 44'h00000000000;
    \8066 [376] = 44'h00000000000;
    \8066 [377] = 44'h00000000000;
    \8066 [378] = 44'h00000000000;
    \8066 [379] = 44'h00000000000;
    \8066 [380] = 44'h00000000000;
    \8066 [381] = 44'h00000000000;
    \8066 [382] = 44'h00000000000;
    \8066 [383] = 44'h00000000000;
    \8066 [384] = 44'h00000000000;
    \8066 [385] = 44'h00000000000;
    \8066 [386] = 44'h00000000000;
    \8066 [387] = 44'h00000000000;
    \8066 [388] = 44'h00000000000;
    \8066 [389] = 44'h00000000000;
    \8066 [390] = 44'h00000000000;
    \8066 [391] = 44'h00000000000;
    \8066 [392] = 44'h00000000000;
    \8066 [393] = 44'h00000000000;
    \8066 [394] = 44'h00000000000;
    \8066 [395] = 44'h00000000000;
    \8066 [396] = 44'h00000000000;
    \8066 [397] = 44'h00000000000;
    \8066 [398] = 44'h00000000000;
    \8066 [399] = 44'h00000000000;
    \8066 [400] = 44'h00000000000;
    \8066 [401] = 44'h00000000000;
    \8066 [402] = 44'h00000000000;
    \8066 [403] = 44'h00000000000;
    \8066 [404] = 44'h00000000000;
    \8066 [405] = 44'h00000000000;
    \8066 [406] = 44'h00000000000;
    \8066 [407] = 44'h00000000000;
    \8066 [408] = 44'h00000000000;
    \8066 [409] = 44'h00000000000;
    \8066 [410] = 44'h00000000000;
    \8066 [411] = 44'h00000000000;
    \8066 [412] = 44'h00000000000;
    \8066 [413] = 44'h00000000000;
    \8066 [414] = 44'h00000000000;
    \8066 [415] = 44'h00000000000;
    \8066 [416] = 44'h00000000000;
    \8066 [417] = 44'h00000000000;
    \8066 [418] = 44'h00000000000;
    \8066 [419] = 44'h00000000000;
    \8066 [420] = 44'h00000000000;
    \8066 [421] = 44'h00000000000;
    \8066 [422] = 44'h00000000000;
    \8066 [423] = 44'h00000000000;
    \8066 [424] = 44'h00000000000;
    \8066 [425] = 44'h00000000000;
    \8066 [426] = 44'h00000000000;
    \8066 [427] = 44'h00000000000;
    \8066 [428] = 44'h00000000000;
    \8066 [429] = 44'h00000000000;
    \8066 [430] = 44'h00000000000;
    \8066 [431] = 44'h00000000000;
    \8066 [432] = 44'h00000000000;
    \8066 [433] = 44'h00000000000;
    \8066 [434] = 44'h00000000000;
    \8066 [435] = 44'h00000000000;
    \8066 [436] = 44'h00000000000;
    \8066 [437] = 44'h00000000000;
    \8066 [438] = 44'h00000000000;
    \8066 [439] = 44'h00000000000;
    \8066 [440] = 44'h00000000000;
    \8066 [441] = 44'h00000000000;
    \8066 [442] = 44'h00000000000;
    \8066 [443] = 44'h00000000000;
    \8066 [444] = 44'h00000000000;
    \8066 [445] = 44'h00000000000;
    \8066 [446] = 44'h00000000000;
    \8066 [447] = 44'h00000000000;
    \8066 [448] = 44'h00000000000;
    \8066 [449] = 44'h00000000000;
    \8066 [450] = 44'h00000000000;
    \8066 [451] = 44'h00000000000;
    \8066 [452] = 44'h00000000000;
    \8066 [453] = 44'h00000000000;
    \8066 [454] = 44'h00000000000;
    \8066 [455] = 44'h00000000000;
    \8066 [456] = 44'h00000000000;
    \8066 [457] = 44'h00000000000;
    \8066 [458] = 44'h00000000000;
    \8066 [459] = 44'h00000000000;
    \8066 [460] = 44'h00000000000;
    \8066 [461] = 44'h00000000000;
    \8066 [462] = 44'h00000000000;
    \8066 [463] = 44'h00000000000;
    \8066 [464] = 44'h00000000000;
    \8066 [465] = 44'h00000000000;
    \8066 [466] = 44'h00000000000;
    \8066 [467] = 44'h00000000000;
    \8066 [468] = 44'h00000000000;
    \8066 [469] = 44'h00000000000;
    \8066 [470] = 44'h00000000000;
    \8066 [471] = 44'h00000000000;
    \8066 [472] = 44'h00000000000;
    \8066 [473] = 44'h00000000000;
    \8066 [474] = 44'h00000000000;
    \8066 [475] = 44'h00000000000;
    \8066 [476] = 44'h00000000000;
    \8066 [477] = 44'h00000000000;
    \8066 [478] = 44'h00000000000;
    \8066 [479] = 44'h00000000000;
    \8066 [480] = 44'h00000000000;
    \8066 [481] = 44'h00000000000;
    \8066 [482] = 44'h00000000000;
    \8066 [483] = 44'h00000000000;
    \8066 [484] = 44'h00000000000;
    \8066 [485] = 44'h00000000000;
    \8066 [486] = 44'h00000000000;
    \8066 [487] = 44'h00000000000;
    \8066 [488] = 44'h00000000000;
    \8066 [489] = 44'h00000000000;
    \8066 [490] = 44'h00000000000;
    \8066 [491] = 44'h00000000000;
    \8066 [492] = 44'h00000000000;
    \8066 [493] = 44'h00000000000;
    \8066 [494] = 44'h00000000000;
    \8066 [495] = 44'h00000000000;
    \8066 [496] = 44'h00000000000;
    \8066 [497] = 44'h00000000000;
    \8066 [498] = 44'h00000000000;
    \8066 [499] = 44'h00000000000;
    \8066 [500] = 44'h00000000000;
    \8066 [501] = 44'h00000000000;
    \8066 [502] = 44'h00000000000;
    \8066 [503] = 44'h00000000000;
    \8066 [504] = 44'h00000000000;
    \8066 [505] = 44'h00000000000;
    \8066 [506] = 44'h0000080f0cf;
    \8066 [507] = 44'h0000080facf;
    \8066 [508] = 44'h00000000000;
    \8066 [509] = 44'h000008000cf;
    \8066 [510] = 44'h0000080facf;
    \8066 [511] = 44'h0000080facf;
  end
  assign _209_ = \8066 [_151_];
  reg [43:0] \8068  [16:0];
  initial begin
    \8068 [0] = 44'h00000000000;
    \8068 [1] = 44'h0800023facf;
    \8068 [2] = 44'h0800023facf;
    \8068 [3] = 44'h0800023facf;
    \8068 [4] = 44'h0800023facf;
    \8068 [5] = 44'h00000000000;
    \8068 [6] = 44'h0800020f0cf;
    \8068 [7] = 44'h08000230acf;
    \8068 [8] = 44'h0800020f0cf;
    \8068 [9] = 44'h0800023facf;
    \8068 [10] = 44'h0800020f0cf;
    \8068 [11] = 44'h0800020facf;
    \8068 [12] = 44'h0800020facf;
    \8068 [13] = 44'h00000000000;
    \8068 [14] = 44'h0800020facf;
    \8068 [15] = 44'h00000000000;
    \8068 [16] = 44'h00000000000;
  end
  assign _211_ = \8068 [_152_];
  assign _000_ = ~ stall_in;
  assign _001_ = _000_ ? s : r;
  assign _002_ = _000_ ? 1'h0 : s[0];
  assign _003_ = _000_ ? si : ri;
  assign _004_ = rin[0] & r[0];
  assign _005_ = _004_ & stall_in;
  assign _006_ = ~ r[0];
  assign _007_ = ~ stall_in;
  assign _008_ = _006_ | _007_;
  assign _009_ = _008_ ? rin : r;
  assign _010_ = _008_ ? ri_in : ri;
  assign _011_ = s[0] ? _001_ : _009_;
  assign _012_ = s[0] ? _002_ : _005_;
  assign _013_ = s[0] ? s[164:1] : rin[164:1];
  assign _014_ = s[0] ? _003_ : _010_;
  assign _015_ = s[0] ? si : ri_in;
  assign _016_ = flush_in ? 1'h0 : _011_[0];
  assign _017_ = flush_in ? r[164:1] : _011_[164:1];
  assign _018_ = flush_in ? 1'h0 : _012_;
  assign _019_ = flush_in ? s[164:1] : _013_;
  assign _020_ = flush_in ? ri : _014_;
  assign _021_ = flush_in ? si : _015_;
  assign _022_ = rst ? 165'h000000000000000000000000000000000000000000 : { _017_, _016_ };
  assign _023_ = rst ? 165'h000000000000000000000000000000000000000000 : { _019_, _018_ };
  assign _024_ = rst ? 47'h000000000000 : _020_;
  assign _025_ = rst ? 47'h000000000000 : _021_;
  assign _026_ = rst ? 87'h0000000000000000000000 : br_in;
  always @(posedge clk)
    _027_ <= _022_;
  always @(posedge clk)
    _028_ <= _023_;
  always @(posedge clk)
    _029_ <= _024_;
  always @(posedge clk)
    _030_ <= _025_;
  always @(posedge clk)
    _031_ <= _026_;
  assign _032_ = 6'h3f - \f_in.insn [31:26];
  assign _033_ = 11'h7ff - { \f_in.insn [5:0], \f_in.insn [10:6] };
  assign _034_ = ~ _191_;
  assign _035_ = 6'h3f - \f_in.insn [5:0];
  assign _036_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h00000004;
  assign _037_ = 10'h3ff - \f_in.insn [10:1];
  assign _038_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h008;
  assign _039_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h009;
  assign _040_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h01a;
  assign _041_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h01b;
  assign _042_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h13a;
  assign _043_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h13b;
  assign _044_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h110;
  assign _045_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h111;
  assign _046_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h112;
  assign _047_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h113;
  assign _048_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h103;
  assign _049_ = _047_ | _048_;
  assign _050_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h130;
  assign _051_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h131;
  assign _052_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h001;
  assign _053_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h32f;
  function [0:0] \7567 ;
    input [0:0] a;
    input [13:0] b;
    input [13:0] s;
    (* parallel_case *)
    casez (s)
      14'b?????????????1:
        \7567  = b[0:0];
      14'b????????????1?:
        \7567  = b[1:1];
      14'b???????????1??:
        \7567  = b[2:2];
      14'b??????????1???:
        \7567  = b[3:3];
      14'b?????????1????:
        \7567  = b[4:4];
      14'b????????1?????:
        \7567  = b[5:5];
      14'b???????1??????:
        \7567  = b[6:6];
      14'b??????1???????:
        \7567  = b[7:7];
      14'b?????1????????:
        \7567  = b[8:8];
      14'b????1?????????:
        \7567  = b[9:9];
      14'b???1??????????:
        \7567  = b[10:10];
      14'b??1???????????:
        \7567  = b[11:11];
      14'b?1????????????:
        \7567  = b[12:12];
      14'b1?????????????:
        \7567  = b[13:13];
      default:
        \7567  = a;
    endcase
  endfunction
  assign _054_ = \7567 (1'h0, 14'h3fff, { _053_, _052_, _051_, _050_, _049_, _046_, _045_, _044_, _043_, _042_, _041_, _040_, _039_, _038_ });
  function [6:0] \7573 ;
    input [6:0] a;
    input [97:0] b;
    input [13:0] s;
    (* parallel_case *)
    casez (s)
      14'b?????????????1:
        \7573  = b[6:0];
      14'b????????????1?:
        \7573  = b[13:7];
      14'b???????????1??:
        \7573  = b[20:14];
      14'b??????????1???:
        \7573  = b[27:21];
      14'b?????????1????:
        \7573  = b[34:28];
      14'b????????1?????:
        \7573  = b[41:35];
      14'b???????1??????:
        \7573  = b[48:42];
      14'b??????1???????:
        \7573  = b[55:49];
      14'b?????1????????:
        \7573  = b[62:56];
      14'b????1?????????:
        \7573  = b[69:63];
      14'b???1??????????:
        \7573  = b[76:70];
      14'b??1???????????:
        \7573  = b[83:77];
      14'b?1????????????:
        \7573  = b[90:84];
      14'b1?????????????:
        \7573  = b[97:91];
      default:
        \7573  = a;
    endcase
  endfunction
  assign _055_ = \7573 (7'h00, 98'hxxxxxxxxxxxxxxxxxxxxxxxxx, { _053_, _052_, _051_, _050_, _049_, _046_, _045_, _044_, _043_, _042_, _041_, _040_, _039_, _038_ });
  function [4:0] \7589 ;
    input [4:0] a;
    input [69:0] b;
    input [13:0] s;
    (* parallel_case *)
    casez (s)
      14'b?????????????1:
        \7589  = b[4:0];
      14'b????????????1?:
        \7589  = b[9:5];
      14'b???????????1??:
        \7589  = b[14:10];
      14'b??????????1???:
        \7589  = b[19:15];
      14'b?????????1????:
        \7589  = b[24:20];
      14'b????????1?????:
        \7589  = b[29:25];
      14'b???????1??????:
        \7589  = b[34:30];
      14'b??????1???????:
        \7589  = b[39:35];
      14'b?????1????????:
        \7589  = b[44:40];
      14'b????1?????????:
        \7589  = b[49:45];
      14'b???1??????????:
        \7589  = b[54:50];
      14'b??1???????????:
        \7589  = b[59:55];
      14'b?1????????????:
        \7589  = b[64:60];
      14'b1?????????????:
        \7589  = b[69:65];
      default:
        \7589  = a;
    endcase
  endfunction
  assign _056_ = \7589 (5'h00, 70'h1ac5a928398a418820, { _053_, _052_, _051_, _050_, _049_, _046_, _045_, _044_, _043_, _042_, _041_, _040_, _039_, _038_ });
  assign _057_ = _054_ ? _056_ : 5'hxx;
  assign _058_ = _054_ ? { 2'h1, _057_ } : _055_;
  assign _059_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h008;
  assign _060_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h009;
  assign _061_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h01a;
  assign _062_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h01b;
  assign _063_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h13a;
  assign _064_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h13b;
  assign _065_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h110;
  assign _066_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h111;
  assign _067_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h112;
  assign _068_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h113;
  assign _069_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h103;
  assign _070_ = _068_ | _069_;
  assign _071_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h130;
  assign _072_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h131;
  assign _073_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h001;
  assign _074_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h32f;
  function [0:0] \7644 ;
    input [0:0] a;
    input [13:0] b;
    input [13:0] s;
    (* parallel_case *)
    casez (s)
      14'b?????????????1:
        \7644  = b[0:0];
      14'b????????????1?:
        \7644  = b[1:1];
      14'b???????????1??:
        \7644  = b[2:2];
      14'b??????????1???:
        \7644  = b[3:3];
      14'b?????????1????:
        \7644  = b[4:4];
      14'b????????1?????:
        \7644  = b[5:5];
      14'b???????1??????:
        \7644  = b[6:6];
      14'b??????1???????:
        \7644  = b[7:7];
      14'b?????1????????:
        \7644  = b[8:8];
      14'b????1?????????:
        \7644  = b[9:9];
      14'b???1??????????:
        \7644  = b[10:10];
      14'b??1???????????:
        \7644  = b[11:11];
      14'b?1????????????:
        \7644  = b[12:12];
      14'b1?????????????:
        \7644  = b[13:13];
      default:
        \7644  = a;
    endcase
  endfunction
  assign _075_ = \7644 (1'h0, 14'h3fff, { _074_, _073_, _072_, _071_, _070_, _067_, _066_, _065_, _064_, _063_, _062_, _061_, _060_, _059_ });
  function [6:0] \7650 ;
    input [6:0] a;
    input [97:0] b;
    input [13:0] s;
    (* parallel_case *)
    casez (s)
      14'b?????????????1:
        \7650  = b[6:0];
      14'b????????????1?:
        \7650  = b[13:7];
      14'b???????????1??:
        \7650  = b[20:14];
      14'b??????????1???:
        \7650  = b[27:21];
      14'b?????????1????:
        \7650  = b[34:28];
      14'b????????1?????:
        \7650  = b[41:35];
      14'b???????1??????:
        \7650  = b[48:42];
      14'b??????1???????:
        \7650  = b[55:49];
      14'b?????1????????:
        \7650  = b[62:56];
      14'b????1?????????:
        \7650  = b[69:63];
      14'b???1??????????:
        \7650  = b[76:70];
      14'b??1???????????:
        \7650  = b[83:77];
      14'b?1????????????:
        \7650  = b[90:84];
      14'b1?????????????:
        \7650  = b[97:91];
      default:
        \7650  = a;
    endcase
  endfunction
  assign _076_ = \7650 (7'h00, 98'hxxxxxxxxxxxxxxxxxxxxxxxxx, { _074_, _073_, _072_, _071_, _070_, _067_, _066_, _065_, _064_, _063_, _062_, _061_, _060_, _059_ });
  function [4:0] \7666 ;
    input [4:0] a;
    input [69:0] b;
    input [13:0] s;
    (* parallel_case *)
    casez (s)
      14'b?????????????1:
        \7666  = b[4:0];
      14'b????????????1?:
        \7666  = b[9:5];
      14'b???????????1??:
        \7666  = b[14:10];
      14'b??????????1???:
        \7666  = b[19:15];
      14'b?????????1????:
        \7666  = b[24:20];
      14'b????????1?????:
        \7666  = b[29:25];
      14'b???????1??????:
        \7666  = b[34:30];
      14'b??????1???????:
        \7666  = b[39:35];
      14'b?????1????????:
        \7666  = b[44:40];
      14'b????1?????????:
        \7666  = b[49:45];
      14'b???1??????????:
        \7666  = b[54:50];
      14'b??1???????????:
        \7666  = b[59:55];
      14'b?1????????????:
        \7666  = b[64:60];
      14'b1?????????????:
        \7666  = b[69:65];
      default:
        \7666  = a;
    endcase
  endfunction
  assign _077_ = \7666 (5'h00, 70'h1ac5a928398a418820, { _074_, _073_, _072_, _071_, _070_, _067_, _066_, _065_, _064_, _063_, _062_, _061_, _060_, _059_ });
  assign _078_ = _075_ ? _077_ : 5'hxx;
  assign _079_ = _075_ ? { 2'h1, _078_ } : _076_;
  assign _080_ = \f_in.insn [10:1] & 10'h37f;
  assign _081_ = _080_ == 10'h153;
  assign _082_ = ~ _058_[5];
  assign _083_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h013;
  assign _084_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h012;
  assign _085_ = _083_ | _084_;
  assign _086_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h030;
  assign _087_ = _085_ | _086_;
  assign _088_ = { \f_in.insn [15:11], \f_in.insn [20:16] } == 10'h1d0;
  assign _089_ = _087_ | _088_;
  function [1:0] \7709 ;
    input [1:0] a;
    input [1:0] b;
    input [0:0] s;
    (* parallel_case *)
    casez (s)
      1'b1:
        \7709  = b[1:0];
      default:
        \7709  = a;
    endcase
  endfunction
  assign _090_ = \7709 (2'h0, 2'h2, _089_);
  function [0:0] \7711 ;
    input [0:0] a;
    input [0:0] b;
    input [0:0] s;
    (* parallel_case *)
    casez (s)
      1'b1:
        \7711  = b[0:0];
      default:
        \7711  = a;
    endcase
  endfunction
  assign _091_ = \7711 (1'h0, 1'h1, _089_);
  assign _092_ = _082_ ? _090_ : 2'h0;
  assign _093_ = _082_ ? { 1'h1, _091_ } : 2'h0;
  assign _094_ = _081_ ? _092_ : 2'h0;
  assign _095_ = _081_ ? _093_ : 2'h0;
  assign _096_ = \f_in.insn [10:1] & 10'h3ff;
  assign _097_ = _096_ == 10'h114;
  assign _098_ = \f_in.insn [25:21] == \f_in.insn [20:16];
  assign _099_ = \f_in.insn [25:21] == \f_in.insn [15:11];
  assign _100_ = _098_ | _099_;
  assign _101_ = _100_ ? 1'h1 : 1'h0;
  assign _102_ = _097_ ? _101_ : 1'h0;
  assign _103_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h0000001f;
  assign _104_ = ~ \f_in.insn [23];
  assign _105_ = \f_in.insn [0] ? 7'h20 : 7'h00;
  assign _106_ = _104_ ? 7'h21 : 7'h00;
  assign _107_ = _104_ ? 7'h21 : _105_;
  assign _108_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h00000010;
  assign _109_ = \f_in.insn [0] ? 7'h20 : 7'h00;
  assign _110_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h00000012;
  assign _111_ = 10'h3ff - { \f_in.insn [5:1], \f_in.insn [10:6] };
  assign _112_ = ~ _197_;
  assign _113_ = 3'h7 - { \f_in.insn [5], \f_in.insn [3:2] };
  assign _114_ = ~ \f_in.insn [2];
  assign _115_ = ~ \f_in.insn [23];
  assign _116_ = ~ \f_in.insn [10];
  assign _117_ = _116_ | \f_in.insn [6];
  assign _118_ = _115_ & _117_;
  assign _119_ = \f_in.insn [0] ? 7'h20 : 7'h00;
  assign _120_ = _118_ ? 7'h21 : 7'h00;
  assign _121_ = _118_ ? 7'h21 : _119_;
  assign _122_ = ~ \f_in.insn [10];
  assign _123_ = ~ \f_in.insn [6];
  assign _124_ = _123_ ? 7'h21 : 7'h2d;
  assign _125_ = _122_ ? 7'h20 : _124_;
  assign _126_ = _114_ ? { _125_, _120_ } : 14'h1123;
  assign _127_ = _114_ ? _121_ : 7'h00;
  assign _128_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h00000013;
  assign _129_ = \f_in.insn  & 32'd4294967295;
  assign _130_ = _129_ == 32'd1610612736;
  assign _131_ = _130_ ? 45'h000000000013 : 45'h000000000000;
  assign _132_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h00000018;
  assign _133_ = 4'hf - \f_in.insn [4:1];
  assign _134_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h0000001e;
  assign _135_ = \f_in.insn [25:21] == \f_in.insn [20:16];
  assign _136_ = _135_ ? 1'h1 : 1'h0;
  assign _137_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h00000038;
  assign _138_ = 2'h3 - \f_in.insn [1:0];
  assign _139_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h0000003a;
  assign _140_ = 5'h1f - \f_in.insn [5:1];
  assign _141_ = ~ \f_in.insn [5];
  assign _142_ = \f_in.insn [10:1] & 10'h37f;
  assign _143_ = _142_ == 10'h34e;
  assign _144_ = ~ _143_;
  assign _145_ = _141_ & _144_;
  assign _146_ = _145_ ? 1'h1 : 1'h0;
  assign _147_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h0000003b;
  assign _148_ = 2'h3 - \f_in.insn [1:0];
  assign _149_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h0000003e;
  assign _150_ = ~ \f_in.insn [5];
  assign _151_ = 9'h1ff - { \f_in.insn [4:1], \f_in.insn [10:6] };
  assign _152_ = 5'h10 - { 1'h0, \f_in.insn [4:1] };
  assign _153_ = _150_ ? _209_ : _211_;
  assign _154_ = { 25'h0000000, \f_in.insn [31:26] } == 31'h0000003f;
  function [6:0] \7928 ;
    input [6:0] a;
    input [83:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7928  = b[6:0];
      12'b??????????1?:
        \7928  = b[13:7];
      12'b?????????1??:
        \7928  = b[20:14];
      12'b????????1???:
        \7928  = b[27:21];
      12'b???????1????:
        \7928  = b[34:28];
      12'b??????1?????:
        \7928  = b[41:35];
      12'b?????1??????:
        \7928  = b[48:42];
      12'b????1???????:
        \7928  = b[55:49];
      12'b???1????????:
        \7928  = b[62:56];
      12'b??1?????????:
        \7928  = b[69:63];
      12'b?1??????????:
        \7928  = b[76:70];
      12'b1???????????:
        \7928  = b[83:77];
      default:
        \7928  = a;
    endcase
  endfunction
  assign _155_ = \7928 (7'h00, { 49'h0000000000000, _126_[6:0], 7'h00, _106_, _058_, 7'h00 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [6:0] \7931 ;
    input [6:0] a;
    input [83:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7931  = b[6:0];
      12'b??????????1?:
        \7931  = b[13:7];
      12'b?????????1??:
        \7931  = b[20:14];
      12'b????????1???:
        \7931  = b[27:21];
      12'b???????1????:
        \7931  = b[34:28];
      12'b??????1?????:
        \7931  = b[41:35];
      12'b?????1??????:
        \7931  = b[48:42];
      12'b????1???????:
        \7931  = b[55:49];
      12'b???1????????:
        \7931  = b[62:56];
      12'b??1?????????:
        \7931  = b[69:63];
      12'b?1??????????:
        \7931  = b[76:70];
      12'b1???????????:
        \7931  = b[83:77];
      default:
        \7931  = a;
    endcase
  endfunction
  assign _156_ = \7931 (7'h00, { 49'h0000000000000, _126_[13:7], 28'h0000000 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [6:0] \7933 ;
    input [6:0] a;
    input [83:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7933  = b[6:0];
      12'b??????????1?:
        \7933  = b[13:7];
      12'b?????????1??:
        \7933  = b[20:14];
      12'b????????1???:
        \7933  = b[27:21];
      12'b???????1????:
        \7933  = b[34:28];
      12'b??????1?????:
        \7933  = b[41:35];
      12'b?????1??????:
        \7933  = b[48:42];
      12'b????1???????:
        \7933  = b[55:49];
      12'b???1????????:
        \7933  = b[62:56];
      12'b??1?????????:
        \7933  = b[69:63];
      12'b?1??????????:
        \7933  = b[76:70];
      12'b1???????????:
        \7933  = b[83:77];
      default:
        \7933  = a;
    endcase
  endfunction
  assign _157_ = \7933 (7'h00, { 49'h0000000000000, _127_, _109_, _107_, _079_, 7'h00 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [43:0] \7934 ;
    input [43:0] a;
    input [527:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7934  = b[43:0];
      12'b??????????1?:
        \7934  = b[87:44];
      12'b?????????1??:
        \7934  = b[131:88];
      12'b????????1???:
        \7934  = b[175:132];
      12'b???????1????:
        \7934  = b[219:176];
      12'b??????1?????:
        \7934  = b[263:220];
      12'b?????1??????:
        \7934  = b[307:264];
      12'b????1???????:
        \7934  = b[351:308];
      12'b???1????????:
        \7934  = b[395:352];
      12'b??1?????????:
        \7934  = b[439:396];
      12'b?1??????????:
        \7934  = b[483:440];
      12'b1???????????:
        \7934  = b[527:484];
      default:
        \7934  = a;
    endcase
  endfunction
  assign _158_ = \7934 (_189_, { _153_, _207_, _205_, _203_, _189_, _201_, _189_, _199_, _189_, _189_, _195_, _193_ }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [0:0] \7935 ;
    input [0:0] a;
    input [11:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7935  = b[0:0];
      12'b??????????1?:
        \7935  = b[1:1];
      12'b?????????1??:
        \7935  = b[2:2];
      12'b????????1???:
        \7935  = b[3:3];
      12'b???????1????:
        \7935  = b[4:4];
      12'b??????1?????:
        \7935  = b[5:5];
      12'b?????1??????:
        \7935  = b[6:6];
      12'b????1???????:
        \7935  = b[7:7];
      12'b???1????????:
        \7935  = b[8:8];
      12'b??1?????????:
        \7935  = b[9:9];
      12'b?1??????????:
        \7935  = b[10:10];
      12'b1???????????:
        \7935  = b[11:11];
      default:
        \7935  = a;
    endcase
  endfunction
  assign _159_ = \7935 (1'h0, { 9'h001, \f_in.insn [15], 2'h0 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [0:0] \7940 ;
    input [0:0] a;
    input [11:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7940  = b[0:0];
      12'b??????????1?:
        \7940  = b[1:1];
      12'b?????????1??:
        \7940  = b[2:2];
      12'b????????1???:
        \7940  = b[3:3];
      12'b???????1????:
        \7940  = b[4:4];
      12'b??????1?????:
        \7940  = b[5:5];
      12'b?????1??????:
        \7940  = b[6:6];
      12'b????1???????:
        \7940  = b[7:7];
      12'b???1????????:
        \7940  = b[8:8];
      12'b??1?????????:
        \7940  = b[9:9];
      12'b?1??????????:
        \7940  = b[10:10];
      12'b1???????????:
        \7940  = b[11:11];
      default:
        \7940  = a;
    endcase
  endfunction
  assign _160_ = \7940 (1'h0, { 2'h0, _146_, 1'h0, _136_, 1'h0, _131_[0], _112_, 2'h0, _102_, _034_ }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [1:0] \7943 ;
    input [1:0] a;
    input [23:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7943  = b[1:0];
      12'b??????????1?:
        \7943  = b[3:2];
      12'b?????????1??:
        \7943  = b[5:4];
      12'b????????1???:
        \7943  = b[7:6];
      12'b???????1????:
        \7943  = b[9:8];
      12'b??????1?????:
        \7943  = b[11:10];
      12'b?????1??????:
        \7943  = b[13:12];
      12'b????1???????:
        \7943  = b[15:14];
      12'b???1????????:
        \7943  = b[17:16];
      12'b??1?????????:
        \7943  = b[19:18];
      12'b?1??????????:
        \7943  = b[21:20];
      12'b1???????????:
        \7943  = b[23:22];
      default:
        \7943  = a;
    endcase
  endfunction
  assign _161_ = \7943 (2'h0, { 12'h000, _131_[2:1], 6'h00, _094_, 2'h0 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [41:0] \7946 ;
    input [41:0] a;
    input [503:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7946  = b[41:0];
      12'b??????????1?:
        \7946  = b[83:42];
      12'b?????????1??:
        \7946  = b[125:84];
      12'b????????1???:
        \7946  = b[167:126];
      12'b???????1????:
        \7946  = b[209:168];
      12'b??????1?????:
        \7946  = b[251:210];
      12'b?????1??????:
        \7946  = b[293:252];
      12'b????1???????:
        \7946  = b[335:294];
      12'b???1????????:
        \7946  = b[377:336];
      12'b??1?????????:
        \7946  = b[419:378];
      12'b?1??????????:
        \7946  = b[461:420];
      12'b1???????????:
        \7946  = b[503:462];
      default:
        \7946  = a;
    endcase
  endfunction
  assign _162_ = \7946 (42'h00000000000, { 252'h000000000000000000000000000000000000000000000000000000000000000, _131_[44:3], 210'h00000000000000000000000000000000000000000000000000000 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [1:0] \7948 ;
    input [1:0] a;
    input [23:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7948  = b[1:0];
      12'b??????????1?:
        \7948  = b[3:2];
      12'b?????????1??:
        \7948  = b[5:4];
      12'b????????1???:
        \7948  = b[7:6];
      12'b???????1????:
        \7948  = b[9:8];
      12'b??????1?????:
        \7948  = b[11:10];
      12'b?????1??????:
        \7948  = b[13:12];
      12'b????1???????:
        \7948  = b[15:14];
      12'b???1????????:
        \7948  = b[17:16];
      12'b??1?????????:
        \7948  = b[19:18];
      12'b?1??????????:
        \7948  = b[21:20];
      12'b1???????????:
        \7948  = b[23:22];
      default:
        \7948  = a;
    endcase
  endfunction
  assign _163_ = \7948 (2'h0, { 20'h00000, _095_, 2'h0 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  function [23:0] \7957 ;
    input [23:0] a;
    input [287:0] b;
    input [11:0] s;
    (* parallel_case *)
    casez (s)
      12'b???????????1:
        \7957  = b[23:0];
      12'b??????????1?:
        \7957  = b[47:24];
      12'b?????????1??:
        \7957  = b[71:48];
      12'b????????1???:
        \7957  = b[95:72];
      12'b???????1????:
        \7957  = b[119:96];
      12'b??????1?????:
        \7957  = b[143:120];
      12'b?????1??????:
        \7957  = b[167:144];
      12'b????1???????:
        \7957  = b[191:168];
      12'b???1????????:
        \7957  = b[215:192];
      12'b??1?????????:
        \7957  = b[239:216];
      12'b?1??????????:
        \7957  = b[263:240];
      12'b1???????????:
        \7957  = b[287:264];
      default:
        \7957  = a;
    endcase
  endfunction
  assign _164_ = \7957 (24'h000000, { 192'h000000000000000000000000000000000000000000000000, \f_in.insn [25:2], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15], \f_in.insn [15:2], 48'h000000000000 }, { _154_, _149_, _147_, _139_, _137_, _134_, _132_, _128_, _110_, _108_, _103_, _036_ });
  assign _165_ = ri[9:4] == 6'h3d;
  assign _166_ = ri[0] & _165_;
  assign _167_ = _166_ ? 1'h0 : 1'h1;
  assign _168_ = \f_in.fetch_failed  ? _167_ : \f_in.valid ;
  assign _169_ = \f_in.fetch_failed  ? 45'h0000000003d5 : { _162_, _161_, _160_ };
  assign _170_ = \f_in.insn [1] ? 62'h0000000000000000 : \f_in.nia [63:2];
  assign _171_ = \f_in.next_pred_ntaken  ? 1'h0 : _159_;
  assign _172_ = \f_in.next_predicted  ? 1'h1 : _171_;
  assign _173_ = _172_ & \f_in.valid ;
  assign _174_ = ~ flush_in;
  assign _175_ = _173_ & _174_;
  assign _176_ = ~ s[0];
  assign _177_ = _175_ & _176_;
  assign _178_ = ~ \f_in.next_predicted ;
  assign _179_ = _177_ & _178_;
  assign _180_ = br[61:0] + { br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85], br[85:62] };
  assign _181_ = ri[45] ? ri[2:1] : r[120:119];
  assign _182_ = ri[0] ? ri[2:1] : _181_;
  assign _183_ = ri[0] ? ri[42] : r[160];
  assign _184_ = ri[46] ? 1'h1 : _183_;
  assign _185_ = ri[0] ? ri[44:43] : r[162:161];
  assign _186_ = ri[0] ? ri[41:3] : r[159:121];
  assign _187_ = _179_ | br[86];
  assign r = _027_;
  assign rin = { \f_in.big_endian , _172_, _158_, _157_, _156_, _155_, \f_in.insn , \f_in.nia , \f_in.stop_mark , _168_ };
  assign s = _028_;
  assign ri = _029_;
  assign ri_in = { _163_, _169_ };
  assign si = _030_;
  assign br = _031_;
  assign br_in = { _179_, _164_, _170_ };
  assign busy_out = s[0];
  assign flush_out = _187_;
  assign \f_out.redirect  = br[86];
  assign \f_out.redirect_nia  = { _180_, 2'h0 };
  assign \d_out.valid  = r[0];
  assign \d_out.stop_mark  = r[1];
  assign \d_out.nia  = r[65:2];
  assign \d_out.insn  = r[97:66];
  assign \d_out.ispr1  = r[104:98];
  assign \d_out.ispr2  = r[111:105];
  assign \d_out.ispro  = r[118:112];
  assign \d_out.decode  = { _185_, _184_, _186_, _182_ };
  assign \d_out.br_pred  = r[163];
  assign \d_out.big_endian  = r[164];
  assign log_out = 13'hzzzz;
endmodule