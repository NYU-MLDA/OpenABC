module bp_io_cce_05
(
  clk_i,
  reset_i,
  cce_id_i,
  lce_req_i,
  lce_req_v_i,
  lce_req_yumi_o,
  lce_cmd_o,
  lce_cmd_v_o,
  lce_cmd_ready_i,
  io_cmd_o,
  io_cmd_v_o,
  io_cmd_ready_i,
  io_resp_i,
  io_resp_v_i,
  io_resp_yumi_o
);

  input [3:0] cce_id_i;
  input [118:0] lce_req_i;
  output [567:0] lce_cmd_o;
  output [571:0] io_cmd_o;
  input [571:0] io_resp_i;
  input clk_i;
  input reset_i;
  input lce_req_v_i;
  input lce_cmd_ready_i;
  input io_cmd_ready_i;
  input io_resp_v_i;
  output lce_req_yumi_o;
  output lce_cmd_v_o;
  output io_cmd_v_o;
  output io_resp_yumi_o;
  wire [567:0] lce_cmd_o;
  wire [571:0] io_cmd_o;
  wire lce_req_yumi_o,lce_cmd_v_o,io_cmd_v_o,io_resp_yumi_o,N0,N1,N2,N3,N4,
  lce_cmd_o_8_,lce_cmd_o_5_,lce_cmd_o_4_,lce_cmd_o_3_,lce_cmd_o_2_,lce_cmd_o_1_,lce_cmd_o_0_,
  io_cmd_o_123_,io_cmd_o_122_,io_cmd_o_121_,io_cmd_o_120_,io_cmd_o_119_,
  io_cmd_o_118_,io_cmd_o_117_,io_cmd_o_116_,io_cmd_o_115_,io_cmd_o_114_,io_cmd_o_113_,
  io_cmd_o_112_,io_cmd_o_111_,io_cmd_o_110_,io_cmd_o_109_,io_cmd_o_108_,io_cmd_o_107_,
  io_cmd_o_106_,io_cmd_o_105_,io_cmd_o_104_,io_cmd_o_103_,io_cmd_o_102_,
  io_cmd_o_101_,io_cmd_o_100_,io_cmd_o_99_,io_cmd_o_98_,io_cmd_o_97_,io_cmd_o_96_,io_cmd_o_95_,
  io_cmd_o_94_,io_cmd_o_93_,io_cmd_o_92_,io_cmd_o_91_,io_cmd_o_90_,io_cmd_o_89_,
  io_cmd_o_88_,io_cmd_o_87_,io_cmd_o_86_,io_cmd_o_85_,io_cmd_o_84_,io_cmd_o_83_,
  io_cmd_o_82_,io_cmd_o_81_,io_cmd_o_80_,io_cmd_o_79_,io_cmd_o_78_,io_cmd_o_77_,
  io_cmd_o_76_,io_cmd_o_75_,io_cmd_o_74_,io_cmd_o_73_,io_cmd_o_72_,io_cmd_o_71_,
  io_cmd_o_70_,io_cmd_o_69_,io_cmd_o_68_,io_cmd_o_67_,io_cmd_o_66_,io_cmd_o_65_,
  io_cmd_o_64_,io_cmd_o_63_,io_cmd_o_62_,io_cmd_o_61_,io_cmd_o_60_,io_cmd_o_59_,
  io_cmd_o_58_,io_cmd_o_57_,io_cmd_o_56_,io_cmd_o_55_,io_cmd_o_54_,io_cmd_o_43_,io_cmd_o_42_,
  io_cmd_o_41_,io_cmd_o_40_,io_cmd_o_39_,io_cmd_o_38_,io_cmd_o_37_,io_cmd_o_36_,
  io_cmd_o_35_,io_cmd_o_34_,io_cmd_o_33_,io_cmd_o_32_,io_cmd_o_31_,io_cmd_o_30_,
  io_cmd_o_29_,io_cmd_o_28_,io_cmd_o_27_,io_cmd_o_26_,io_cmd_o_25_,io_cmd_o_24_,
  io_cmd_o_23_,io_cmd_o_22_,io_cmd_o_21_,io_cmd_o_20_,io_cmd_o_19_,io_cmd_o_18_,
  io_cmd_o_17_,io_cmd_o_16_,io_cmd_o_15_,io_cmd_o_14_,io_cmd_o_13_,io_cmd_o_12_,
  io_cmd_o_11_,io_cmd_o_10_,io_cmd_o_9_,io_cmd_o_8_,io_cmd_o_7_,io_cmd_o_6_,io_cmd_o_5_,
  io_cmd_o_4_,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,N26;
  assign io_cmd_o[1] = 1'b1;
  assign lce_cmd_o[6] = 1'b1;
  assign io_cmd_o[2] = 1'b0;
  assign io_cmd_o[3] = 1'b0;
  assign io_cmd_o[46] = 1'b0;
  assign io_cmd_o[47] = 1'b0;
  assign io_cmd_o[48] = 1'b0;
  assign io_cmd_o[49] = 1'b0;
  assign io_cmd_o[50] = 1'b0;
  assign io_cmd_o[51] = 1'b0;
  assign io_cmd_o[52] = 1'b0;
  assign io_cmd_o[53] = 1'b0;
  assign io_cmd_o[124] = 1'b0;
  assign io_cmd_o[125] = 1'b0;
  assign io_cmd_o[126] = 1'b0;
  assign io_cmd_o[127] = 1'b0;
  assign io_cmd_o[128] = 1'b0;
  assign io_cmd_o[129] = 1'b0;
  assign io_cmd_o[130] = 1'b0;
  assign io_cmd_o[131] = 1'b0;
  assign io_cmd_o[132] = 1'b0;
  assign io_cmd_o[133] = 1'b0;
  assign io_cmd_o[134] = 1'b0;
  assign io_cmd_o[135] = 1'b0;
  assign io_cmd_o[136] = 1'b0;
  assign io_cmd_o[137] = 1'b0;
  assign io_cmd_o[138] = 1'b0;
  assign io_cmd_o[139] = 1'b0;
  assign io_cmd_o[140] = 1'b0;
  assign io_cmd_o[141] = 1'b0;
  assign io_cmd_o[142] = 1'b0;
  assign io_cmd_o[143] = 1'b0;
  assign io_cmd_o[144] = 1'b0;
  assign io_cmd_o[145] = 1'b0;
  assign io_cmd_o[146] = 1'b0;
  assign io_cmd_o[147] = 1'b0;
  assign io_cmd_o[148] = 1'b0;
  assign io_cmd_o[149] = 1'b0;
  assign io_cmd_o[150] = 1'b0;
  assign io_cmd_o[151] = 1'b0;
  assign io_cmd_o[152] = 1'b0;
  assign io_cmd_o[153] = 1'b0;
  assign io_cmd_o[154] = 1'b0;
  assign io_cmd_o[155] = 1'b0;
  assign io_cmd_o[156] = 1'b0;
  assign io_cmd_o[157] = 1'b0;
  assign io_cmd_o[158] = 1'b0;
  assign io_cmd_o[159] = 1'b0;
  assign io_cmd_o[160] = 1'b0;
  assign io_cmd_o[161] = 1'b0;
  assign io_cmd_o[162] = 1'b0;
  assign io_cmd_o[163] = 1'b0;
  assign io_cmd_o[164] = 1'b0;
  assign io_cmd_o[165] = 1'b0;
  assign io_cmd_o[166] = 1'b0;
  assign io_cmd_o[167] = 1'b0;
  assign io_cmd_o[168] = 1'b0;
  assign io_cmd_o[169] = 1'b0;
  assign io_cmd_o[170] = 1'b0;
  assign io_cmd_o[171] = 1'b0;
  assign io_cmd_o[172] = 1'b0;
  assign io_cmd_o[173] = 1'b0;
  assign io_cmd_o[174] = 1'b0;
  assign io_cmd_o[175] = 1'b0;
  assign io_cmd_o[176] = 1'b0;
  assign io_cmd_o[177] = 1'b0;
  assign io_cmd_o[178] = 1'b0;
  assign io_cmd_o[179] = 1'b0;
  assign io_cmd_o[180] = 1'b0;
  assign io_cmd_o[181] = 1'b0;
  assign io_cmd_o[182] = 1'b0;
  assign io_cmd_o[183] = 1'b0;
  assign io_cmd_o[184] = 1'b0;
  assign io_cmd_o[185] = 1'b0;
  assign io_cmd_o[186] = 1'b0;
  assign io_cmd_o[187] = 1'b0;
  assign io_cmd_o[188] = 1'b0;
  assign io_cmd_o[189] = 1'b0;
  assign io_cmd_o[190] = 1'b0;
  assign io_cmd_o[191] = 1'b0;
  assign io_cmd_o[192] = 1'b0;
  assign io_cmd_o[193] = 1'b0;
  assign io_cmd_o[194] = 1'b0;
  assign io_cmd_o[195] = 1'b0;
  assign io_cmd_o[196] = 1'b0;
  assign io_cmd_o[197] = 1'b0;
  assign io_cmd_o[198] = 1'b0;
  assign io_cmd_o[199] = 1'b0;
  assign io_cmd_o[200] = 1'b0;
  assign io_cmd_o[201] = 1'b0;
  assign io_cmd_o[202] = 1'b0;
  assign io_cmd_o[203] = 1'b0;
  assign io_cmd_o[204] = 1'b0;
  assign io_cmd_o[205] = 1'b0;
  assign io_cmd_o[206] = 1'b0;
  assign io_cmd_o[207] = 1'b0;
  assign io_cmd_o[208] = 1'b0;
  assign io_cmd_o[209] = 1'b0;
  assign io_cmd_o[210] = 1'b0;
  assign io_cmd_o[211] = 1'b0;
  assign io_cmd_o[212] = 1'b0;
  assign io_cmd_o[213] = 1'b0;
  assign io_cmd_o[214] = 1'b0;
  assign io_cmd_o[215] = 1'b0;
  assign io_cmd_o[216] = 1'b0;
  assign io_cmd_o[217] = 1'b0;
  assign io_cmd_o[218] = 1'b0;
  assign io_cmd_o[219] = 1'b0;
  assign io_cmd_o[220] = 1'b0;
  assign io_cmd_o[221] = 1'b0;
  assign io_cmd_o[222] = 1'b0;
  assign io_cmd_o[223] = 1'b0;
  assign io_cmd_o[224] = 1'b0;
  assign io_cmd_o[225] = 1'b0;
  assign io_cmd_o[226] = 1'b0;
  assign io_cmd_o[227] = 1'b0;
  assign io_cmd_o[228] = 1'b0;
  assign io_cmd_o[229] = 1'b0;
  assign io_cmd_o[230] = 1'b0;
  assign io_cmd_o[231] = 1'b0;
  assign io_cmd_o[232] = 1'b0;
  assign io_cmd_o[233] = 1'b0;
  assign io_cmd_o[234] = 1'b0;
  assign io_cmd_o[235] = 1'b0;
  assign io_cmd_o[236] = 1'b0;
  assign io_cmd_o[237] = 1'b0;
  assign io_cmd_o[238] = 1'b0;
  assign io_cmd_o[239] = 1'b0;
  assign io_cmd_o[240] = 1'b0;
  assign io_cmd_o[241] = 1'b0;
  assign io_cmd_o[242] = 1'b0;
  assign io_cmd_o[243] = 1'b0;
  assign io_cmd_o[244] = 1'b0;
  assign io_cmd_o[245] = 1'b0;
  assign io_cmd_o[246] = 1'b0;
  assign io_cmd_o[247] = 1'b0;
  assign io_cmd_o[248] = 1'b0;
  assign io_cmd_o[249] = 1'b0;
  assign io_cmd_o[250] = 1'b0;
  assign io_cmd_o[251] = 1'b0;
  assign io_cmd_o[252] = 1'b0;
  assign io_cmd_o[253] = 1'b0;
  assign io_cmd_o[254] = 1'b0;
  assign io_cmd_o[255] = 1'b0;
  assign io_cmd_o[256] = 1'b0;
  assign io_cmd_o[257] = 1'b0;
  assign io_cmd_o[258] = 1'b0;
  assign io_cmd_o[259] = 1'b0;
  assign io_cmd_o[260] = 1'b0;
  assign io_cmd_o[261] = 1'b0;
  assign io_cmd_o[262] = 1'b0;
  assign io_cmd_o[263] = 1'b0;
  assign io_cmd_o[264] = 1'b0;
  assign io_cmd_o[265] = 1'b0;
  assign io_cmd_o[266] = 1'b0;
  assign io_cmd_o[267] = 1'b0;
  assign io_cmd_o[268] = 1'b0;
  assign io_cmd_o[269] = 1'b0;
  assign io_cmd_o[270] = 1'b0;
  assign io_cmd_o[271] = 1'b0;
  assign io_cmd_o[272] = 1'b0;
  assign io_cmd_o[273] = 1'b0;
  assign io_cmd_o[274] = 1'b0;
  assign io_cmd_o[275] = 1'b0;
  assign io_cmd_o[276] = 1'b0;
  assign io_cmd_o[277] = 1'b0;
  assign io_cmd_o[278] = 1'b0;
  assign io_cmd_o[279] = 1'b0;
  assign io_cmd_o[280] = 1'b0;
  assign io_cmd_o[281] = 1'b0;
  assign io_cmd_o[282] = 1'b0;
  assign io_cmd_o[283] = 1'b0;
  assign io_cmd_o[284] = 1'b0;
  assign io_cmd_o[285] = 1'b0;
  assign io_cmd_o[286] = 1'b0;
  assign io_cmd_o[287] = 1'b0;
  assign io_cmd_o[288] = 1'b0;
  assign io_cmd_o[289] = 1'b0;
  assign io_cmd_o[290] = 1'b0;
  assign io_cmd_o[291] = 1'b0;
  assign io_cmd_o[292] = 1'b0;
  assign io_cmd_o[293] = 1'b0;
  assign io_cmd_o[294] = 1'b0;
  assign io_cmd_o[295] = 1'b0;
  assign io_cmd_o[296] = 1'b0;
  assign io_cmd_o[297] = 1'b0;
  assign io_cmd_o[298] = 1'b0;
  assign io_cmd_o[299] = 1'b0;
  assign io_cmd_o[300] = 1'b0;
  assign io_cmd_o[301] = 1'b0;
  assign io_cmd_o[302] = 1'b0;
  assign io_cmd_o[303] = 1'b0;
  assign io_cmd_o[304] = 1'b0;
  assign io_cmd_o[305] = 1'b0;
  assign io_cmd_o[306] = 1'b0;
  assign io_cmd_o[307] = 1'b0;
  assign io_cmd_o[308] = 1'b0;
  assign io_cmd_o[309] = 1'b0;
  assign io_cmd_o[310] = 1'b0;
  assign io_cmd_o[311] = 1'b0;
  assign io_cmd_o[312] = 1'b0;
  assign io_cmd_o[313] = 1'b0;
  assign io_cmd_o[314] = 1'b0;
  assign io_cmd_o[315] = 1'b0;
  assign io_cmd_o[316] = 1'b0;
  assign io_cmd_o[317] = 1'b0;
  assign io_cmd_o[318] = 1'b0;
  assign io_cmd_o[319] = 1'b0;
  assign io_cmd_o[320] = 1'b0;
  assign io_cmd_o[321] = 1'b0;
  assign io_cmd_o[322] = 1'b0;
  assign io_cmd_o[323] = 1'b0;
  assign io_cmd_o[324] = 1'b0;
  assign io_cmd_o[325] = 1'b0;
  assign io_cmd_o[326] = 1'b0;
  assign io_cmd_o[327] = 1'b0;
  assign io_cmd_o[328] = 1'b0;
  assign io_cmd_o[329] = 1'b0;
  assign io_cmd_o[330] = 1'b0;
  assign io_cmd_o[331] = 1'b0;
  assign io_cmd_o[332] = 1'b0;
  assign io_cmd_o[333] = 1'b0;
  assign io_cmd_o[334] = 1'b0;
  assign io_cmd_o[335] = 1'b0;
  assign io_cmd_o[336] = 1'b0;
  assign io_cmd_o[337] = 1'b0;
  assign io_cmd_o[338] = 1'b0;
  assign io_cmd_o[339] = 1'b0;
  assign io_cmd_o[340] = 1'b0;
  assign io_cmd_o[341] = 1'b0;
  assign io_cmd_o[342] = 1'b0;
  assign io_cmd_o[343] = 1'b0;
  assign io_cmd_o[344] = 1'b0;
  assign io_cmd_o[345] = 1'b0;
  assign io_cmd_o[346] = 1'b0;
  assign io_cmd_o[347] = 1'b0;
  assign io_cmd_o[348] = 1'b0;
  assign io_cmd_o[349] = 1'b0;
  assign io_cmd_o[350] = 1'b0;
  assign io_cmd_o[351] = 1'b0;
  assign io_cmd_o[352] = 1'b0;
  assign io_cmd_o[353] = 1'b0;
  assign io_cmd_o[354] = 1'b0;
  assign io_cmd_o[355] = 1'b0;
  assign io_cmd_o[356] = 1'b0;
  assign io_cmd_o[357] = 1'b0;
  assign io_cmd_o[358] = 1'b0;
  assign io_cmd_o[359] = 1'b0;
  assign io_cmd_o[360] = 1'b0;
  assign io_cmd_o[361] = 1'b0;
  assign io_cmd_o[362] = 1'b0;
  assign io_cmd_o[363] = 1'b0;
  assign io_cmd_o[364] = 1'b0;
  assign io_cmd_o[365] = 1'b0;
  assign io_cmd_o[366] = 1'b0;
  assign io_cmd_o[367] = 1'b0;
  assign io_cmd_o[368] = 1'b0;
  assign io_cmd_o[369] = 1'b0;
  assign io_cmd_o[370] = 1'b0;
  assign io_cmd_o[371] = 1'b0;
  assign io_cmd_o[372] = 1'b0;
  assign io_cmd_o[373] = 1'b0;
  assign io_cmd_o[374] = 1'b0;
  assign io_cmd_o[375] = 1'b0;
  assign io_cmd_o[376] = 1'b0;
  assign io_cmd_o[377] = 1'b0;
  assign io_cmd_o[378] = 1'b0;
  assign io_cmd_o[379] = 1'b0;
  assign io_cmd_o[380] = 1'b0;
  assign io_cmd_o[381] = 1'b0;
  assign io_cmd_o[382] = 1'b0;
  assign io_cmd_o[383] = 1'b0;
  assign io_cmd_o[384] = 1'b0;
  assign io_cmd_o[385] = 1'b0;
  assign io_cmd_o[386] = 1'b0;
  assign io_cmd_o[387] = 1'b0;
  assign io_cmd_o[388] = 1'b0;
  assign io_cmd_o[389] = 1'b0;
  assign io_cmd_o[390] = 1'b0;
  assign io_cmd_o[391] = 1'b0;
  assign io_cmd_o[392] = 1'b0;
  assign io_cmd_o[393] = 1'b0;
  assign io_cmd_o[394] = 1'b0;
  assign io_cmd_o[395] = 1'b0;
  assign io_cmd_o[396] = 1'b0;
  assign io_cmd_o[397] = 1'b0;
  assign io_cmd_o[398] = 1'b0;
  assign io_cmd_o[399] = 1'b0;
  assign io_cmd_o[400] = 1'b0;
  assign io_cmd_o[401] = 1'b0;
  assign io_cmd_o[402] = 1'b0;
  assign io_cmd_o[403] = 1'b0;
  assign io_cmd_o[404] = 1'b0;
  assign io_cmd_o[405] = 1'b0;
  assign io_cmd_o[406] = 1'b0;
  assign io_cmd_o[407] = 1'b0;
  assign io_cmd_o[408] = 1'b0;
  assign io_cmd_o[409] = 1'b0;
  assign io_cmd_o[410] = 1'b0;
  assign io_cmd_o[411] = 1'b0;
  assign io_cmd_o[412] = 1'b0;
  assign io_cmd_o[413] = 1'b0;
  assign io_cmd_o[414] = 1'b0;
  assign io_cmd_o[415] = 1'b0;
  assign io_cmd_o[416] = 1'b0;
  assign io_cmd_o[417] = 1'b0;
  assign io_cmd_o[418] = 1'b0;
  assign io_cmd_o[419] = 1'b0;
  assign io_cmd_o[420] = 1'b0;
  assign io_cmd_o[421] = 1'b0;
  assign io_cmd_o[422] = 1'b0;
  assign io_cmd_o[423] = 1'b0;
  assign io_cmd_o[424] = 1'b0;
  assign io_cmd_o[425] = 1'b0;
  assign io_cmd_o[426] = 1'b0;
  assign io_cmd_o[427] = 1'b0;
  assign io_cmd_o[428] = 1'b0;
  assign io_cmd_o[429] = 1'b0;
  assign io_cmd_o[430] = 1'b0;
  assign io_cmd_o[431] = 1'b0;
  assign io_cmd_o[432] = 1'b0;
  assign io_cmd_o[433] = 1'b0;
  assign io_cmd_o[434] = 1'b0;
  assign io_cmd_o[435] = 1'b0;
  assign io_cmd_o[436] = 1'b0;
  assign io_cmd_o[437] = 1'b0;
  assign io_cmd_o[438] = 1'b0;
  assign io_cmd_o[439] = 1'b0;
  assign io_cmd_o[440] = 1'b0;
  assign io_cmd_o[441] = 1'b0;
  assign io_cmd_o[442] = 1'b0;
  assign io_cmd_o[443] = 1'b0;
  assign io_cmd_o[444] = 1'b0;
  assign io_cmd_o[445] = 1'b0;
  assign io_cmd_o[446] = 1'b0;
  assign io_cmd_o[447] = 1'b0;
  assign io_cmd_o[448] = 1'b0;
  assign io_cmd_o[449] = 1'b0;
  assign io_cmd_o[450] = 1'b0;
  assign io_cmd_o[451] = 1'b0;
  assign io_cmd_o[452] = 1'b0;
  assign io_cmd_o[453] = 1'b0;
  assign io_cmd_o[454] = 1'b0;
  assign io_cmd_o[455] = 1'b0;
  assign io_cmd_o[456] = 1'b0;
  assign io_cmd_o[457] = 1'b0;
  assign io_cmd_o[458] = 1'b0;
  assign io_cmd_o[459] = 1'b0;
  assign io_cmd_o[460] = 1'b0;
  assign io_cmd_o[461] = 1'b0;
  assign io_cmd_o[462] = 1'b0;
  assign io_cmd_o[463] = 1'b0;
  assign io_cmd_o[464] = 1'b0;
  assign io_cmd_o[465] = 1'b0;
  assign io_cmd_o[466] = 1'b0;
  assign io_cmd_o[467] = 1'b0;
  assign io_cmd_o[468] = 1'b0;
  assign io_cmd_o[469] = 1'b0;
  assign io_cmd_o[470] = 1'b0;
  assign io_cmd_o[471] = 1'b0;
  assign io_cmd_o[472] = 1'b0;
  assign io_cmd_o[473] = 1'b0;
  assign io_cmd_o[474] = 1'b0;
  assign io_cmd_o[475] = 1'b0;
  assign io_cmd_o[476] = 1'b0;
  assign io_cmd_o[477] = 1'b0;
  assign io_cmd_o[478] = 1'b0;
  assign io_cmd_o[479] = 1'b0;
  assign io_cmd_o[480] = 1'b0;
  assign io_cmd_o[481] = 1'b0;
  assign io_cmd_o[482] = 1'b0;
  assign io_cmd_o[483] = 1'b0;
  assign io_cmd_o[484] = 1'b0;
  assign io_cmd_o[485] = 1'b0;
  assign io_cmd_o[486] = 1'b0;
  assign io_cmd_o[487] = 1'b0;
  assign io_cmd_o[488] = 1'b0;
  assign io_cmd_o[489] = 1'b0;
  assign io_cmd_o[490] = 1'b0;
  assign io_cmd_o[491] = 1'b0;
  assign io_cmd_o[492] = 1'b0;
  assign io_cmd_o[493] = 1'b0;
  assign io_cmd_o[494] = 1'b0;
  assign io_cmd_o[495] = 1'b0;
  assign io_cmd_o[496] = 1'b0;
  assign io_cmd_o[497] = 1'b0;
  assign io_cmd_o[498] = 1'b0;
  assign io_cmd_o[499] = 1'b0;
  assign io_cmd_o[500] = 1'b0;
  assign io_cmd_o[501] = 1'b0;
  assign io_cmd_o[502] = 1'b0;
  assign io_cmd_o[503] = 1'b0;
  assign io_cmd_o[504] = 1'b0;
  assign io_cmd_o[505] = 1'b0;
  assign io_cmd_o[506] = 1'b0;
  assign io_cmd_o[507] = 1'b0;
  assign io_cmd_o[508] = 1'b0;
  assign io_cmd_o[509] = 1'b0;
  assign io_cmd_o[510] = 1'b0;
  assign io_cmd_o[511] = 1'b0;
  assign io_cmd_o[512] = 1'b0;
  assign io_cmd_o[513] = 1'b0;
  assign io_cmd_o[514] = 1'b0;
  assign io_cmd_o[515] = 1'b0;
  assign io_cmd_o[516] = 1'b0;
  assign io_cmd_o[517] = 1'b0;
  assign io_cmd_o[518] = 1'b0;
  assign io_cmd_o[519] = 1'b0;
  assign io_cmd_o[520] = 1'b0;
  assign io_cmd_o[521] = 1'b0;
  assign io_cmd_o[522] = 1'b0;
  assign io_cmd_o[523] = 1'b0;
  assign io_cmd_o[524] = 1'b0;
  assign io_cmd_o[525] = 1'b0;
  assign io_cmd_o[526] = 1'b0;
  assign io_cmd_o[527] = 1'b0;
  assign io_cmd_o[528] = 1'b0;
  assign io_cmd_o[529] = 1'b0;
  assign io_cmd_o[530] = 1'b0;
  assign io_cmd_o[531] = 1'b0;
  assign io_cmd_o[532] = 1'b0;
  assign io_cmd_o[533] = 1'b0;
  assign io_cmd_o[534] = 1'b0;
  assign io_cmd_o[535] = 1'b0;
  assign io_cmd_o[536] = 1'b0;
  assign io_cmd_o[537] = 1'b0;
  assign io_cmd_o[538] = 1'b0;
  assign io_cmd_o[539] = 1'b0;
  assign io_cmd_o[540] = 1'b0;
  assign io_cmd_o[541] = 1'b0;
  assign io_cmd_o[542] = 1'b0;
  assign io_cmd_o[543] = 1'b0;
  assign io_cmd_o[544] = 1'b0;
  assign io_cmd_o[545] = 1'b0;
  assign io_cmd_o[546] = 1'b0;
  assign io_cmd_o[547] = 1'b0;
  assign io_cmd_o[548] = 1'b0;
  assign io_cmd_o[549] = 1'b0;
  assign io_cmd_o[550] = 1'b0;
  assign io_cmd_o[551] = 1'b0;
  assign io_cmd_o[552] = 1'b0;
  assign io_cmd_o[553] = 1'b0;
  assign io_cmd_o[554] = 1'b0;
  assign io_cmd_o[555] = 1'b0;
  assign io_cmd_o[556] = 1'b0;
  assign io_cmd_o[557] = 1'b0;
  assign io_cmd_o[558] = 1'b0;
  assign io_cmd_o[559] = 1'b0;
  assign io_cmd_o[560] = 1'b0;
  assign io_cmd_o[561] = 1'b0;
  assign io_cmd_o[562] = 1'b0;
  assign io_cmd_o[563] = 1'b0;
  assign io_cmd_o[564] = 1'b0;
  assign io_cmd_o[565] = 1'b0;
  assign io_cmd_o[566] = 1'b0;
  assign io_cmd_o[567] = 1'b0;
  assign io_cmd_o[568] = 1'b0;
  assign io_cmd_o[569] = 1'b0;
  assign io_cmd_o[570] = 1'b0;
  assign io_cmd_o[571] = 1'b0;
  assign lce_cmd_o[10] = 1'b0;
  assign lce_cmd_o[11] = 1'b0;
  assign lce_cmd_o[12] = 1'b0;
  assign io_cmd_v_o = lce_req_yumi_o;
  assign lce_cmd_o[7] = lce_cmd_o_8_;
  assign lce_cmd_o[8] = lce_cmd_o_8_;
  assign lce_cmd_o_5_ = io_resp_i[59];
  assign lce_cmd_o[5] = lce_cmd_o_5_;
  assign lce_cmd_o_4_ = io_resp_i[58];
  assign lce_cmd_o[4] = lce_cmd_o_4_;
  assign lce_cmd_o_3_ = io_resp_i[57];
  assign lce_cmd_o[3] = lce_cmd_o_3_;
  assign lce_cmd_o_2_ = io_resp_i[56];
  assign lce_cmd_o[2] = lce_cmd_o_2_;
  assign lce_cmd_o_1_ = io_resp_i[55];
  assign lce_cmd_o[1] = lce_cmd_o_1_;
  assign lce_cmd_o_0_ = io_resp_i[54];
  assign lce_cmd_o[0] = lce_cmd_o_0_;
  assign io_cmd_o_123_ = lce_req_i[118];
  assign io_cmd_o[123] = io_cmd_o_123_;
  assign io_cmd_o_122_ = lce_req_i[117];
  assign io_cmd_o[122] = io_cmd_o_122_;
  assign io_cmd_o_121_ = lce_req_i[116];
  assign io_cmd_o[121] = io_cmd_o_121_;
  assign io_cmd_o_120_ = lce_req_i[115];
  assign io_cmd_o[120] = io_cmd_o_120_;
  assign io_cmd_o_119_ = lce_req_i[114];
  assign io_cmd_o[119] = io_cmd_o_119_;
  assign io_cmd_o_118_ = lce_req_i[113];
  assign io_cmd_o[118] = io_cmd_o_118_;
  assign io_cmd_o_117_ = lce_req_i[112];
  assign io_cmd_o[117] = io_cmd_o_117_;
  assign io_cmd_o_116_ = lce_req_i[111];
  assign io_cmd_o[116] = io_cmd_o_116_;
  assign io_cmd_o_115_ = lce_req_i[110];
  assign io_cmd_o[115] = io_cmd_o_115_;
  assign io_cmd_o_114_ = lce_req_i[109];
  assign io_cmd_o[114] = io_cmd_o_114_;
  assign io_cmd_o_113_ = lce_req_i[108];
  assign io_cmd_o[113] = io_cmd_o_113_;
  assign io_cmd_o_112_ = lce_req_i[107];
  assign io_cmd_o[112] = io_cmd_o_112_;
  assign io_cmd_o_111_ = lce_req_i[106];
  assign io_cmd_o[111] = io_cmd_o_111_;
  assign io_cmd_o_110_ = lce_req_i[105];
  assign io_cmd_o[110] = io_cmd_o_110_;
  assign io_cmd_o_109_ = lce_req_i[104];
  assign io_cmd_o[109] = io_cmd_o_109_;
  assign io_cmd_o_108_ = lce_req_i[103];
  assign io_cmd_o[108] = io_cmd_o_108_;
  assign io_cmd_o_107_ = lce_req_i[102];
  assign io_cmd_o[107] = io_cmd_o_107_;
  assign io_cmd_o_106_ = lce_req_i[101];
  assign io_cmd_o[106] = io_cmd_o_106_;
  assign io_cmd_o_105_ = lce_req_i[100];
  assign io_cmd_o[105] = io_cmd_o_105_;
  assign io_cmd_o_104_ = lce_req_i[99];
  assign io_cmd_o[104] = io_cmd_o_104_;
  assign io_cmd_o_103_ = lce_req_i[98];
  assign io_cmd_o[103] = io_cmd_o_103_;
  assign io_cmd_o_102_ = lce_req_i[97];
  assign io_cmd_o[102] = io_cmd_o_102_;
  assign io_cmd_o_101_ = lce_req_i[96];
  assign io_cmd_o[101] = io_cmd_o_101_;
  assign io_cmd_o_100_ = lce_req_i[95];
  assign io_cmd_o[100] = io_cmd_o_100_;
  assign io_cmd_o_99_ = lce_req_i[94];
  assign io_cmd_o[99] = io_cmd_o_99_;
  assign io_cmd_o_98_ = lce_req_i[93];
  assign io_cmd_o[98] = io_cmd_o_98_;
  assign io_cmd_o_97_ = lce_req_i[92];
  assign io_cmd_o[97] = io_cmd_o_97_;
  assign io_cmd_o_96_ = lce_req_i[91];
  assign io_cmd_o[96] = io_cmd_o_96_;
  assign io_cmd_o_95_ = lce_req_i[90];
  assign io_cmd_o[95] = io_cmd_o_95_;
  assign io_cmd_o_94_ = lce_req_i[89];
  assign io_cmd_o[94] = io_cmd_o_94_;
  assign io_cmd_o_93_ = lce_req_i[88];
  assign io_cmd_o[93] = io_cmd_o_93_;
  assign io_cmd_o_92_ = lce_req_i[87];
  assign io_cmd_o[92] = io_cmd_o_92_;
  assign io_cmd_o_91_ = lce_req_i[86];
  assign io_cmd_o[91] = io_cmd_o_91_;
  assign io_cmd_o_90_ = lce_req_i[85];
  assign io_cmd_o[90] = io_cmd_o_90_;
  assign io_cmd_o_89_ = lce_req_i[84];
  assign io_cmd_o[89] = io_cmd_o_89_;
  assign io_cmd_o_88_ = lce_req_i[83];
  assign io_cmd_o[88] = io_cmd_o_88_;
  assign io_cmd_o_87_ = lce_req_i[82];
  assign io_cmd_o[87] = io_cmd_o_87_;
  assign io_cmd_o_86_ = lce_req_i[81];
  assign io_cmd_o[86] = io_cmd_o_86_;
  assign io_cmd_o_85_ = lce_req_i[80];
  assign io_cmd_o[85] = io_cmd_o_85_;
  assign io_cmd_o_84_ = lce_req_i[79];
  assign io_cmd_o[84] = io_cmd_o_84_;
  assign io_cmd_o_83_ = lce_req_i[78];
  assign io_cmd_o[83] = io_cmd_o_83_;
  assign io_cmd_o_82_ = lce_req_i[77];
  assign io_cmd_o[82] = io_cmd_o_82_;
  assign io_cmd_o_81_ = lce_req_i[76];
  assign io_cmd_o[81] = io_cmd_o_81_;
  assign io_cmd_o_80_ = lce_req_i[75];
  assign io_cmd_o[80] = io_cmd_o_80_;
  assign io_cmd_o_79_ = lce_req_i[74];
  assign io_cmd_o[79] = io_cmd_o_79_;
  assign io_cmd_o_78_ = lce_req_i[73];
  assign io_cmd_o[78] = io_cmd_o_78_;
  assign io_cmd_o_77_ = lce_req_i[72];
  assign io_cmd_o[77] = io_cmd_o_77_;
  assign io_cmd_o_76_ = lce_req_i[71];
  assign io_cmd_o[76] = io_cmd_o_76_;
  assign io_cmd_o_75_ = lce_req_i[70];
  assign io_cmd_o[75] = io_cmd_o_75_;
  assign io_cmd_o_74_ = lce_req_i[69];
  assign io_cmd_o[74] = io_cmd_o_74_;
  assign io_cmd_o_73_ = lce_req_i[68];
  assign io_cmd_o[73] = io_cmd_o_73_;
  assign io_cmd_o_72_ = lce_req_i[67];
  assign io_cmd_o[72] = io_cmd_o_72_;
  assign io_cmd_o_71_ = lce_req_i[66];
  assign io_cmd_o[71] = io_cmd_o_71_;
  assign io_cmd_o_70_ = lce_req_i[65];
  assign io_cmd_o[70] = io_cmd_o_70_;
  assign io_cmd_o_69_ = lce_req_i[64];
  assign io_cmd_o[69] = io_cmd_o_69_;
  assign io_cmd_o_68_ = lce_req_i[63];
  assign io_cmd_o[68] = io_cmd_o_68_;
  assign io_cmd_o_67_ = lce_req_i[62];
  assign io_cmd_o[67] = io_cmd_o_67_;
  assign io_cmd_o_66_ = lce_req_i[61];
  assign io_cmd_o[66] = io_cmd_o_66_;
  assign io_cmd_o_65_ = lce_req_i[60];
  assign io_cmd_o[65] = io_cmd_o_65_;
  assign io_cmd_o_64_ = lce_req_i[59];
  assign io_cmd_o[64] = io_cmd_o_64_;
  assign io_cmd_o_63_ = lce_req_i[58];
  assign io_cmd_o[63] = io_cmd_o_63_;
  assign io_cmd_o_62_ = lce_req_i[57];
  assign io_cmd_o[62] = io_cmd_o_62_;
  assign io_cmd_o_61_ = lce_req_i[56];
  assign io_cmd_o[61] = io_cmd_o_61_;
  assign io_cmd_o_60_ = lce_req_i[55];
  assign io_cmd_o[60] = io_cmd_o_60_;
  assign io_cmd_o_59_ = lce_req_i[9];
  assign io_cmd_o[59] = io_cmd_o_59_;
  assign io_cmd_o_58_ = lce_req_i[8];
  assign io_cmd_o[58] = io_cmd_o_58_;
  assign io_cmd_o_57_ = lce_req_i[7];
  assign io_cmd_o[57] = io_cmd_o_57_;
  assign io_cmd_o_56_ = lce_req_i[6];
  assign io_cmd_o[56] = io_cmd_o_56_;
  assign io_cmd_o_55_ = lce_req_i[5];
  assign io_cmd_o[55] = io_cmd_o_55_;
  assign io_cmd_o_54_ = lce_req_i[4];
  assign io_cmd_o[54] = io_cmd_o_54_;
  assign io_cmd_o_43_ = lce_req_i[52];
  assign io_cmd_o[43] = io_cmd_o_43_;
  assign io_cmd_o_42_ = lce_req_i[51];
  assign io_cmd_o[42] = io_cmd_o_42_;
  assign io_cmd_o_41_ = lce_req_i[50];
  assign io_cmd_o[41] = io_cmd_o_41_;
  assign io_cmd_o_40_ = lce_req_i[49];
  assign io_cmd_o[40] = io_cmd_o_40_;
  assign io_cmd_o_39_ = lce_req_i[48];
  assign io_cmd_o[39] = io_cmd_o_39_;
  assign io_cmd_o_38_ = lce_req_i[47];
  assign io_cmd_o[38] = io_cmd_o_38_;
  assign io_cmd_o_37_ = lce_req_i[46];
  assign io_cmd_o[37] = io_cmd_o_37_;
  assign io_cmd_o_36_ = lce_req_i[45];
  assign io_cmd_o[36] = io_cmd_o_36_;
  assign io_cmd_o_35_ = lce_req_i[44];
  assign io_cmd_o[35] = io_cmd_o_35_;
  assign io_cmd_o_34_ = lce_req_i[43];
  assign io_cmd_o[34] = io_cmd_o_34_;
  assign io_cmd_o_33_ = lce_req_i[42];
  assign io_cmd_o[33] = io_cmd_o_33_;
  assign io_cmd_o_32_ = lce_req_i[41];
  assign io_cmd_o[32] = io_cmd_o_32_;
  assign io_cmd_o_31_ = lce_req_i[40];
  assign io_cmd_o[31] = io_cmd_o_31_;
  assign io_cmd_o_30_ = lce_req_i[39];
  assign io_cmd_o[30] = io_cmd_o_30_;
  assign io_cmd_o_29_ = lce_req_i[38];
  assign io_cmd_o[29] = io_cmd_o_29_;
  assign io_cmd_o_28_ = lce_req_i[37];
  assign io_cmd_o[28] = io_cmd_o_28_;
  assign io_cmd_o_27_ = lce_req_i[36];
  assign io_cmd_o[27] = io_cmd_o_27_;
  assign io_cmd_o_26_ = lce_req_i[35];
  assign io_cmd_o[26] = io_cmd_o_26_;
  assign io_cmd_o_25_ = lce_req_i[34];
  assign io_cmd_o[25] = io_cmd_o_25_;
  assign io_cmd_o_24_ = lce_req_i[33];
  assign io_cmd_o[24] = io_cmd_o_24_;
  assign io_cmd_o_23_ = lce_req_i[32];
  assign io_cmd_o[23] = io_cmd_o_23_;
  assign io_cmd_o_22_ = lce_req_i[31];
  assign io_cmd_o[22] = io_cmd_o_22_;
  assign io_cmd_o_21_ = lce_req_i[30];
  assign io_cmd_o[21] = io_cmd_o_21_;
  assign io_cmd_o_20_ = lce_req_i[29];
  assign io_cmd_o[20] = io_cmd_o_20_;
  assign io_cmd_o_19_ = lce_req_i[28];
  assign io_cmd_o[19] = io_cmd_o_19_;
  assign io_cmd_o_18_ = lce_req_i[27];
  assign io_cmd_o[18] = io_cmd_o_18_;
  assign io_cmd_o_17_ = lce_req_i[26];
  assign io_cmd_o[17] = io_cmd_o_17_;
  assign io_cmd_o_16_ = lce_req_i[25];
  assign io_cmd_o[16] = io_cmd_o_16_;
  assign io_cmd_o_15_ = lce_req_i[24];
  assign io_cmd_o[15] = io_cmd_o_15_;
  assign io_cmd_o_14_ = lce_req_i[23];
  assign io_cmd_o[14] = io_cmd_o_14_;
  assign io_cmd_o_13_ = lce_req_i[22];
  assign io_cmd_o[13] = io_cmd_o_13_;
  assign io_cmd_o_12_ = lce_req_i[21];
  assign io_cmd_o[12] = io_cmd_o_12_;
  assign io_cmd_o_11_ = lce_req_i[20];
  assign io_cmd_o[11] = io_cmd_o_11_;
  assign io_cmd_o_10_ = lce_req_i[19];
  assign io_cmd_o[10] = io_cmd_o_10_;
  assign io_cmd_o_9_ = lce_req_i[18];
  assign io_cmd_o[9] = io_cmd_o_9_;
  assign io_cmd_o_8_ = lce_req_i[17];
  assign io_cmd_o[8] = io_cmd_o_8_;
  assign io_cmd_o_7_ = lce_req_i[16];
  assign io_cmd_o[7] = io_cmd_o_7_;
  assign io_cmd_o_6_ = lce_req_i[15];
  assign io_cmd_o[6] = io_cmd_o_6_;
  assign io_cmd_o_5_ = lce_req_i[14];
  assign io_cmd_o[5] = io_cmd_o_5_;
  assign io_cmd_o_4_ = lce_req_i[13];
  assign io_cmd_o[4] = io_cmd_o_4_;
  assign lce_cmd_v_o = io_resp_yumi_o;
  assign N8 = ~io_resp_i[1];
  assign N9 = ~io_resp_i[0];
  assign N10 = io_resp_i[2] | io_resp_i[3];
  assign N11 = N8 | N10;
  assign N12 = N9 | N11;
  assign N13 = ~N12;
  assign N14 = ~lce_req_i[11];
  assign N15 = ~lce_req_i[10];
  assign N16 = N14 | lce_req_i[12];
  assign N17 = N15 | N16;
  assign N18 = ~N17;
  assign N19 = ~lce_req_i[54];
  assign N20 = lce_req_i[53] | N19;
  assign N21 = ~N20;
  assign N22 = ~lce_req_i[53];
  assign N23 = N22 | lce_req_i[54];
  assign N24 = ~N23;
  assign N25 = lce_req_i[53] | lce_req_i[54];
  assign N26 = ~N25;
  assign io_cmd_o[45:44] = (N0)? { 1'b0, 1'b0 } : 
                           (N1)? { 1'b0, 1'b1 } : 
                           (N2)? { 1'b1, 1'b0 } : 
                           (N7)? { 1'b1, 1'b1 } : 1'b0;
  assign N0 = N26;
  assign N1 = N24;
  assign N2 = N21;
  assign lce_cmd_o[567:13] = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, io_resp_i[43:4], cce_id_i } : 
                             (N4)? { io_resp_i[571:60], 1'b0, 1'b0, 1'b0, io_resp_i[43:4] } : 1'b0;
  assign N3 = lce_cmd_o_8_;
  assign N4 = lce_cmd_o[9];
  assign N5 = N24 | N26;
  assign N6 = N21 | N5;
  assign N7 = ~N6;
  assign lce_req_yumi_o = lce_req_v_i & io_cmd_ready_i;
  assign io_cmd_o[0] = N18;
  assign io_resp_yumi_o = io_resp_v_i & lce_cmd_ready_i;
  assign lce_cmd_o_8_ = N13;
  assign lce_cmd_o[9] = N12;

endmodule