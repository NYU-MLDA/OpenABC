module PTW( // @[:freechips.rocketchip.system.TinyConfig.fir@115493.2]
  output        io_requestor_0_pmp_0_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_0_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_0_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_0_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_0_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_0_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_0_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_1_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_1_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_1_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_1_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_1_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_1_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_1_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_2_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_2_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_2_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_2_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_2_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_2_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_2_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_3_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_3_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_3_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_3_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_3_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_3_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_3_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_4_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_4_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_4_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_4_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_4_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_4_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_4_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_5_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_5_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_5_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_5_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_5_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_5_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_5_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_6_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_6_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_6_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_6_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_6_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_6_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_6_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_7_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_0_pmp_7_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_7_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_7_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_0_pmp_7_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_0_pmp_7_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_0_pmp_7_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_0_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_0_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_0_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_0_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_0_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_0_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_0_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_1_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_1_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_1_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_1_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_1_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_1_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_1_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_2_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_2_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_2_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_2_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_2_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_2_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_2_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_3_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_3_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_3_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_3_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_3_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_3_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_3_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_4_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_4_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_4_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_4_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_4_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_4_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_4_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_5_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_5_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_5_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_5_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_5_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_5_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_5_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_6_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_6_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_6_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_6_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_6_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_6_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_6_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_7_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [1:0]  io_requestor_1_pmp_7_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_7_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_7_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output        io_requestor_1_pmp_7_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [29:0] io_requestor_1_pmp_7_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  output [31:0] io_requestor_1_pmp_7_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_0_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_0_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_0_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_0_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_0_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_0_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_0_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_1_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_1_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_1_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_1_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_1_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_1_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_1_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_2_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_2_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_2_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_2_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_2_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_2_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_2_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_3_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_3_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_3_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_3_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_3_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_3_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_3_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_4_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_4_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_4_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_4_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_4_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_4_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_4_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_5_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_5_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_5_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_5_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_5_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_5_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_5_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_6_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_6_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_6_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_6_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_6_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_6_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_6_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_7_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [1:0]  io_dpath_pmp_7_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_7_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_7_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input         io_dpath_pmp_7_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [29:0] io_dpath_pmp_7_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
  input  [31:0] io_dpath_pmp_7_mask // @[:freechips.rocketchip.system.TinyConfig.fir@115496.4]
);
  assign io_requestor_0_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_0_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116344.4]
  assign io_requestor_1_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
  assign io_requestor_1_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 277:25:freechips.rocketchip.system.TinyConfig.fir@116356.4]
endmodule