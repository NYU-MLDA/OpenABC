module bp_be_dcache_lce_tr_num_lce_p2_num_cce_p1_data_width_p64_paddr_width_p22_lce_data_width_p512_ways_p8_sets_p64
(
  tr_received_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_yumi_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [538:0] lce_tr_resp_i;
  output [521:0] data_mem_pkt_o;
  input lce_tr_resp_v_i;
  input data_mem_pkt_yumi_i;
  output tr_received_o;
  output lce_tr_resp_yumi_o;
  output data_mem_pkt_v_o;
  wire [521:0] data_mem_pkt_o;
  wire tr_received_o,lce_tr_resp_yumi_o,data_mem_pkt_v_o,data_mem_pkt_yumi_i,
  lce_tr_resp_v_i;
  assign data_mem_pkt_o[0] = 1'b1;
  assign tr_received_o = data_mem_pkt_yumi_i;
  assign lce_tr_resp_yumi_o = data_mem_pkt_yumi_i;
  assign data_mem_pkt_v_o = lce_tr_resp_v_i;
  assign data_mem_pkt_o[521] = lce_tr_resp_i[523];
  assign data_mem_pkt_o[520] = lce_tr_resp_i[522];
  assign data_mem_pkt_o[519] = lce_tr_resp_i[521];
  assign data_mem_pkt_o[518] = lce_tr_resp_i[520];
  assign data_mem_pkt_o[517] = lce_tr_resp_i[519];
  assign data_mem_pkt_o[516] = lce_tr_resp_i[518];
  assign data_mem_pkt_o[515] = lce_tr_resp_i[536];
  assign data_mem_pkt_o[514] = lce_tr_resp_i[535];
  assign data_mem_pkt_o[513] = lce_tr_resp_i[534];
  assign data_mem_pkt_o[512] = lce_tr_resp_i[511];
  assign data_mem_pkt_o[511] = lce_tr_resp_i[510];
  assign data_mem_pkt_o[510] = lce_tr_resp_i[509];
  assign data_mem_pkt_o[509] = lce_tr_resp_i[508];
  assign data_mem_pkt_o[508] = lce_tr_resp_i[507];
  assign data_mem_pkt_o[507] = lce_tr_resp_i[506];
  assign data_mem_pkt_o[506] = lce_tr_resp_i[505];
  assign data_mem_pkt_o[505] = lce_tr_resp_i[504];
  assign data_mem_pkt_o[504] = lce_tr_resp_i[503];
  assign data_mem_pkt_o[503] = lce_tr_resp_i[502];
  assign data_mem_pkt_o[502] = lce_tr_resp_i[501];
  assign data_mem_pkt_o[501] = lce_tr_resp_i[500];
  assign data_mem_pkt_o[500] = lce_tr_resp_i[499];
  assign data_mem_pkt_o[499] = lce_tr_resp_i[498];
  assign data_mem_pkt_o[498] = lce_tr_resp_i[497];
  assign data_mem_pkt_o[497] = lce_tr_resp_i[496];
  assign data_mem_pkt_o[496] = lce_tr_resp_i[495];
  assign data_mem_pkt_o[495] = lce_tr_resp_i[494];
  assign data_mem_pkt_o[494] = lce_tr_resp_i[493];
  assign data_mem_pkt_o[493] = lce_tr_resp_i[492];
  assign data_mem_pkt_o[492] = lce_tr_resp_i[491];
  assign data_mem_pkt_o[491] = lce_tr_resp_i[490];
  assign data_mem_pkt_o[490] = lce_tr_resp_i[489];
  assign data_mem_pkt_o[489] = lce_tr_resp_i[488];
  assign data_mem_pkt_o[488] = lce_tr_resp_i[487];
  assign data_mem_pkt_o[487] = lce_tr_resp_i[486];
  assign data_mem_pkt_o[486] = lce_tr_resp_i[485];
  assign data_mem_pkt_o[485] = lce_tr_resp_i[484];
  assign data_mem_pkt_o[484] = lce_tr_resp_i[483];
  assign data_mem_pkt_o[483] = lce_tr_resp_i[482];
  assign data_mem_pkt_o[482] = lce_tr_resp_i[481];
  assign data_mem_pkt_o[481] = lce_tr_resp_i[480];
  assign data_mem_pkt_o[480] = lce_tr_resp_i[479];
  assign data_mem_pkt_o[479] = lce_tr_resp_i[478];
  assign data_mem_pkt_o[478] = lce_tr_resp_i[477];
  assign data_mem_pkt_o[477] = lce_tr_resp_i[476];
  assign data_mem_pkt_o[476] = lce_tr_resp_i[475];
  assign data_mem_pkt_o[475] = lce_tr_resp_i[474];
  assign data_mem_pkt_o[474] = lce_tr_resp_i[473];
  assign data_mem_pkt_o[473] = lce_tr_resp_i[472];
  assign data_mem_pkt_o[472] = lce_tr_resp_i[471];
  assign data_mem_pkt_o[471] = lce_tr_resp_i[470];
  assign data_mem_pkt_o[470] = lce_tr_resp_i[469];
  assign data_mem_pkt_o[469] = lce_tr_resp_i[468];
  assign data_mem_pkt_o[468] = lce_tr_resp_i[467];
  assign data_mem_pkt_o[467] = lce_tr_resp_i[466];
  assign data_mem_pkt_o[466] = lce_tr_resp_i[465];
  assign data_mem_pkt_o[465] = lce_tr_resp_i[464];
  assign data_mem_pkt_o[464] = lce_tr_resp_i[463];
  assign data_mem_pkt_o[463] = lce_tr_resp_i[462];
  assign data_mem_pkt_o[462] = lce_tr_resp_i[461];
  assign data_mem_pkt_o[461] = lce_tr_resp_i[460];
  assign data_mem_pkt_o[460] = lce_tr_resp_i[459];
  assign data_mem_pkt_o[459] = lce_tr_resp_i[458];
  assign data_mem_pkt_o[458] = lce_tr_resp_i[457];
  assign data_mem_pkt_o[457] = lce_tr_resp_i[456];
  assign data_mem_pkt_o[456] = lce_tr_resp_i[455];
  assign data_mem_pkt_o[455] = lce_tr_resp_i[454];
  assign data_mem_pkt_o[454] = lce_tr_resp_i[453];
  assign data_mem_pkt_o[453] = lce_tr_resp_i[452];
  assign data_mem_pkt_o[452] = lce_tr_resp_i[451];
  assign data_mem_pkt_o[451] = lce_tr_resp_i[450];
  assign data_mem_pkt_o[450] = lce_tr_resp_i[449];
  assign data_mem_pkt_o[449] = lce_tr_resp_i[448];
  assign data_mem_pkt_o[448] = lce_tr_resp_i[447];
  assign data_mem_pkt_o[447] = lce_tr_resp_i[446];
  assign data_mem_pkt_o[446] = lce_tr_resp_i[445];
  assign data_mem_pkt_o[445] = lce_tr_resp_i[444];
  assign data_mem_pkt_o[444] = lce_tr_resp_i[443];
  assign data_mem_pkt_o[443] = lce_tr_resp_i[442];
  assign data_mem_pkt_o[442] = lce_tr_resp_i[441];
  assign data_mem_pkt_o[441] = lce_tr_resp_i[440];
  assign data_mem_pkt_o[440] = lce_tr_resp_i[439];
  assign data_mem_pkt_o[439] = lce_tr_resp_i[438];
  assign data_mem_pkt_o[438] = lce_tr_resp_i[437];
  assign data_mem_pkt_o[437] = lce_tr_resp_i[436];
  assign data_mem_pkt_o[436] = lce_tr_resp_i[435];
  assign data_mem_pkt_o[435] = lce_tr_resp_i[434];
  assign data_mem_pkt_o[434] = lce_tr_resp_i[433];
  assign data_mem_pkt_o[433] = lce_tr_resp_i[432];
  assign data_mem_pkt_o[432] = lce_tr_resp_i[431];
  assign data_mem_pkt_o[431] = lce_tr_resp_i[430];
  assign data_mem_pkt_o[430] = lce_tr_resp_i[429];
  assign data_mem_pkt_o[429] = lce_tr_resp_i[428];
  assign data_mem_pkt_o[428] = lce_tr_resp_i[427];
  assign data_mem_pkt_o[427] = lce_tr_resp_i[426];
  assign data_mem_pkt_o[426] = lce_tr_resp_i[425];
  assign data_mem_pkt_o[425] = lce_tr_resp_i[424];
  assign data_mem_pkt_o[424] = lce_tr_resp_i[423];
  assign data_mem_pkt_o[423] = lce_tr_resp_i[422];
  assign data_mem_pkt_o[422] = lce_tr_resp_i[421];
  assign data_mem_pkt_o[421] = lce_tr_resp_i[420];
  assign data_mem_pkt_o[420] = lce_tr_resp_i[419];
  assign data_mem_pkt_o[419] = lce_tr_resp_i[418];
  assign data_mem_pkt_o[418] = lce_tr_resp_i[417];
  assign data_mem_pkt_o[417] = lce_tr_resp_i[416];
  assign data_mem_pkt_o[416] = lce_tr_resp_i[415];
  assign data_mem_pkt_o[415] = lce_tr_resp_i[414];
  assign data_mem_pkt_o[414] = lce_tr_resp_i[413];
  assign data_mem_pkt_o[413] = lce_tr_resp_i[412];
  assign data_mem_pkt_o[412] = lce_tr_resp_i[411];
  assign data_mem_pkt_o[411] = lce_tr_resp_i[410];
  assign data_mem_pkt_o[410] = lce_tr_resp_i[409];
  assign data_mem_pkt_o[409] = lce_tr_resp_i[408];
  assign data_mem_pkt_o[408] = lce_tr_resp_i[407];
  assign data_mem_pkt_o[407] = lce_tr_resp_i[406];
  assign data_mem_pkt_o[406] = lce_tr_resp_i[405];
  assign data_mem_pkt_o[405] = lce_tr_resp_i[404];
  assign data_mem_pkt_o[404] = lce_tr_resp_i[403];
  assign data_mem_pkt_o[403] = lce_tr_resp_i[402];
  assign data_mem_pkt_o[402] = lce_tr_resp_i[401];
  assign data_mem_pkt_o[401] = lce_tr_resp_i[400];
  assign data_mem_pkt_o[400] = lce_tr_resp_i[399];
  assign data_mem_pkt_o[399] = lce_tr_resp_i[398];
  assign data_mem_pkt_o[398] = lce_tr_resp_i[397];
  assign data_mem_pkt_o[397] = lce_tr_resp_i[396];
  assign data_mem_pkt_o[396] = lce_tr_resp_i[395];
  assign data_mem_pkt_o[395] = lce_tr_resp_i[394];
  assign data_mem_pkt_o[394] = lce_tr_resp_i[393];
  assign data_mem_pkt_o[393] = lce_tr_resp_i[392];
  assign data_mem_pkt_o[392] = lce_tr_resp_i[391];
  assign data_mem_pkt_o[391] = lce_tr_resp_i[390];
  assign data_mem_pkt_o[390] = lce_tr_resp_i[389];
  assign data_mem_pkt_o[389] = lce_tr_resp_i[388];
  assign data_mem_pkt_o[388] = lce_tr_resp_i[387];
  assign data_mem_pkt_o[387] = lce_tr_resp_i[386];
  assign data_mem_pkt_o[386] = lce_tr_resp_i[385];
  assign data_mem_pkt_o[385] = lce_tr_resp_i[384];
  assign data_mem_pkt_o[384] = lce_tr_resp_i[383];
  assign data_mem_pkt_o[383] = lce_tr_resp_i[382];
  assign data_mem_pkt_o[382] = lce_tr_resp_i[381];
  assign data_mem_pkt_o[381] = lce_tr_resp_i[380];
  assign data_mem_pkt_o[380] = lce_tr_resp_i[379];
  assign data_mem_pkt_o[379] = lce_tr_resp_i[378];
  assign data_mem_pkt_o[378] = lce_tr_resp_i[377];
  assign data_mem_pkt_o[377] = lce_tr_resp_i[376];
  assign data_mem_pkt_o[376] = lce_tr_resp_i[375];
  assign data_mem_pkt_o[375] = lce_tr_resp_i[374];
  assign data_mem_pkt_o[374] = lce_tr_resp_i[373];
  assign data_mem_pkt_o[373] = lce_tr_resp_i[372];
  assign data_mem_pkt_o[372] = lce_tr_resp_i[371];
  assign data_mem_pkt_o[371] = lce_tr_resp_i[370];
  assign data_mem_pkt_o[370] = lce_tr_resp_i[369];
  assign data_mem_pkt_o[369] = lce_tr_resp_i[368];
  assign data_mem_pkt_o[368] = lce_tr_resp_i[367];
  assign data_mem_pkt_o[367] = lce_tr_resp_i[366];
  assign data_mem_pkt_o[366] = lce_tr_resp_i[365];
  assign data_mem_pkt_o[365] = lce_tr_resp_i[364];
  assign data_mem_pkt_o[364] = lce_tr_resp_i[363];
  assign data_mem_pkt_o[363] = lce_tr_resp_i[362];
  assign data_mem_pkt_o[362] = lce_tr_resp_i[361];
  assign data_mem_pkt_o[361] = lce_tr_resp_i[360];
  assign data_mem_pkt_o[360] = lce_tr_resp_i[359];
  assign data_mem_pkt_o[359] = lce_tr_resp_i[358];
  assign data_mem_pkt_o[358] = lce_tr_resp_i[357];
  assign data_mem_pkt_o[357] = lce_tr_resp_i[356];
  assign data_mem_pkt_o[356] = lce_tr_resp_i[355];
  assign data_mem_pkt_o[355] = lce_tr_resp_i[354];
  assign data_mem_pkt_o[354] = lce_tr_resp_i[353];
  assign data_mem_pkt_o[353] = lce_tr_resp_i[352];
  assign data_mem_pkt_o[352] = lce_tr_resp_i[351];
  assign data_mem_pkt_o[351] = lce_tr_resp_i[350];
  assign data_mem_pkt_o[350] = lce_tr_resp_i[349];
  assign data_mem_pkt_o[349] = lce_tr_resp_i[348];
  assign data_mem_pkt_o[348] = lce_tr_resp_i[347];
  assign data_mem_pkt_o[347] = lce_tr_resp_i[346];
  assign data_mem_pkt_o[346] = lce_tr_resp_i[345];
  assign data_mem_pkt_o[345] = lce_tr_resp_i[344];
  assign data_mem_pkt_o[344] = lce_tr_resp_i[343];
  assign data_mem_pkt_o[343] = lce_tr_resp_i[342];
  assign data_mem_pkt_o[342] = lce_tr_resp_i[341];
  assign data_mem_pkt_o[341] = lce_tr_resp_i[340];
  assign data_mem_pkt_o[340] = lce_tr_resp_i[339];
  assign data_mem_pkt_o[339] = lce_tr_resp_i[338];
  assign data_mem_pkt_o[338] = lce_tr_resp_i[337];
  assign data_mem_pkt_o[337] = lce_tr_resp_i[336];
  assign data_mem_pkt_o[336] = lce_tr_resp_i[335];
  assign data_mem_pkt_o[335] = lce_tr_resp_i[334];
  assign data_mem_pkt_o[334] = lce_tr_resp_i[333];
  assign data_mem_pkt_o[333] = lce_tr_resp_i[332];
  assign data_mem_pkt_o[332] = lce_tr_resp_i[331];
  assign data_mem_pkt_o[331] = lce_tr_resp_i[330];
  assign data_mem_pkt_o[330] = lce_tr_resp_i[329];
  assign data_mem_pkt_o[329] = lce_tr_resp_i[328];
  assign data_mem_pkt_o[328] = lce_tr_resp_i[327];
  assign data_mem_pkt_o[327] = lce_tr_resp_i[326];
  assign data_mem_pkt_o[326] = lce_tr_resp_i[325];
  assign data_mem_pkt_o[325] = lce_tr_resp_i[324];
  assign data_mem_pkt_o[324] = lce_tr_resp_i[323];
  assign data_mem_pkt_o[323] = lce_tr_resp_i[322];
  assign data_mem_pkt_o[322] = lce_tr_resp_i[321];
  assign data_mem_pkt_o[321] = lce_tr_resp_i[320];
  assign data_mem_pkt_o[320] = lce_tr_resp_i[319];
  assign data_mem_pkt_o[319] = lce_tr_resp_i[318];
  assign data_mem_pkt_o[318] = lce_tr_resp_i[317];
  assign data_mem_pkt_o[317] = lce_tr_resp_i[316];
  assign data_mem_pkt_o[316] = lce_tr_resp_i[315];
  assign data_mem_pkt_o[315] = lce_tr_resp_i[314];
  assign data_mem_pkt_o[314] = lce_tr_resp_i[313];
  assign data_mem_pkt_o[313] = lce_tr_resp_i[312];
  assign data_mem_pkt_o[312] = lce_tr_resp_i[311];
  assign data_mem_pkt_o[311] = lce_tr_resp_i[310];
  assign data_mem_pkt_o[310] = lce_tr_resp_i[309];
  assign data_mem_pkt_o[309] = lce_tr_resp_i[308];
  assign data_mem_pkt_o[308] = lce_tr_resp_i[307];
  assign data_mem_pkt_o[307] = lce_tr_resp_i[306];
  assign data_mem_pkt_o[306] = lce_tr_resp_i[305];
  assign data_mem_pkt_o[305] = lce_tr_resp_i[304];
  assign data_mem_pkt_o[304] = lce_tr_resp_i[303];
  assign data_mem_pkt_o[303] = lce_tr_resp_i[302];
  assign data_mem_pkt_o[302] = lce_tr_resp_i[301];
  assign data_mem_pkt_o[301] = lce_tr_resp_i[300];
  assign data_mem_pkt_o[300] = lce_tr_resp_i[299];
  assign data_mem_pkt_o[299] = lce_tr_resp_i[298];
  assign data_mem_pkt_o[298] = lce_tr_resp_i[297];
  assign data_mem_pkt_o[297] = lce_tr_resp_i[296];
  assign data_mem_pkt_o[296] = lce_tr_resp_i[295];
  assign data_mem_pkt_o[295] = lce_tr_resp_i[294];
  assign data_mem_pkt_o[294] = lce_tr_resp_i[293];
  assign data_mem_pkt_o[293] = lce_tr_resp_i[292];
  assign data_mem_pkt_o[292] = lce_tr_resp_i[291];
  assign data_mem_pkt_o[291] = lce_tr_resp_i[290];
  assign data_mem_pkt_o[290] = lce_tr_resp_i[289];
  assign data_mem_pkt_o[289] = lce_tr_resp_i[288];
  assign data_mem_pkt_o[288] = lce_tr_resp_i[287];
  assign data_mem_pkt_o[287] = lce_tr_resp_i[286];
  assign data_mem_pkt_o[286] = lce_tr_resp_i[285];
  assign data_mem_pkt_o[285] = lce_tr_resp_i[284];
  assign data_mem_pkt_o[284] = lce_tr_resp_i[283];
  assign data_mem_pkt_o[283] = lce_tr_resp_i[282];
  assign data_mem_pkt_o[282] = lce_tr_resp_i[281];
  assign data_mem_pkt_o[281] = lce_tr_resp_i[280];
  assign data_mem_pkt_o[280] = lce_tr_resp_i[279];
  assign data_mem_pkt_o[279] = lce_tr_resp_i[278];
  assign data_mem_pkt_o[278] = lce_tr_resp_i[277];
  assign data_mem_pkt_o[277] = lce_tr_resp_i[276];
  assign data_mem_pkt_o[276] = lce_tr_resp_i[275];
  assign data_mem_pkt_o[275] = lce_tr_resp_i[274];
  assign data_mem_pkt_o[274] = lce_tr_resp_i[273];
  assign data_mem_pkt_o[273] = lce_tr_resp_i[272];
  assign data_mem_pkt_o[272] = lce_tr_resp_i[271];
  assign data_mem_pkt_o[271] = lce_tr_resp_i[270];
  assign data_mem_pkt_o[270] = lce_tr_resp_i[269];
  assign data_mem_pkt_o[269] = lce_tr_resp_i[268];
  assign data_mem_pkt_o[268] = lce_tr_resp_i[267];
  assign data_mem_pkt_o[267] = lce_tr_resp_i[266];
  assign data_mem_pkt_o[266] = lce_tr_resp_i[265];
  assign data_mem_pkt_o[265] = lce_tr_resp_i[264];
  assign data_mem_pkt_o[264] = lce_tr_resp_i[263];
  assign data_mem_pkt_o[263] = lce_tr_resp_i[262];
  assign data_mem_pkt_o[262] = lce_tr_resp_i[261];
  assign data_mem_pkt_o[261] = lce_tr_resp_i[260];
  assign data_mem_pkt_o[260] = lce_tr_resp_i[259];
  assign data_mem_pkt_o[259] = lce_tr_resp_i[258];
  assign data_mem_pkt_o[258] = lce_tr_resp_i[257];
  assign data_mem_pkt_o[257] = lce_tr_resp_i[256];
  assign data_mem_pkt_o[256] = lce_tr_resp_i[255];
  assign data_mem_pkt_o[255] = lce_tr_resp_i[254];
  assign data_mem_pkt_o[254] = lce_tr_resp_i[253];
  assign data_mem_pkt_o[253] = lce_tr_resp_i[252];
  assign data_mem_pkt_o[252] = lce_tr_resp_i[251];
  assign data_mem_pkt_o[251] = lce_tr_resp_i[250];
  assign data_mem_pkt_o[250] = lce_tr_resp_i[249];
  assign data_mem_pkt_o[249] = lce_tr_resp_i[248];
  assign data_mem_pkt_o[248] = lce_tr_resp_i[247];
  assign data_mem_pkt_o[247] = lce_tr_resp_i[246];
  assign data_mem_pkt_o[246] = lce_tr_resp_i[245];
  assign data_mem_pkt_o[245] = lce_tr_resp_i[244];
  assign data_mem_pkt_o[244] = lce_tr_resp_i[243];
  assign data_mem_pkt_o[243] = lce_tr_resp_i[242];
  assign data_mem_pkt_o[242] = lce_tr_resp_i[241];
  assign data_mem_pkt_o[241] = lce_tr_resp_i[240];
  assign data_mem_pkt_o[240] = lce_tr_resp_i[239];
  assign data_mem_pkt_o[239] = lce_tr_resp_i[238];
  assign data_mem_pkt_o[238] = lce_tr_resp_i[237];
  assign data_mem_pkt_o[237] = lce_tr_resp_i[236];
  assign data_mem_pkt_o[236] = lce_tr_resp_i[235];
  assign data_mem_pkt_o[235] = lce_tr_resp_i[234];
  assign data_mem_pkt_o[234] = lce_tr_resp_i[233];
  assign data_mem_pkt_o[233] = lce_tr_resp_i[232];
  assign data_mem_pkt_o[232] = lce_tr_resp_i[231];
  assign data_mem_pkt_o[231] = lce_tr_resp_i[230];
  assign data_mem_pkt_o[230] = lce_tr_resp_i[229];
  assign data_mem_pkt_o[229] = lce_tr_resp_i[228];
  assign data_mem_pkt_o[228] = lce_tr_resp_i[227];
  assign data_mem_pkt_o[227] = lce_tr_resp_i[226];
  assign data_mem_pkt_o[226] = lce_tr_resp_i[225];
  assign data_mem_pkt_o[225] = lce_tr_resp_i[224];
  assign data_mem_pkt_o[224] = lce_tr_resp_i[223];
  assign data_mem_pkt_o[223] = lce_tr_resp_i[222];
  assign data_mem_pkt_o[222] = lce_tr_resp_i[221];
  assign data_mem_pkt_o[221] = lce_tr_resp_i[220];
  assign data_mem_pkt_o[220] = lce_tr_resp_i[219];
  assign data_mem_pkt_o[219] = lce_tr_resp_i[218];
  assign data_mem_pkt_o[218] = lce_tr_resp_i[217];
  assign data_mem_pkt_o[217] = lce_tr_resp_i[216];
  assign data_mem_pkt_o[216] = lce_tr_resp_i[215];
  assign data_mem_pkt_o[215] = lce_tr_resp_i[214];
  assign data_mem_pkt_o[214] = lce_tr_resp_i[213];
  assign data_mem_pkt_o[213] = lce_tr_resp_i[212];
  assign data_mem_pkt_o[212] = lce_tr_resp_i[211];
  assign data_mem_pkt_o[211] = lce_tr_resp_i[210];
  assign data_mem_pkt_o[210] = lce_tr_resp_i[209];
  assign data_mem_pkt_o[209] = lce_tr_resp_i[208];
  assign data_mem_pkt_o[208] = lce_tr_resp_i[207];
  assign data_mem_pkt_o[207] = lce_tr_resp_i[206];
  assign data_mem_pkt_o[206] = lce_tr_resp_i[205];
  assign data_mem_pkt_o[205] = lce_tr_resp_i[204];
  assign data_mem_pkt_o[204] = lce_tr_resp_i[203];
  assign data_mem_pkt_o[203] = lce_tr_resp_i[202];
  assign data_mem_pkt_o[202] = lce_tr_resp_i[201];
  assign data_mem_pkt_o[201] = lce_tr_resp_i[200];
  assign data_mem_pkt_o[200] = lce_tr_resp_i[199];
  assign data_mem_pkt_o[199] = lce_tr_resp_i[198];
  assign data_mem_pkt_o[198] = lce_tr_resp_i[197];
  assign data_mem_pkt_o[197] = lce_tr_resp_i[196];
  assign data_mem_pkt_o[196] = lce_tr_resp_i[195];
  assign data_mem_pkt_o[195] = lce_tr_resp_i[194];
  assign data_mem_pkt_o[194] = lce_tr_resp_i[193];
  assign data_mem_pkt_o[193] = lce_tr_resp_i[192];
  assign data_mem_pkt_o[192] = lce_tr_resp_i[191];
  assign data_mem_pkt_o[191] = lce_tr_resp_i[190];
  assign data_mem_pkt_o[190] = lce_tr_resp_i[189];
  assign data_mem_pkt_o[189] = lce_tr_resp_i[188];
  assign data_mem_pkt_o[188] = lce_tr_resp_i[187];
  assign data_mem_pkt_o[187] = lce_tr_resp_i[186];
  assign data_mem_pkt_o[186] = lce_tr_resp_i[185];
  assign data_mem_pkt_o[185] = lce_tr_resp_i[184];
  assign data_mem_pkt_o[184] = lce_tr_resp_i[183];
  assign data_mem_pkt_o[183] = lce_tr_resp_i[182];
  assign data_mem_pkt_o[182] = lce_tr_resp_i[181];
  assign data_mem_pkt_o[181] = lce_tr_resp_i[180];
  assign data_mem_pkt_o[180] = lce_tr_resp_i[179];
  assign data_mem_pkt_o[179] = lce_tr_resp_i[178];
  assign data_mem_pkt_o[178] = lce_tr_resp_i[177];
  assign data_mem_pkt_o[177] = lce_tr_resp_i[176];
  assign data_mem_pkt_o[176] = lce_tr_resp_i[175];
  assign data_mem_pkt_o[175] = lce_tr_resp_i[174];
  assign data_mem_pkt_o[174] = lce_tr_resp_i[173];
  assign data_mem_pkt_o[173] = lce_tr_resp_i[172];
  assign data_mem_pkt_o[172] = lce_tr_resp_i[171];
  assign data_mem_pkt_o[171] = lce_tr_resp_i[170];
  assign data_mem_pkt_o[170] = lce_tr_resp_i[169];
  assign data_mem_pkt_o[169] = lce_tr_resp_i[168];
  assign data_mem_pkt_o[168] = lce_tr_resp_i[167];
  assign data_mem_pkt_o[167] = lce_tr_resp_i[166];
  assign data_mem_pkt_o[166] = lce_tr_resp_i[165];
  assign data_mem_pkt_o[165] = lce_tr_resp_i[164];
  assign data_mem_pkt_o[164] = lce_tr_resp_i[163];
  assign data_mem_pkt_o[163] = lce_tr_resp_i[162];
  assign data_mem_pkt_o[162] = lce_tr_resp_i[161];
  assign data_mem_pkt_o[161] = lce_tr_resp_i[160];
  assign data_mem_pkt_o[160] = lce_tr_resp_i[159];
  assign data_mem_pkt_o[159] = lce_tr_resp_i[158];
  assign data_mem_pkt_o[158] = lce_tr_resp_i[157];
  assign data_mem_pkt_o[157] = lce_tr_resp_i[156];
  assign data_mem_pkt_o[156] = lce_tr_resp_i[155];
  assign data_mem_pkt_o[155] = lce_tr_resp_i[154];
  assign data_mem_pkt_o[154] = lce_tr_resp_i[153];
  assign data_mem_pkt_o[153] = lce_tr_resp_i[152];
  assign data_mem_pkt_o[152] = lce_tr_resp_i[151];
  assign data_mem_pkt_o[151] = lce_tr_resp_i[150];
  assign data_mem_pkt_o[150] = lce_tr_resp_i[149];
  assign data_mem_pkt_o[149] = lce_tr_resp_i[148];
  assign data_mem_pkt_o[148] = lce_tr_resp_i[147];
  assign data_mem_pkt_o[147] = lce_tr_resp_i[146];
  assign data_mem_pkt_o[146] = lce_tr_resp_i[145];
  assign data_mem_pkt_o[145] = lce_tr_resp_i[144];
  assign data_mem_pkt_o[144] = lce_tr_resp_i[143];
  assign data_mem_pkt_o[143] = lce_tr_resp_i[142];
  assign data_mem_pkt_o[142] = lce_tr_resp_i[141];
  assign data_mem_pkt_o[141] = lce_tr_resp_i[140];
  assign data_mem_pkt_o[140] = lce_tr_resp_i[139];
  assign data_mem_pkt_o[139] = lce_tr_resp_i[138];
  assign data_mem_pkt_o[138] = lce_tr_resp_i[137];
  assign data_mem_pkt_o[137] = lce_tr_resp_i[136];
  assign data_mem_pkt_o[136] = lce_tr_resp_i[135];
  assign data_mem_pkt_o[135] = lce_tr_resp_i[134];
  assign data_mem_pkt_o[134] = lce_tr_resp_i[133];
  assign data_mem_pkt_o[133] = lce_tr_resp_i[132];
  assign data_mem_pkt_o[132] = lce_tr_resp_i[131];
  assign data_mem_pkt_o[131] = lce_tr_resp_i[130];
  assign data_mem_pkt_o[130] = lce_tr_resp_i[129];
  assign data_mem_pkt_o[129] = lce_tr_resp_i[128];
  assign data_mem_pkt_o[128] = lce_tr_resp_i[127];
  assign data_mem_pkt_o[127] = lce_tr_resp_i[126];
  assign data_mem_pkt_o[126] = lce_tr_resp_i[125];
  assign data_mem_pkt_o[125] = lce_tr_resp_i[124];
  assign data_mem_pkt_o[124] = lce_tr_resp_i[123];
  assign data_mem_pkt_o[123] = lce_tr_resp_i[122];
  assign data_mem_pkt_o[122] = lce_tr_resp_i[121];
  assign data_mem_pkt_o[121] = lce_tr_resp_i[120];
  assign data_mem_pkt_o[120] = lce_tr_resp_i[119];
  assign data_mem_pkt_o[119] = lce_tr_resp_i[118];
  assign data_mem_pkt_o[118] = lce_tr_resp_i[117];
  assign data_mem_pkt_o[117] = lce_tr_resp_i[116];
  assign data_mem_pkt_o[116] = lce_tr_resp_i[115];
  assign data_mem_pkt_o[115] = lce_tr_resp_i[114];
  assign data_mem_pkt_o[114] = lce_tr_resp_i[113];
  assign data_mem_pkt_o[113] = lce_tr_resp_i[112];
  assign data_mem_pkt_o[112] = lce_tr_resp_i[111];
  assign data_mem_pkt_o[111] = lce_tr_resp_i[110];
  assign data_mem_pkt_o[110] = lce_tr_resp_i[109];
  assign data_mem_pkt_o[109] = lce_tr_resp_i[108];
  assign data_mem_pkt_o[108] = lce_tr_resp_i[107];
  assign data_mem_pkt_o[107] = lce_tr_resp_i[106];
  assign data_mem_pkt_o[106] = lce_tr_resp_i[105];
  assign data_mem_pkt_o[105] = lce_tr_resp_i[104];
  assign data_mem_pkt_o[104] = lce_tr_resp_i[103];
  assign data_mem_pkt_o[103] = lce_tr_resp_i[102];
  assign data_mem_pkt_o[102] = lce_tr_resp_i[101];
  assign data_mem_pkt_o[101] = lce_tr_resp_i[100];
  assign data_mem_pkt_o[100] = lce_tr_resp_i[99];
  assign data_mem_pkt_o[99] = lce_tr_resp_i[98];
  assign data_mem_pkt_o[98] = lce_tr_resp_i[97];
  assign data_mem_pkt_o[97] = lce_tr_resp_i[96];
  assign data_mem_pkt_o[96] = lce_tr_resp_i[95];
  assign data_mem_pkt_o[95] = lce_tr_resp_i[94];
  assign data_mem_pkt_o[94] = lce_tr_resp_i[93];
  assign data_mem_pkt_o[93] = lce_tr_resp_i[92];
  assign data_mem_pkt_o[92] = lce_tr_resp_i[91];
  assign data_mem_pkt_o[91] = lce_tr_resp_i[90];
  assign data_mem_pkt_o[90] = lce_tr_resp_i[89];
  assign data_mem_pkt_o[89] = lce_tr_resp_i[88];
  assign data_mem_pkt_o[88] = lce_tr_resp_i[87];
  assign data_mem_pkt_o[87] = lce_tr_resp_i[86];
  assign data_mem_pkt_o[86] = lce_tr_resp_i[85];
  assign data_mem_pkt_o[85] = lce_tr_resp_i[84];
  assign data_mem_pkt_o[84] = lce_tr_resp_i[83];
  assign data_mem_pkt_o[83] = lce_tr_resp_i[82];
  assign data_mem_pkt_o[82] = lce_tr_resp_i[81];
  assign data_mem_pkt_o[81] = lce_tr_resp_i[80];
  assign data_mem_pkt_o[80] = lce_tr_resp_i[79];
  assign data_mem_pkt_o[79] = lce_tr_resp_i[78];
  assign data_mem_pkt_o[78] = lce_tr_resp_i[77];
  assign data_mem_pkt_o[77] = lce_tr_resp_i[76];
  assign data_mem_pkt_o[76] = lce_tr_resp_i[75];
  assign data_mem_pkt_o[75] = lce_tr_resp_i[74];
  assign data_mem_pkt_o[74] = lce_tr_resp_i[73];
  assign data_mem_pkt_o[73] = lce_tr_resp_i[72];
  assign data_mem_pkt_o[72] = lce_tr_resp_i[71];
  assign data_mem_pkt_o[71] = lce_tr_resp_i[70];
  assign data_mem_pkt_o[70] = lce_tr_resp_i[69];
  assign data_mem_pkt_o[69] = lce_tr_resp_i[68];
  assign data_mem_pkt_o[68] = lce_tr_resp_i[67];
  assign data_mem_pkt_o[67] = lce_tr_resp_i[66];
  assign data_mem_pkt_o[66] = lce_tr_resp_i[65];
  assign data_mem_pkt_o[65] = lce_tr_resp_i[64];
  assign data_mem_pkt_o[64] = lce_tr_resp_i[63];
  assign data_mem_pkt_o[63] = lce_tr_resp_i[62];
  assign data_mem_pkt_o[62] = lce_tr_resp_i[61];
  assign data_mem_pkt_o[61] = lce_tr_resp_i[60];
  assign data_mem_pkt_o[60] = lce_tr_resp_i[59];
  assign data_mem_pkt_o[59] = lce_tr_resp_i[58];
  assign data_mem_pkt_o[58] = lce_tr_resp_i[57];
  assign data_mem_pkt_o[57] = lce_tr_resp_i[56];
  assign data_mem_pkt_o[56] = lce_tr_resp_i[55];
  assign data_mem_pkt_o[55] = lce_tr_resp_i[54];
  assign data_mem_pkt_o[54] = lce_tr_resp_i[53];
  assign data_mem_pkt_o[53] = lce_tr_resp_i[52];
  assign data_mem_pkt_o[52] = lce_tr_resp_i[51];
  assign data_mem_pkt_o[51] = lce_tr_resp_i[50];
  assign data_mem_pkt_o[50] = lce_tr_resp_i[49];
  assign data_mem_pkt_o[49] = lce_tr_resp_i[48];
  assign data_mem_pkt_o[48] = lce_tr_resp_i[47];
  assign data_mem_pkt_o[47] = lce_tr_resp_i[46];
  assign data_mem_pkt_o[46] = lce_tr_resp_i[45];
  assign data_mem_pkt_o[45] = lce_tr_resp_i[44];
  assign data_mem_pkt_o[44] = lce_tr_resp_i[43];
  assign data_mem_pkt_o[43] = lce_tr_resp_i[42];
  assign data_mem_pkt_o[42] = lce_tr_resp_i[41];
  assign data_mem_pkt_o[41] = lce_tr_resp_i[40];
  assign data_mem_pkt_o[40] = lce_tr_resp_i[39];
  assign data_mem_pkt_o[39] = lce_tr_resp_i[38];
  assign data_mem_pkt_o[38] = lce_tr_resp_i[37];
  assign data_mem_pkt_o[37] = lce_tr_resp_i[36];
  assign data_mem_pkt_o[36] = lce_tr_resp_i[35];
  assign data_mem_pkt_o[35] = lce_tr_resp_i[34];
  assign data_mem_pkt_o[34] = lce_tr_resp_i[33];
  assign data_mem_pkt_o[33] = lce_tr_resp_i[32];
  assign data_mem_pkt_o[32] = lce_tr_resp_i[31];
  assign data_mem_pkt_o[31] = lce_tr_resp_i[30];
  assign data_mem_pkt_o[30] = lce_tr_resp_i[29];
  assign data_mem_pkt_o[29] = lce_tr_resp_i[28];
  assign data_mem_pkt_o[28] = lce_tr_resp_i[27];
  assign data_mem_pkt_o[27] = lce_tr_resp_i[26];
  assign data_mem_pkt_o[26] = lce_tr_resp_i[25];
  assign data_mem_pkt_o[25] = lce_tr_resp_i[24];
  assign data_mem_pkt_o[24] = lce_tr_resp_i[23];
  assign data_mem_pkt_o[23] = lce_tr_resp_i[22];
  assign data_mem_pkt_o[22] = lce_tr_resp_i[21];
  assign data_mem_pkt_o[21] = lce_tr_resp_i[20];
  assign data_mem_pkt_o[20] = lce_tr_resp_i[19];
  assign data_mem_pkt_o[19] = lce_tr_resp_i[18];
  assign data_mem_pkt_o[18] = lce_tr_resp_i[17];
  assign data_mem_pkt_o[17] = lce_tr_resp_i[16];
  assign data_mem_pkt_o[16] = lce_tr_resp_i[15];
  assign data_mem_pkt_o[15] = lce_tr_resp_i[14];
  assign data_mem_pkt_o[14] = lce_tr_resp_i[13];
  assign data_mem_pkt_o[13] = lce_tr_resp_i[12];
  assign data_mem_pkt_o[12] = lce_tr_resp_i[11];
  assign data_mem_pkt_o[11] = lce_tr_resp_i[10];
  assign data_mem_pkt_o[10] = lce_tr_resp_i[9];
  assign data_mem_pkt_o[9] = lce_tr_resp_i[8];
  assign data_mem_pkt_o[8] = lce_tr_resp_i[7];
  assign data_mem_pkt_o[7] = lce_tr_resp_i[6];
  assign data_mem_pkt_o[6] = lce_tr_resp_i[5];
  assign data_mem_pkt_o[5] = lce_tr_resp_i[4];
  assign data_mem_pkt_o[4] = lce_tr_resp_i[3];
  assign data_mem_pkt_o[3] = lce_tr_resp_i[2];
  assign data_mem_pkt_o[2] = lce_tr_resp_i[1];
  assign data_mem_pkt_o[1] = lce_tr_resp_i[0];

endmodule