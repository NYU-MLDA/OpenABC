module rvbradder
(
  pc,
  offset,
  dout
);

  input [31:1] pc;
  input [12:1] offset;
  output [31:1] dout;
  wire [31:1] dout;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,cout,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153;
  wire [31:13] pc_inc,pc_dec;
  assign { cout, dout[12:1] } = pc[12:1] + offset;
  assign pc_inc = pc[31:13] + 1'b1;
  assign pc_dec = pc[31:13] - 1'b1;
  assign dout[31] = N24 | N27;
  assign N24 = N20 | N23;
  assign N20 = N19 & pc[31];
  assign N0 = offset[12] ^ cout;
  assign N19 = ~N0;
  assign N23 = N22 & pc_inc[31];
  assign N22 = N21 & cout;
  assign N21 = ~offset[12];
  assign N27 = N26 & pc_dec[31];
  assign N26 = offset[12] & N25;
  assign N25 = ~cout;
  assign dout[30] = N32 | N34;
  assign N32 = N29 | N31;
  assign N29 = N28 & pc[30];
  assign N1 = offset[12] ^ cout;
  assign N28 = ~N1;
  assign N31 = N30 & pc_inc[30];
  assign N30 = N21 & cout;
  assign N34 = N33 & pc_dec[30];
  assign N33 = offset[12] & N25;
  assign dout[29] = N39 | N41;
  assign N39 = N36 | N38;
  assign N36 = N35 & pc[29];
  assign N2 = offset[12] ^ cout;
  assign N35 = ~N2;
  assign N38 = N37 & pc_inc[29];
  assign N37 = N21 & cout;
  assign N41 = N40 & pc_dec[29];
  assign N40 = offset[12] & N25;
  assign dout[28] = N46 | N48;
  assign N46 = N43 | N45;
  assign N43 = N42 & pc[28];
  assign N3 = offset[12] ^ cout;
  assign N42 = ~N3;
  assign N45 = N44 & pc_inc[28];
  assign N44 = N21 & cout;
  assign N48 = N47 & pc_dec[28];
  assign N47 = offset[12] & N25;
  assign dout[27] = N53 | N55;
  assign N53 = N50 | N52;
  assign N50 = N49 & pc[27];
  assign N4 = offset[12] ^ cout;
  assign N49 = ~N4;
  assign N52 = N51 & pc_inc[27];
  assign N51 = N21 & cout;
  assign N55 = N54 & pc_dec[27];
  assign N54 = offset[12] & N25;
  assign dout[26] = N60 | N62;
  assign N60 = N57 | N59;
  assign N57 = N56 & pc[26];
  assign N5 = offset[12] ^ cout;
  assign N56 = ~N5;
  assign N59 = N58 & pc_inc[26];
  assign N58 = N21 & cout;
  assign N62 = N61 & pc_dec[26];
  assign N61 = offset[12] & N25;
  assign dout[25] = N67 | N69;
  assign N67 = N64 | N66;
  assign N64 = N63 & pc[25];
  assign N6 = offset[12] ^ cout;
  assign N63 = ~N6;
  assign N66 = N65 & pc_inc[25];
  assign N65 = N21 & cout;
  assign N69 = N68 & pc_dec[25];
  assign N68 = offset[12] & N25;
  assign dout[24] = N74 | N76;
  assign N74 = N71 | N73;
  assign N71 = N70 & pc[24];
  assign N7 = offset[12] ^ cout;
  assign N70 = ~N7;
  assign N73 = N72 & pc_inc[24];
  assign N72 = N21 & cout;
  assign N76 = N75 & pc_dec[24];
  assign N75 = offset[12] & N25;
  assign dout[23] = N81 | N83;
  assign N81 = N78 | N80;
  assign N78 = N77 & pc[23];
  assign N8 = offset[12] ^ cout;
  assign N77 = ~N8;
  assign N80 = N79 & pc_inc[23];
  assign N79 = N21 & cout;
  assign N83 = N82 & pc_dec[23];
  assign N82 = offset[12] & N25;
  assign dout[22] = N88 | N90;
  assign N88 = N85 | N87;
  assign N85 = N84 & pc[22];
  assign N9 = offset[12] ^ cout;
  assign N84 = ~N9;
  assign N87 = N86 & pc_inc[22];
  assign N86 = N21 & cout;
  assign N90 = N89 & pc_dec[22];
  assign N89 = offset[12] & N25;
  assign dout[21] = N95 | N97;
  assign N95 = N92 | N94;
  assign N92 = N91 & pc[21];
  assign N10 = offset[12] ^ cout;
  assign N91 = ~N10;
  assign N94 = N93 & pc_inc[21];
  assign N93 = N21 & cout;
  assign N97 = N96 & pc_dec[21];
  assign N96 = offset[12] & N25;
  assign dout[20] = N102 | N104;
  assign N102 = N99 | N101;
  assign N99 = N98 & pc[20];
  assign N11 = offset[12] ^ cout;
  assign N98 = ~N11;
  assign N101 = N100 & pc_inc[20];
  assign N100 = N21 & cout;
  assign N104 = N103 & pc_dec[20];
  assign N103 = offset[12] & N25;
  assign dout[19] = N109 | N111;
  assign N109 = N106 | N108;
  assign N106 = N105 & pc[19];
  assign N12 = offset[12] ^ cout;
  assign N105 = ~N12;
  assign N108 = N107 & pc_inc[19];
  assign N107 = N21 & cout;
  assign N111 = N110 & pc_dec[19];
  assign N110 = offset[12] & N25;
  assign dout[18] = N116 | N118;
  assign N116 = N113 | N115;
  assign N113 = N112 & pc[18];
  assign N13 = offset[12] ^ cout;
  assign N112 = ~N13;
  assign N115 = N114 & pc_inc[18];
  assign N114 = N21 & cout;
  assign N118 = N117 & pc_dec[18];
  assign N117 = offset[12] & N25;
  assign dout[17] = N123 | N125;
  assign N123 = N120 | N122;
  assign N120 = N119 & pc[17];
  assign N14 = offset[12] ^ cout;
  assign N119 = ~N14;
  assign N122 = N121 & pc_inc[17];
  assign N121 = N21 & cout;
  assign N125 = N124 & pc_dec[17];
  assign N124 = offset[12] & N25;
  assign dout[16] = N130 | N132;
  assign N130 = N127 | N129;
  assign N127 = N126 & pc[16];
  assign N15 = offset[12] ^ cout;
  assign N126 = ~N15;
  assign N129 = N128 & pc_inc[16];
  assign N128 = N21 & cout;
  assign N132 = N131 & pc_dec[16];
  assign N131 = offset[12] & N25;
  assign dout[15] = N137 | N139;
  assign N137 = N134 | N136;
  assign N134 = N133 & pc[15];
  assign N16 = offset[12] ^ cout;
  assign N133 = ~N16;
  assign N136 = N135 & pc_inc[15];
  assign N135 = N21 & cout;
  assign N139 = N138 & pc_dec[15];
  assign N138 = offset[12] & N25;
  assign dout[14] = N144 | N146;
  assign N144 = N141 | N143;
  assign N141 = N140 & pc[14];
  assign N17 = offset[12] ^ cout;
  assign N140 = ~N17;
  assign N143 = N142 & pc_inc[14];
  assign N142 = N21 & cout;
  assign N146 = N145 & pc_dec[14];
  assign N145 = offset[12] & N25;
  assign dout[13] = N151 | N153;
  assign N151 = N148 | N150;
  assign N148 = N147 & pc[13];
  assign N18 = offset[12] ^ cout;
  assign N147 = ~N18;
  assign N150 = N149 & pc_inc[13];
  assign N149 = N21 & cout;
  assign N153 = N152 & pc_dec[13];
  assign N152 = offset[12] & N25;

endmodule