module pipe_reg_simple_Depth0
(
  clk_i,
  rst_ni,
  d_i,
  d_o
);

  input [196:0] d_i;
  output [196:0] d_o;
  input clk_i;
  input rst_ni;
  wire [196:0] d_o;
  assign d_o[196] = d_i[196];
  assign d_o[195] = d_i[195];
  assign d_o[194] = d_i[194];
  assign d_o[193] = d_i[193];
  assign d_o[192] = d_i[192];
  assign d_o[191] = d_i[191];
  assign d_o[190] = d_i[190];
  assign d_o[189] = d_i[189];
  assign d_o[188] = d_i[188];
  assign d_o[187] = d_i[187];
  assign d_o[186] = d_i[186];
  assign d_o[185] = d_i[185];
  assign d_o[184] = d_i[184];
  assign d_o[183] = d_i[183];
  assign d_o[182] = d_i[182];
  assign d_o[181] = d_i[181];
  assign d_o[180] = d_i[180];
  assign d_o[179] = d_i[179];
  assign d_o[178] = d_i[178];
  assign d_o[177] = d_i[177];
  assign d_o[176] = d_i[176];
  assign d_o[175] = d_i[175];
  assign d_o[174] = d_i[174];
  assign d_o[173] = d_i[173];
  assign d_o[172] = d_i[172];
  assign d_o[171] = d_i[171];
  assign d_o[170] = d_i[170];
  assign d_o[169] = d_i[169];
  assign d_o[168] = d_i[168];
  assign d_o[167] = d_i[167];
  assign d_o[166] = d_i[166];
  assign d_o[165] = d_i[165];
  assign d_o[164] = d_i[164];
  assign d_o[163] = d_i[163];
  assign d_o[162] = d_i[162];
  assign d_o[161] = d_i[161];
  assign d_o[160] = d_i[160];
  assign d_o[159] = d_i[159];
  assign d_o[158] = d_i[158];
  assign d_o[157] = d_i[157];
  assign d_o[156] = d_i[156];
  assign d_o[155] = d_i[155];
  assign d_o[154] = d_i[154];
  assign d_o[153] = d_i[153];
  assign d_o[152] = d_i[152];
  assign d_o[151] = d_i[151];
  assign d_o[150] = d_i[150];
  assign d_o[149] = d_i[149];
  assign d_o[148] = d_i[148];
  assign d_o[147] = d_i[147];
  assign d_o[146] = d_i[146];
  assign d_o[145] = d_i[145];
  assign d_o[144] = d_i[144];
  assign d_o[143] = d_i[143];
  assign d_o[142] = d_i[142];
  assign d_o[141] = d_i[141];
  assign d_o[140] = d_i[140];
  assign d_o[139] = d_i[139];
  assign d_o[138] = d_i[138];
  assign d_o[137] = d_i[137];
  assign d_o[136] = d_i[136];
  assign d_o[135] = d_i[135];
  assign d_o[134] = d_i[134];
  assign d_o[133] = d_i[133];
  assign d_o[132] = d_i[132];
  assign d_o[131] = d_i[131];
  assign d_o[130] = d_i[130];
  assign d_o[129] = d_i[129];
  assign d_o[128] = d_i[128];
  assign d_o[127] = d_i[127];
  assign d_o[126] = d_i[126];
  assign d_o[125] = d_i[125];
  assign d_o[124] = d_i[124];
  assign d_o[123] = d_i[123];
  assign d_o[122] = d_i[122];
  assign d_o[121] = d_i[121];
  assign d_o[120] = d_i[120];
  assign d_o[119] = d_i[119];
  assign d_o[118] = d_i[118];
  assign d_o[117] = d_i[117];
  assign d_o[116] = d_i[116];
  assign d_o[115] = d_i[115];
  assign d_o[114] = d_i[114];
  assign d_o[113] = d_i[113];
  assign d_o[112] = d_i[112];
  assign d_o[111] = d_i[111];
  assign d_o[110] = d_i[110];
  assign d_o[109] = d_i[109];
  assign d_o[108] = d_i[108];
  assign d_o[107] = d_i[107];
  assign d_o[106] = d_i[106];
  assign d_o[105] = d_i[105];
  assign d_o[104] = d_i[104];
  assign d_o[103] = d_i[103];
  assign d_o[102] = d_i[102];
  assign d_o[101] = d_i[101];
  assign d_o[100] = d_i[100];
  assign d_o[99] = d_i[99];
  assign d_o[98] = d_i[98];
  assign d_o[97] = d_i[97];
  assign d_o[96] = d_i[96];
  assign d_o[95] = d_i[95];
  assign d_o[94] = d_i[94];
  assign d_o[93] = d_i[93];
  assign d_o[92] = d_i[92];
  assign d_o[91] = d_i[91];
  assign d_o[90] = d_i[90];
  assign d_o[89] = d_i[89];
  assign d_o[88] = d_i[88];
  assign d_o[87] = d_i[87];
  assign d_o[86] = d_i[86];
  assign d_o[85] = d_i[85];
  assign d_o[84] = d_i[84];
  assign d_o[83] = d_i[83];
  assign d_o[82] = d_i[82];
  assign d_o[81] = d_i[81];
  assign d_o[80] = d_i[80];
  assign d_o[79] = d_i[79];
  assign d_o[78] = d_i[78];
  assign d_o[77] = d_i[77];
  assign d_o[76] = d_i[76];
  assign d_o[75] = d_i[75];
  assign d_o[74] = d_i[74];
  assign d_o[73] = d_i[73];
  assign d_o[72] = d_i[72];
  assign d_o[71] = d_i[71];
  assign d_o[70] = d_i[70];
  assign d_o[69] = d_i[69];
  assign d_o[68] = d_i[68];
  assign d_o[67] = d_i[67];
  assign d_o[66] = d_i[66];
  assign d_o[65] = d_i[65];
  assign d_o[64] = d_i[64];
  assign d_o[63] = d_i[63];
  assign d_o[62] = d_i[62];
  assign d_o[61] = d_i[61];
  assign d_o[60] = d_i[60];
  assign d_o[59] = d_i[59];
  assign d_o[58] = d_i[58];
  assign d_o[57] = d_i[57];
  assign d_o[56] = d_i[56];
  assign d_o[55] = d_i[55];
  assign d_o[54] = d_i[54];
  assign d_o[53] = d_i[53];
  assign d_o[52] = d_i[52];
  assign d_o[51] = d_i[51];
  assign d_o[50] = d_i[50];
  assign d_o[49] = d_i[49];
  assign d_o[48] = d_i[48];
  assign d_o[47] = d_i[47];
  assign d_o[46] = d_i[46];
  assign d_o[45] = d_i[45];
  assign d_o[44] = d_i[44];
  assign d_o[43] = d_i[43];
  assign d_o[42] = d_i[42];
  assign d_o[41] = d_i[41];
  assign d_o[40] = d_i[40];
  assign d_o[39] = d_i[39];
  assign d_o[38] = d_i[38];
  assign d_o[37] = d_i[37];
  assign d_o[36] = d_i[36];
  assign d_o[35] = d_i[35];
  assign d_o[34] = d_i[34];
  assign d_o[33] = d_i[33];
  assign d_o[32] = d_i[32];
  assign d_o[31] = d_i[31];
  assign d_o[30] = d_i[30];
  assign d_o[29] = d_i[29];
  assign d_o[28] = d_i[28];
  assign d_o[27] = d_i[27];
  assign d_o[26] = d_i[26];
  assign d_o[25] = d_i[25];
  assign d_o[24] = d_i[24];
  assign d_o[23] = d_i[23];
  assign d_o[22] = d_i[22];
  assign d_o[21] = d_i[21];
  assign d_o[20] = d_i[20];
  assign d_o[19] = d_i[19];
  assign d_o[18] = d_i[18];
  assign d_o[17] = d_i[17];
  assign d_o[16] = d_i[16];
  assign d_o[15] = d_i[15];
  assign d_o[14] = d_i[14];
  assign d_o[13] = d_i[13];
  assign d_o[12] = d_i[12];
  assign d_o[11] = d_i[11];
  assign d_o[10] = d_i[10];
  assign d_o[9] = d_i[9];
  assign d_o[8] = d_i[8];
  assign d_o[7] = d_i[7];
  assign d_o[6] = d_i[6];
  assign d_o[5] = d_i[5];
  assign d_o[4] = d_i[4];
  assign d_o[3] = d_i[3];
  assign d_o[2] = d_i[2];
  assign d_o[1] = d_i[1];
  assign d_o[0] = d_i[0];

endmodule