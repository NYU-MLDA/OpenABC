module Htif
(
  clk,
  reset,
  io_host_in_ready,
  io_host_in_valid,
  io_host_in_bits,
  io_host_out_ready,
  io_host_out_valid,
  io_host_out_bits,
  io_host_debug_stats_csr,
  io_cpu_0_reset,
  io_cpu_0_id,
  io_cpu_0_csr_req_ready,
  io_cpu_0_csr_req_valid,
  io_cpu_0_csr_req_bits_rw,
  io_cpu_0_csr_req_bits_addr,
  io_cpu_0_csr_req_bits_data,
  io_cpu_0_csr_resp_ready,
  io_cpu_0_csr_resp_valid,
  io_cpu_0_csr_resp_bits,
  io_cpu_0_debug_stats_csr,
  io_mem_acquire_ready,
  io_mem_acquire_valid,
  io_mem_acquire_bits_addr_block,
  io_mem_acquire_bits_client_xact_id,
  io_mem_acquire_bits_addr_beat,
  io_mem_acquire_bits_is_builtin_type,
  io_mem_acquire_bits_a_type,
  io_mem_acquire_bits_union,
  io_mem_acquire_bits_data,
  io_mem_grant_ready,
  io_mem_grant_valid,
  io_mem_grant_bits_addr_beat,
  io_mem_grant_bits_client_xact_id,
  io_mem_grant_bits_manager_xact_id,
  io_mem_grant_bits_is_builtin_type,
  io_mem_grant_bits_g_type,
  io_mem_grant_bits_data,
  io_scr_req_ready,
  io_scr_req_valid,
  io_scr_req_bits_rw,
  io_scr_req_bits_addr,
  io_scr_req_bits_data,
  io_scr_resp_ready,
  io_scr_resp_valid,
  io_scr_resp_bits
);

  input [15:0] io_host_in_bits;
  output [15:0] io_host_out_bits;
  output [11:0] io_cpu_0_csr_req_bits_addr;
  output [63:0] io_cpu_0_csr_req_bits_data;
  input [63:0] io_cpu_0_csr_resp_bits;
  output [25:0] io_mem_acquire_bits_addr_block;
  output [5:0] io_mem_acquire_bits_client_xact_id;
  output [1:0] io_mem_acquire_bits_addr_beat;
  output [2:0] io_mem_acquire_bits_a_type;
  output [16:0] io_mem_acquire_bits_union;
  output [127:0] io_mem_acquire_bits_data;
  input [1:0] io_mem_grant_bits_addr_beat;
  input [5:0] io_mem_grant_bits_client_xact_id;
  input [3:0] io_mem_grant_bits_manager_xact_id;
  input [3:0] io_mem_grant_bits_g_type;
  input [127:0] io_mem_grant_bits_data;
  output [5:0] io_scr_req_bits_addr;
  output [63:0] io_scr_req_bits_data;
  input [63:0] io_scr_resp_bits;
  input clk;
  input reset;
  input io_host_in_valid;
  input io_host_out_ready;
  input io_cpu_0_csr_req_ready;
  input io_cpu_0_csr_resp_valid;
  input io_cpu_0_debug_stats_csr;
  input io_mem_acquire_ready;
  input io_mem_grant_valid;
  input io_mem_grant_bits_is_builtin_type;
  input io_scr_req_ready;
  input io_scr_resp_valid;
  output io_host_in_ready;
  output io_host_out_valid;
  output io_host_debug_stats_csr;
  output io_cpu_0_reset;
  output io_cpu_0_id;
  output io_cpu_0_csr_req_valid;
  output io_cpu_0_csr_req_bits_rw;
  output io_cpu_0_csr_resp_ready;
  output io_mem_acquire_valid;
  output io_mem_acquire_bits_is_builtin_type;
  output io_mem_grant_ready;
  output io_scr_req_valid;
  output io_scr_req_bits_rw;
  output io_scr_resp_ready;
  wire [15:0] io_host_out_bits;
  wire [63:0] io_cpu_0_csr_req_bits_data,tx_data,T195,T196;
  wire [5:0] io_mem_acquire_bits_client_xact_id;
  wire [1:0] io_mem_acquire_bits_addr_beat,T82;
  wire [2:0] io_mem_acquire_bits_a_type,T15,T16,packet_ram_raddr,T142;
  wire [16:0] io_mem_acquire_bits_union;
  wire [127:0] io_mem_acquire_bits_data,T152;
  wire io_host_in_ready,io_host_out_valid,io_host_debug_stats_csr,io_cpu_0_id,
  io_cpu_0_csr_req_valid,io_cpu_0_csr_req_bits_rw,io_cpu_0_csr_resp_ready,
  io_mem_acquire_valid,io_mem_acquire_bits_is_builtin_type,io_mem_grant_ready,io_scr_req_valid,
  io_scr_req_bits_rw,io_scr_resp_ready,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,io_cpu_0_debug_stats_csr,T2,T132,T131,T129,
  T124,T123,T113,T107,T101,T89,T79,T66,T18,N63,T21,T61,T26,T27,T32,N64,T38,T33,T35,
  nack,T54,N65,bad_mem_packet,T39,T41,N66,T60,rx_done,rx_word_done,T67,T72,T68,T71,
  cnt_done,T83,T86,T84,T92,T104,T110,tx_done,T120,T114,T119,T115,T118,T116,T126,
  T137,T141,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,T185,T190,tx_header_0,T200,N95,N96,N97,
  N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,
  N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
  N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,
  N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,
  N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,
  N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,
  N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,
  N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
  N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,
  N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,
  N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,
  N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
  N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,
  N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,
  N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,
  N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,
  N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,
  N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,
  N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,
  N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,
  N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,
  N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,
  N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
  N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
  N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,
  N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,
  N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
  N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,
  N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,
  N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,
  N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,
  N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,
  N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,
  N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,
  N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,
  N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,
  N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
  N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,
  N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,
  N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,
  N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,
  N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,
  N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,
  N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,
  N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,
  N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,
  N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,
  N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,
  N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,
  N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,
  N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,
  N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,
  N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,
  N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,
  N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,
  N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,
  N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,
  N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,
  N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,
  N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,
  N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,
  N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,
  N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,
  N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,
  N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,
  N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,
  N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,
  N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,
  N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,
  N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,
  N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,
  N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,
  N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,
  N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,
  N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,
  N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,
  N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,
  N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,
  N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,
  N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,
  N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,
  N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,
  N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,
  N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,
  N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,
  N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,
  N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,
  N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,
  N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,
  N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,
  N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,
  N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,
  N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,
  N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,
  N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,
  N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,
  N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,
  N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,
  N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,
  N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,
  N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,
  N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,
  N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,
  N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,
  N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,
  N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,
  N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,
  N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,
  N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,
  N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,
  N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,
  N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,
  N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,
  N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,
  N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,
  N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,
  N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,
  N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,
  N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,
  N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,
  N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,
  N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,
  N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,
  N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,
  N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,
  N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,
  N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,
  N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,
  N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,
  N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,
  N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,
  N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,
  N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,
  N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,
  N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,
  N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,
  N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,
  N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,
  N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,
  N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,
  N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,
  N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,
  N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,
  N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,
  N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
  N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,
  N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,
  N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,
  N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,
  N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,
  N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,
  N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,
  N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,
  N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,
  N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,
  N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,
  N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,
  N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,
  N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,
  N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,
  N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,
  N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,
  N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,
  N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,
  N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2510,N2511,N2512,N2514,N2515,N2516,
  N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,
  N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,
  N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,
  N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,
  N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,
  N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,
  N2597,N2598,N2599,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,
  N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,N2651,
  N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,
  N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
  N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,N2691,
  N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,N2705,
  N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,
  N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,
  N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
  N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,
  N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,N2771,
  N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785,
  N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  io_cpu_0_id_snps_wire,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,
  SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11,SV2V_UNCONNECTED_12,SV2V_UNCONNECTED_13,
  SV2V_UNCONNECTED_14,SV2V_UNCONNECTED_15,SV2V_UNCONNECTED_16,
  SV2V_UNCONNECTED_17,SV2V_UNCONNECTED_18,SV2V_UNCONNECTED_19,
  SV2V_UNCONNECTED_20,SV2V_UNCONNECTED_21,SV2V_UNCONNECTED_22,SV2V_UNCONNECTED_23,
  SV2V_UNCONNECTED_24,SV2V_UNCONNECTED_25,SV2V_UNCONNECTED_26,
  SV2V_UNCONNECTED_27,SV2V_UNCONNECTED_28,SV2V_UNCONNECTED_29,
  SV2V_UNCONNECTED_30,SV2V_UNCONNECTED_31,SV2V_UNCONNECTED_32,SV2V_UNCONNECTED_33,
  SV2V_UNCONNECTED_34,SV2V_UNCONNECTED_35,SV2V_UNCONNECTED_36,
  SV2V_UNCONNECTED_37,SV2V_UNCONNECTED_38,SV2V_UNCONNECTED_39,
  SV2V_UNCONNECTED_40,SV2V_UNCONNECTED_41,SV2V_UNCONNECTED_42,SV2V_UNCONNECTED_43,
  SV2V_UNCONNECTED_44,SV2V_UNCONNECTED_45,SV2V_UNCONNECTED_46,
  SV2V_UNCONNECTED_47,SV2V_UNCONNECTED_48;
  wire [1:1] T109;
  wire [2:2] T103,T91,T17;
  wire [3:0] rx_cmd;
  wire [14:0] T25,T59;
  wire [11:0] T212;
  wire [39:0] T51,T50;
  wire [8:0] T99,T98;
  reg packet_ram_7__63_,packet_ram_7__62_,packet_ram_7__61_,packet_ram_7__60_,
  packet_ram_7__59_,packet_ram_7__58_,packet_ram_7__57_,packet_ram_7__56_,
  packet_ram_7__55_,packet_ram_7__54_,packet_ram_7__53_,packet_ram_7__52_,packet_ram_7__51_,
  packet_ram_7__50_,packet_ram_7__49_,packet_ram_7__48_,packet_ram_7__47_,
  packet_ram_7__46_,packet_ram_7__45_,packet_ram_7__44_,packet_ram_7__43_,packet_ram_7__42_,
  packet_ram_7__41_,packet_ram_7__40_,packet_ram_7__39_,packet_ram_7__38_,
  packet_ram_7__37_,packet_ram_7__36_,packet_ram_7__35_,packet_ram_7__34_,packet_ram_7__33_,
  packet_ram_7__32_,packet_ram_7__31_,packet_ram_7__30_,packet_ram_7__29_,
  packet_ram_7__28_,packet_ram_7__27_,packet_ram_7__26_,packet_ram_7__25_,packet_ram_7__24_,
  packet_ram_7__23_,packet_ram_7__22_,packet_ram_7__21_,packet_ram_7__20_,
  packet_ram_7__19_,packet_ram_7__18_,packet_ram_7__17_,packet_ram_7__16_,
  packet_ram_7__15_,packet_ram_7__14_,packet_ram_7__13_,packet_ram_7__12_,packet_ram_7__11_,
  packet_ram_7__10_,packet_ram_7__9_,packet_ram_7__8_,packet_ram_7__7_,packet_ram_7__6_,
  packet_ram_7__5_,packet_ram_7__4_,packet_ram_7__3_,packet_ram_7__2_,
  packet_ram_7__1_,packet_ram_7__0_,packet_ram_6__63_,packet_ram_6__62_,packet_ram_6__61_,
  packet_ram_6__60_,packet_ram_6__59_,packet_ram_6__58_,packet_ram_6__57_,
  packet_ram_6__56_,packet_ram_6__55_,packet_ram_6__54_,packet_ram_6__53_,packet_ram_6__52_,
  packet_ram_6__51_,packet_ram_6__50_,packet_ram_6__49_,packet_ram_6__48_,
  packet_ram_6__47_,packet_ram_6__46_,packet_ram_6__45_,packet_ram_6__44_,packet_ram_6__43_,
  packet_ram_6__42_,packet_ram_6__41_,packet_ram_6__40_,packet_ram_6__39_,
  packet_ram_6__38_,packet_ram_6__37_,packet_ram_6__36_,packet_ram_6__35_,
  packet_ram_6__34_,packet_ram_6__33_,packet_ram_6__32_,packet_ram_6__31_,packet_ram_6__30_,
  packet_ram_6__29_,packet_ram_6__28_,packet_ram_6__27_,packet_ram_6__26_,
  packet_ram_6__25_,packet_ram_6__24_,packet_ram_6__23_,packet_ram_6__22_,packet_ram_6__21_,
  packet_ram_6__20_,packet_ram_6__19_,packet_ram_6__18_,packet_ram_6__17_,
  packet_ram_6__16_,packet_ram_6__15_,packet_ram_6__14_,packet_ram_6__13_,packet_ram_6__12_,
  packet_ram_6__11_,packet_ram_6__10_,packet_ram_6__9_,packet_ram_6__8_,
  packet_ram_6__7_,packet_ram_6__6_,packet_ram_6__5_,packet_ram_6__4_,packet_ram_6__3_,
  packet_ram_6__2_,packet_ram_6__1_,packet_ram_6__0_,packet_ram_5__63_,packet_ram_5__62_,
  packet_ram_5__61_,packet_ram_5__60_,packet_ram_5__59_,packet_ram_5__58_,
  packet_ram_5__57_,packet_ram_5__56_,packet_ram_5__55_,packet_ram_5__54_,
  packet_ram_5__53_,packet_ram_5__52_,packet_ram_5__51_,packet_ram_5__50_,packet_ram_5__49_,
  packet_ram_5__48_,packet_ram_5__47_,packet_ram_5__46_,packet_ram_5__45_,
  packet_ram_5__44_,packet_ram_5__43_,packet_ram_5__42_,packet_ram_5__41_,packet_ram_5__40_,
  packet_ram_5__39_,packet_ram_5__38_,packet_ram_5__37_,packet_ram_5__36_,
  packet_ram_5__35_,packet_ram_5__34_,packet_ram_5__33_,packet_ram_5__32_,packet_ram_5__31_,
  packet_ram_5__30_,packet_ram_5__29_,packet_ram_5__28_,packet_ram_5__27_,
  packet_ram_5__26_,packet_ram_5__25_,packet_ram_5__24_,packet_ram_5__23_,packet_ram_5__22_,
  packet_ram_5__21_,packet_ram_5__20_,packet_ram_5__19_,packet_ram_5__18_,
  packet_ram_5__17_,packet_ram_5__16_,packet_ram_5__15_,packet_ram_5__14_,
  packet_ram_5__13_,packet_ram_5__12_,packet_ram_5__11_,packet_ram_5__10_,packet_ram_5__9_,
  packet_ram_5__8_,packet_ram_5__7_,packet_ram_5__6_,packet_ram_5__5_,packet_ram_5__4_,
  packet_ram_5__3_,packet_ram_5__2_,packet_ram_5__1_,packet_ram_5__0_,
  packet_ram_4__63_,packet_ram_4__62_,packet_ram_4__61_,packet_ram_4__60_,packet_ram_4__59_,
  packet_ram_4__58_,packet_ram_4__57_,packet_ram_4__56_,packet_ram_4__55_,
  packet_ram_4__54_,packet_ram_4__53_,packet_ram_4__52_,packet_ram_4__51_,packet_ram_4__50_,
  packet_ram_4__49_,packet_ram_4__48_,packet_ram_4__47_,packet_ram_4__46_,
  packet_ram_4__45_,packet_ram_4__44_,packet_ram_4__43_,packet_ram_4__42_,packet_ram_4__41_,
  packet_ram_4__40_,packet_ram_4__39_,packet_ram_4__38_,packet_ram_4__37_,
  packet_ram_4__36_,packet_ram_4__35_,packet_ram_4__34_,packet_ram_4__33_,
  packet_ram_4__32_,packet_ram_4__31_,packet_ram_4__30_,packet_ram_4__29_,packet_ram_4__28_,
  packet_ram_4__27_,packet_ram_4__26_,packet_ram_4__25_,packet_ram_4__24_,
  packet_ram_4__23_,packet_ram_4__22_,packet_ram_4__21_,packet_ram_4__20_,packet_ram_4__19_,
  packet_ram_4__18_,packet_ram_4__17_,packet_ram_4__16_,packet_ram_4__15_,
  packet_ram_4__14_,packet_ram_4__13_,packet_ram_4__12_,packet_ram_4__11_,packet_ram_4__10_,
  packet_ram_4__9_,packet_ram_4__8_,packet_ram_4__7_,packet_ram_4__6_,
  packet_ram_4__5_,packet_ram_4__4_,packet_ram_4__3_,packet_ram_4__2_,packet_ram_4__1_,
  packet_ram_4__0_,packet_ram_3__63_,packet_ram_3__62_,packet_ram_3__61_,packet_ram_3__60_,
  packet_ram_3__59_,packet_ram_3__58_,packet_ram_3__57_,packet_ram_3__56_,
  packet_ram_3__55_,packet_ram_3__54_,packet_ram_3__53_,packet_ram_3__52_,
  packet_ram_3__51_,packet_ram_3__50_,packet_ram_3__49_,packet_ram_3__48_,packet_ram_3__47_,
  packet_ram_3__46_,packet_ram_3__45_,packet_ram_3__44_,packet_ram_3__43_,
  packet_ram_3__42_,packet_ram_3__41_,packet_ram_3__40_,packet_ram_3__39_,packet_ram_3__38_,
  packet_ram_3__37_,packet_ram_3__36_,packet_ram_3__35_,packet_ram_3__34_,
  packet_ram_3__33_,packet_ram_3__32_,packet_ram_3__31_,packet_ram_3__30_,packet_ram_3__29_,
  packet_ram_3__28_,packet_ram_3__27_,packet_ram_3__26_,packet_ram_3__25_,
  packet_ram_3__24_,packet_ram_3__23_,packet_ram_3__22_,packet_ram_3__21_,packet_ram_3__20_,
  packet_ram_3__19_,packet_ram_3__18_,packet_ram_3__17_,packet_ram_3__16_,
  packet_ram_3__15_,packet_ram_3__14_,packet_ram_3__13_,packet_ram_3__12_,
  packet_ram_3__11_,packet_ram_3__10_,packet_ram_3__9_,packet_ram_3__8_,packet_ram_3__7_,
  packet_ram_3__6_,packet_ram_3__5_,packet_ram_3__4_,packet_ram_3__3_,packet_ram_3__2_,
  packet_ram_3__1_,packet_ram_3__0_,packet_ram_2__63_,packet_ram_2__62_,
  packet_ram_2__61_,packet_ram_2__60_,packet_ram_2__59_,packet_ram_2__58_,packet_ram_2__57_,
  packet_ram_2__56_,packet_ram_2__55_,packet_ram_2__54_,packet_ram_2__53_,
  packet_ram_2__52_,packet_ram_2__51_,packet_ram_2__50_,packet_ram_2__49_,packet_ram_2__48_,
  packet_ram_2__47_,packet_ram_2__46_,packet_ram_2__45_,packet_ram_2__44_,
  packet_ram_2__43_,packet_ram_2__42_,packet_ram_2__41_,packet_ram_2__40_,packet_ram_2__39_,
  packet_ram_2__38_,packet_ram_2__37_,packet_ram_2__36_,packet_ram_2__35_,
  packet_ram_2__34_,packet_ram_2__33_,packet_ram_2__32_,packet_ram_2__31_,
  packet_ram_2__30_,packet_ram_2__29_,packet_ram_2__28_,packet_ram_2__27_,packet_ram_2__26_,
  packet_ram_2__25_,packet_ram_2__24_,packet_ram_2__23_,packet_ram_2__22_,
  packet_ram_2__21_,packet_ram_2__20_,packet_ram_2__19_,packet_ram_2__18_,packet_ram_2__17_,
  packet_ram_2__16_,packet_ram_2__15_,packet_ram_2__14_,packet_ram_2__13_,
  packet_ram_2__12_,packet_ram_2__11_,packet_ram_2__10_,packet_ram_2__9_,packet_ram_2__8_,
  packet_ram_2__7_,packet_ram_2__6_,packet_ram_2__5_,packet_ram_2__4_,
  packet_ram_2__3_,packet_ram_2__2_,packet_ram_2__1_,packet_ram_2__0_,packet_ram_1__63_,
  packet_ram_1__62_,packet_ram_1__61_,packet_ram_1__60_,packet_ram_1__59_,packet_ram_1__58_,
  packet_ram_1__57_,packet_ram_1__56_,packet_ram_1__55_,packet_ram_1__54_,
  packet_ram_1__53_,packet_ram_1__52_,packet_ram_1__51_,packet_ram_1__50_,
  packet_ram_1__49_,packet_ram_1__48_,packet_ram_1__47_,packet_ram_1__46_,packet_ram_1__45_,
  packet_ram_1__44_,packet_ram_1__43_,packet_ram_1__42_,packet_ram_1__41_,
  packet_ram_1__40_,packet_ram_1__39_,packet_ram_1__38_,packet_ram_1__37_,packet_ram_1__36_,
  packet_ram_1__35_,packet_ram_1__34_,packet_ram_1__33_,packet_ram_1__32_,
  packet_ram_1__31_,packet_ram_1__30_,packet_ram_1__29_,packet_ram_1__28_,packet_ram_1__27_,
  packet_ram_1__26_,packet_ram_1__25_,packet_ram_1__24_,packet_ram_1__23_,
  packet_ram_1__22_,packet_ram_1__21_,packet_ram_1__20_,packet_ram_1__19_,packet_ram_1__18_,
  packet_ram_1__17_,packet_ram_1__16_,packet_ram_1__15_,packet_ram_1__14_,
  packet_ram_1__13_,packet_ram_1__12_,packet_ram_1__11_,packet_ram_1__10_,
  packet_ram_1__9_,packet_ram_1__8_,packet_ram_1__7_,packet_ram_1__6_,packet_ram_1__5_,
  packet_ram_1__4_,packet_ram_1__3_,packet_ram_1__2_,packet_ram_1__1_,packet_ram_1__0_,
  rx_shifter_in_3,rx_shifter_in_2,rx_shifter_in_1,rx_shifter_in_0,io_cpu_0_reset;
  reg [63:0] io_scr_req_bits_data,csrReadData;
  reg [2:0] state,T53;
  reg [3:0] cmd;
  reg [12:0] rx_word_count,tx_word_count;
  reg [1:0] T77,tx_subword_count;
  reg [11:3] T214;
  reg [47:16] rx_shifter_in;
  reg [11:0] T29,io_cpu_0_csr_req_bits_addr;
  reg [36:26] init_addr;
  reg [25:0] io_mem_acquire_bits_addr_block;
  reg [5:0] io_scr_req_bits_addr;
  reg [2:1] T154;
  reg [8:0] pos;
  reg [23:16] tx_header;
  assign io_mem_acquire_bits_is_builtin_type = 1'b1;
  assign io_mem_acquire_bits_a_type[0] = 1'b1;
  assign io_mem_acquire_bits_union[8] = 1'b1;
  assign io_mem_acquire_bits_union[7] = 1'b1;
  assign io_mem_acquire_bits_union[6] = 1'b1;
  assign io_mem_acquire_bits_union[0] = 1'b1;
  assign io_cpu_0_csr_resp_ready = 1'b1;
  assign io_mem_grant_ready = 1'b1;
  assign io_scr_resp_ready = 1'b1;
  assign io_mem_acquire_bits_client_xact_id[5] = 1'b0;
  assign io_mem_acquire_bits_client_xact_id[4] = 1'b0;
  assign io_mem_acquire_bits_client_xact_id[3] = 1'b0;
  assign io_mem_acquire_bits_client_xact_id[2] = 1'b0;
  assign io_mem_acquire_bits_client_xact_id[1] = 1'b0;
  assign io_mem_acquire_bits_client_xact_id[0] = 1'b0;
  assign io_mem_acquire_bits_a_type[2] = 1'b0;
  assign io_mem_acquire_bits_union[1] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[2] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[3] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[4] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[5] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[9] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[10] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[11] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[12] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[13] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[14] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[15] = io_mem_acquire_bits_a_type[1];
  assign io_mem_acquire_bits_union[16] = io_mem_acquire_bits_a_type[1];
  assign io_host_debug_stats_csr = io_cpu_0_debug_stats_csr;
  assign io_mem_acquire_bits_addr_block[8] = io_cpu_0_csr_req_bits_addr[11];
  assign io_mem_acquire_bits_addr_block[7] = io_cpu_0_csr_req_bits_addr[10];
  assign io_mem_acquire_bits_addr_block[6] = io_cpu_0_csr_req_bits_addr[9];
  assign io_mem_acquire_bits_addr_block[5] = io_cpu_0_csr_req_bits_addr[8];
  assign io_mem_acquire_bits_addr_block[4] = io_cpu_0_csr_req_bits_addr[7];
  assign io_mem_acquire_bits_addr_block[3] = io_cpu_0_csr_req_bits_addr[6];
  assign io_mem_acquire_bits_addr_block[2] = io_scr_req_bits_addr[5];
  assign io_cpu_0_csr_req_bits_addr[5] = io_scr_req_bits_addr[5];
  assign io_mem_acquire_bits_addr_block[1] = io_scr_req_bits_addr[4];
  assign io_cpu_0_csr_req_bits_addr[4] = io_scr_req_bits_addr[4];
  assign io_mem_acquire_bits_addr_block[0] = io_scr_req_bits_addr[3];
  assign io_cpu_0_csr_req_bits_addr[3] = io_scr_req_bits_addr[3];
  assign io_cpu_0_csr_req_bits_addr[2] = io_scr_req_bits_addr[2];
  assign io_cpu_0_csr_req_bits_addr[1] = io_scr_req_bits_addr[1];
  assign io_cpu_0_csr_req_bits_addr[0] = io_scr_req_bits_addr[0];
  assign io_cpu_0_csr_req_bits_data[63] = io_scr_req_bits_data[63];
  assign io_cpu_0_csr_req_bits_data[62] = io_scr_req_bits_data[62];
  assign io_cpu_0_csr_req_bits_data[61] = io_scr_req_bits_data[61];
  assign io_cpu_0_csr_req_bits_data[60] = io_scr_req_bits_data[60];
  assign io_cpu_0_csr_req_bits_data[59] = io_scr_req_bits_data[59];
  assign io_cpu_0_csr_req_bits_data[58] = io_scr_req_bits_data[58];
  assign io_cpu_0_csr_req_bits_data[57] = io_scr_req_bits_data[57];
  assign io_cpu_0_csr_req_bits_data[56] = io_scr_req_bits_data[56];
  assign io_cpu_0_csr_req_bits_data[55] = io_scr_req_bits_data[55];
  assign io_cpu_0_csr_req_bits_data[54] = io_scr_req_bits_data[54];
  assign io_cpu_0_csr_req_bits_data[53] = io_scr_req_bits_data[53];
  assign io_cpu_0_csr_req_bits_data[52] = io_scr_req_bits_data[52];
  assign io_cpu_0_csr_req_bits_data[51] = io_scr_req_bits_data[51];
  assign io_cpu_0_csr_req_bits_data[50] = io_scr_req_bits_data[50];
  assign io_cpu_0_csr_req_bits_data[49] = io_scr_req_bits_data[49];
  assign io_cpu_0_csr_req_bits_data[48] = io_scr_req_bits_data[48];
  assign io_cpu_0_csr_req_bits_data[47] = io_scr_req_bits_data[47];
  assign io_cpu_0_csr_req_bits_data[46] = io_scr_req_bits_data[46];
  assign io_cpu_0_csr_req_bits_data[45] = io_scr_req_bits_data[45];
  assign io_cpu_0_csr_req_bits_data[44] = io_scr_req_bits_data[44];
  assign io_cpu_0_csr_req_bits_data[43] = io_scr_req_bits_data[43];
  assign io_cpu_0_csr_req_bits_data[42] = io_scr_req_bits_data[42];
  assign io_cpu_0_csr_req_bits_data[41] = io_scr_req_bits_data[41];
  assign io_cpu_0_csr_req_bits_data[40] = io_scr_req_bits_data[40];
  assign io_cpu_0_csr_req_bits_data[39] = io_scr_req_bits_data[39];
  assign io_cpu_0_csr_req_bits_data[38] = io_scr_req_bits_data[38];
  assign io_cpu_0_csr_req_bits_data[37] = io_scr_req_bits_data[37];
  assign io_cpu_0_csr_req_bits_data[36] = io_scr_req_bits_data[36];
  assign io_cpu_0_csr_req_bits_data[35] = io_scr_req_bits_data[35];
  assign io_cpu_0_csr_req_bits_data[34] = io_scr_req_bits_data[34];
  assign io_cpu_0_csr_req_bits_data[33] = io_scr_req_bits_data[33];
  assign io_cpu_0_csr_req_bits_data[32] = io_scr_req_bits_data[32];
  assign io_cpu_0_csr_req_bits_data[31] = io_scr_req_bits_data[31];
  assign io_cpu_0_csr_req_bits_data[30] = io_scr_req_bits_data[30];
  assign io_cpu_0_csr_req_bits_data[29] = io_scr_req_bits_data[29];
  assign io_cpu_0_csr_req_bits_data[28] = io_scr_req_bits_data[28];
  assign io_cpu_0_csr_req_bits_data[27] = io_scr_req_bits_data[27];
  assign io_cpu_0_csr_req_bits_data[26] = io_scr_req_bits_data[26];
  assign io_cpu_0_csr_req_bits_data[25] = io_scr_req_bits_data[25];
  assign io_cpu_0_csr_req_bits_data[24] = io_scr_req_bits_data[24];
  assign io_cpu_0_csr_req_bits_data[23] = io_scr_req_bits_data[23];
  assign io_cpu_0_csr_req_bits_data[22] = io_scr_req_bits_data[22];
  assign io_cpu_0_csr_req_bits_data[21] = io_scr_req_bits_data[21];
  assign io_cpu_0_csr_req_bits_data[20] = io_scr_req_bits_data[20];
  assign io_cpu_0_csr_req_bits_data[19] = io_scr_req_bits_data[19];
  assign io_cpu_0_csr_req_bits_data[18] = io_scr_req_bits_data[18];
  assign io_cpu_0_csr_req_bits_data[17] = io_scr_req_bits_data[17];
  assign io_cpu_0_csr_req_bits_data[16] = io_scr_req_bits_data[16];
  assign io_cpu_0_csr_req_bits_data[15] = io_scr_req_bits_data[15];
  assign io_cpu_0_csr_req_bits_data[14] = io_scr_req_bits_data[14];
  assign io_cpu_0_csr_req_bits_data[13] = io_scr_req_bits_data[13];
  assign io_cpu_0_csr_req_bits_data[12] = io_scr_req_bits_data[12];
  assign io_cpu_0_csr_req_bits_data[11] = io_scr_req_bits_data[11];
  assign io_cpu_0_csr_req_bits_data[10] = io_scr_req_bits_data[10];
  assign io_cpu_0_csr_req_bits_data[9] = io_scr_req_bits_data[9];
  assign io_cpu_0_csr_req_bits_data[8] = io_scr_req_bits_data[8];
  assign io_cpu_0_csr_req_bits_data[7] = io_scr_req_bits_data[7];
  assign io_cpu_0_csr_req_bits_data[6] = io_scr_req_bits_data[6];
  assign io_cpu_0_csr_req_bits_data[5] = io_scr_req_bits_data[5];
  assign io_cpu_0_csr_req_bits_data[4] = io_scr_req_bits_data[4];
  assign io_cpu_0_csr_req_bits_data[3] = io_scr_req_bits_data[3];
  assign io_cpu_0_csr_req_bits_data[2] = io_scr_req_bits_data[2];
  assign io_cpu_0_csr_req_bits_data[1] = io_scr_req_bits_data[1];
  assign io_cpu_0_csr_req_bits_data[0] = io_scr_req_bits_data[0];
  assign T27 = tx_word_count == { 1'b0, T212 };
  assign T71 = rx_word_count == { 1'b0, T214, T53 };
  assign T116 = packet_ram_raddr == { 1'b1, 1'b1, 1'b1 };
  assign T118 = 1'b0 < tx_word_count;
  assign T119 = tx_word_count == { 1'b0, T212 };
  assign T152[63] = (N74)? io_scr_req_bits_data[63] : 
                    (N76)? packet_ram_1__63_ : 
                    (N78)? packet_ram_2__63_ : 
                    (N80)? packet_ram_3__63_ : 
                    (N75)? packet_ram_4__63_ : 
                    (N77)? packet_ram_5__63_ : 
                    (N79)? packet_ram_6__63_ : 
                    (N81)? packet_ram_7__63_ : 1'b0;
  assign T152[62] = (N74)? io_scr_req_bits_data[62] : 
                    (N76)? packet_ram_1__62_ : 
                    (N78)? packet_ram_2__62_ : 
                    (N80)? packet_ram_3__62_ : 
                    (N75)? packet_ram_4__62_ : 
                    (N77)? packet_ram_5__62_ : 
                    (N79)? packet_ram_6__62_ : 
                    (N81)? packet_ram_7__62_ : 1'b0;
  assign T152[61] = (N74)? io_scr_req_bits_data[61] : 
                    (N76)? packet_ram_1__61_ : 
                    (N78)? packet_ram_2__61_ : 
                    (N80)? packet_ram_3__61_ : 
                    (N75)? packet_ram_4__61_ : 
                    (N77)? packet_ram_5__61_ : 
                    (N79)? packet_ram_6__61_ : 
                    (N81)? packet_ram_7__61_ : 1'b0;
  assign T152[60] = (N74)? io_scr_req_bits_data[60] : 
                    (N76)? packet_ram_1__60_ : 
                    (N78)? packet_ram_2__60_ : 
                    (N80)? packet_ram_3__60_ : 
                    (N75)? packet_ram_4__60_ : 
                    (N77)? packet_ram_5__60_ : 
                    (N79)? packet_ram_6__60_ : 
                    (N81)? packet_ram_7__60_ : 1'b0;
  assign T152[59] = (N74)? io_scr_req_bits_data[59] : 
                    (N76)? packet_ram_1__59_ : 
                    (N78)? packet_ram_2__59_ : 
                    (N80)? packet_ram_3__59_ : 
                    (N75)? packet_ram_4__59_ : 
                    (N77)? packet_ram_5__59_ : 
                    (N79)? packet_ram_6__59_ : 
                    (N81)? packet_ram_7__59_ : 1'b0;
  assign T152[58] = (N74)? io_scr_req_bits_data[58] : 
                    (N76)? packet_ram_1__58_ : 
                    (N78)? packet_ram_2__58_ : 
                    (N80)? packet_ram_3__58_ : 
                    (N75)? packet_ram_4__58_ : 
                    (N77)? packet_ram_5__58_ : 
                    (N79)? packet_ram_6__58_ : 
                    (N81)? packet_ram_7__58_ : 1'b0;
  assign T152[57] = (N74)? io_scr_req_bits_data[57] : 
                    (N76)? packet_ram_1__57_ : 
                    (N78)? packet_ram_2__57_ : 
                    (N80)? packet_ram_3__57_ : 
                    (N75)? packet_ram_4__57_ : 
                    (N77)? packet_ram_5__57_ : 
                    (N79)? packet_ram_6__57_ : 
                    (N81)? packet_ram_7__57_ : 1'b0;
  assign T152[56] = (N74)? io_scr_req_bits_data[56] : 
                    (N76)? packet_ram_1__56_ : 
                    (N78)? packet_ram_2__56_ : 
                    (N80)? packet_ram_3__56_ : 
                    (N75)? packet_ram_4__56_ : 
                    (N77)? packet_ram_5__56_ : 
                    (N79)? packet_ram_6__56_ : 
                    (N81)? packet_ram_7__56_ : 1'b0;
  assign T152[55] = (N74)? io_scr_req_bits_data[55] : 
                    (N76)? packet_ram_1__55_ : 
                    (N78)? packet_ram_2__55_ : 
                    (N80)? packet_ram_3__55_ : 
                    (N75)? packet_ram_4__55_ : 
                    (N77)? packet_ram_5__55_ : 
                    (N79)? packet_ram_6__55_ : 
                    (N81)? packet_ram_7__55_ : 1'b0;
  assign T152[54] = (N74)? io_scr_req_bits_data[54] : 
                    (N76)? packet_ram_1__54_ : 
                    (N78)? packet_ram_2__54_ : 
                    (N80)? packet_ram_3__54_ : 
                    (N75)? packet_ram_4__54_ : 
                    (N77)? packet_ram_5__54_ : 
                    (N79)? packet_ram_6__54_ : 
                    (N81)? packet_ram_7__54_ : 1'b0;
  assign T152[53] = (N74)? io_scr_req_bits_data[53] : 
                    (N76)? packet_ram_1__53_ : 
                    (N78)? packet_ram_2__53_ : 
                    (N80)? packet_ram_3__53_ : 
                    (N75)? packet_ram_4__53_ : 
                    (N77)? packet_ram_5__53_ : 
                    (N79)? packet_ram_6__53_ : 
                    (N81)? packet_ram_7__53_ : 1'b0;
  assign T152[52] = (N74)? io_scr_req_bits_data[52] : 
                    (N76)? packet_ram_1__52_ : 
                    (N78)? packet_ram_2__52_ : 
                    (N80)? packet_ram_3__52_ : 
                    (N75)? packet_ram_4__52_ : 
                    (N77)? packet_ram_5__52_ : 
                    (N79)? packet_ram_6__52_ : 
                    (N81)? packet_ram_7__52_ : 1'b0;
  assign T152[51] = (N74)? io_scr_req_bits_data[51] : 
                    (N76)? packet_ram_1__51_ : 
                    (N78)? packet_ram_2__51_ : 
                    (N80)? packet_ram_3__51_ : 
                    (N75)? packet_ram_4__51_ : 
                    (N77)? packet_ram_5__51_ : 
                    (N79)? packet_ram_6__51_ : 
                    (N81)? packet_ram_7__51_ : 1'b0;
  assign T152[50] = (N74)? io_scr_req_bits_data[50] : 
                    (N76)? packet_ram_1__50_ : 
                    (N78)? packet_ram_2__50_ : 
                    (N80)? packet_ram_3__50_ : 
                    (N75)? packet_ram_4__50_ : 
                    (N77)? packet_ram_5__50_ : 
                    (N79)? packet_ram_6__50_ : 
                    (N81)? packet_ram_7__50_ : 1'b0;
  assign T152[49] = (N74)? io_scr_req_bits_data[49] : 
                    (N76)? packet_ram_1__49_ : 
                    (N78)? packet_ram_2__49_ : 
                    (N80)? packet_ram_3__49_ : 
                    (N75)? packet_ram_4__49_ : 
                    (N77)? packet_ram_5__49_ : 
                    (N79)? packet_ram_6__49_ : 
                    (N81)? packet_ram_7__49_ : 1'b0;
  assign T152[48] = (N74)? io_scr_req_bits_data[48] : 
                    (N76)? packet_ram_1__48_ : 
                    (N78)? packet_ram_2__48_ : 
                    (N80)? packet_ram_3__48_ : 
                    (N75)? packet_ram_4__48_ : 
                    (N77)? packet_ram_5__48_ : 
                    (N79)? packet_ram_6__48_ : 
                    (N81)? packet_ram_7__48_ : 1'b0;
  assign T152[47] = (N74)? io_scr_req_bits_data[47] : 
                    (N76)? packet_ram_1__47_ : 
                    (N78)? packet_ram_2__47_ : 
                    (N80)? packet_ram_3__47_ : 
                    (N75)? packet_ram_4__47_ : 
                    (N77)? packet_ram_5__47_ : 
                    (N79)? packet_ram_6__47_ : 
                    (N81)? packet_ram_7__47_ : 1'b0;
  assign T152[46] = (N74)? io_scr_req_bits_data[46] : 
                    (N76)? packet_ram_1__46_ : 
                    (N78)? packet_ram_2__46_ : 
                    (N80)? packet_ram_3__46_ : 
                    (N75)? packet_ram_4__46_ : 
                    (N77)? packet_ram_5__46_ : 
                    (N79)? packet_ram_6__46_ : 
                    (N81)? packet_ram_7__46_ : 1'b0;
  assign T152[45] = (N74)? io_scr_req_bits_data[45] : 
                    (N76)? packet_ram_1__45_ : 
                    (N78)? packet_ram_2__45_ : 
                    (N80)? packet_ram_3__45_ : 
                    (N75)? packet_ram_4__45_ : 
                    (N77)? packet_ram_5__45_ : 
                    (N79)? packet_ram_6__45_ : 
                    (N81)? packet_ram_7__45_ : 1'b0;
  assign T152[44] = (N74)? io_scr_req_bits_data[44] : 
                    (N76)? packet_ram_1__44_ : 
                    (N78)? packet_ram_2__44_ : 
                    (N80)? packet_ram_3__44_ : 
                    (N75)? packet_ram_4__44_ : 
                    (N77)? packet_ram_5__44_ : 
                    (N79)? packet_ram_6__44_ : 
                    (N81)? packet_ram_7__44_ : 1'b0;
  assign T152[43] = (N74)? io_scr_req_bits_data[43] : 
                    (N76)? packet_ram_1__43_ : 
                    (N78)? packet_ram_2__43_ : 
                    (N80)? packet_ram_3__43_ : 
                    (N75)? packet_ram_4__43_ : 
                    (N77)? packet_ram_5__43_ : 
                    (N79)? packet_ram_6__43_ : 
                    (N81)? packet_ram_7__43_ : 1'b0;
  assign T152[42] = (N74)? io_scr_req_bits_data[42] : 
                    (N76)? packet_ram_1__42_ : 
                    (N78)? packet_ram_2__42_ : 
                    (N80)? packet_ram_3__42_ : 
                    (N75)? packet_ram_4__42_ : 
                    (N77)? packet_ram_5__42_ : 
                    (N79)? packet_ram_6__42_ : 
                    (N81)? packet_ram_7__42_ : 1'b0;
  assign T152[41] = (N74)? io_scr_req_bits_data[41] : 
                    (N76)? packet_ram_1__41_ : 
                    (N78)? packet_ram_2__41_ : 
                    (N80)? packet_ram_3__41_ : 
                    (N75)? packet_ram_4__41_ : 
                    (N77)? packet_ram_5__41_ : 
                    (N79)? packet_ram_6__41_ : 
                    (N81)? packet_ram_7__41_ : 1'b0;
  assign T152[40] = (N74)? io_scr_req_bits_data[40] : 
                    (N76)? packet_ram_1__40_ : 
                    (N78)? packet_ram_2__40_ : 
                    (N80)? packet_ram_3__40_ : 
                    (N75)? packet_ram_4__40_ : 
                    (N77)? packet_ram_5__40_ : 
                    (N79)? packet_ram_6__40_ : 
                    (N81)? packet_ram_7__40_ : 1'b0;
  assign T152[39] = (N74)? io_scr_req_bits_data[39] : 
                    (N76)? packet_ram_1__39_ : 
                    (N78)? packet_ram_2__39_ : 
                    (N80)? packet_ram_3__39_ : 
                    (N75)? packet_ram_4__39_ : 
                    (N77)? packet_ram_5__39_ : 
                    (N79)? packet_ram_6__39_ : 
                    (N81)? packet_ram_7__39_ : 1'b0;
  assign T152[38] = (N74)? io_scr_req_bits_data[38] : 
                    (N76)? packet_ram_1__38_ : 
                    (N78)? packet_ram_2__38_ : 
                    (N80)? packet_ram_3__38_ : 
                    (N75)? packet_ram_4__38_ : 
                    (N77)? packet_ram_5__38_ : 
                    (N79)? packet_ram_6__38_ : 
                    (N81)? packet_ram_7__38_ : 1'b0;
  assign T152[37] = (N74)? io_scr_req_bits_data[37] : 
                    (N76)? packet_ram_1__37_ : 
                    (N78)? packet_ram_2__37_ : 
                    (N80)? packet_ram_3__37_ : 
                    (N75)? packet_ram_4__37_ : 
                    (N77)? packet_ram_5__37_ : 
                    (N79)? packet_ram_6__37_ : 
                    (N81)? packet_ram_7__37_ : 1'b0;
  assign T152[36] = (N74)? io_scr_req_bits_data[36] : 
                    (N76)? packet_ram_1__36_ : 
                    (N78)? packet_ram_2__36_ : 
                    (N80)? packet_ram_3__36_ : 
                    (N75)? packet_ram_4__36_ : 
                    (N77)? packet_ram_5__36_ : 
                    (N79)? packet_ram_6__36_ : 
                    (N81)? packet_ram_7__36_ : 1'b0;
  assign T152[35] = (N74)? io_scr_req_bits_data[35] : 
                    (N76)? packet_ram_1__35_ : 
                    (N78)? packet_ram_2__35_ : 
                    (N80)? packet_ram_3__35_ : 
                    (N75)? packet_ram_4__35_ : 
                    (N77)? packet_ram_5__35_ : 
                    (N79)? packet_ram_6__35_ : 
                    (N81)? packet_ram_7__35_ : 1'b0;
  assign T152[34] = (N74)? io_scr_req_bits_data[34] : 
                    (N76)? packet_ram_1__34_ : 
                    (N78)? packet_ram_2__34_ : 
                    (N80)? packet_ram_3__34_ : 
                    (N75)? packet_ram_4__34_ : 
                    (N77)? packet_ram_5__34_ : 
                    (N79)? packet_ram_6__34_ : 
                    (N81)? packet_ram_7__34_ : 1'b0;
  assign T152[33] = (N74)? io_scr_req_bits_data[33] : 
                    (N76)? packet_ram_1__33_ : 
                    (N78)? packet_ram_2__33_ : 
                    (N80)? packet_ram_3__33_ : 
                    (N75)? packet_ram_4__33_ : 
                    (N77)? packet_ram_5__33_ : 
                    (N79)? packet_ram_6__33_ : 
                    (N81)? packet_ram_7__33_ : 1'b0;
  assign T152[32] = (N74)? io_scr_req_bits_data[32] : 
                    (N76)? packet_ram_1__32_ : 
                    (N78)? packet_ram_2__32_ : 
                    (N80)? packet_ram_3__32_ : 
                    (N75)? packet_ram_4__32_ : 
                    (N77)? packet_ram_5__32_ : 
                    (N79)? packet_ram_6__32_ : 
                    (N81)? packet_ram_7__32_ : 1'b0;
  assign T152[31] = (N74)? io_scr_req_bits_data[31] : 
                    (N76)? packet_ram_1__31_ : 
                    (N78)? packet_ram_2__31_ : 
                    (N80)? packet_ram_3__31_ : 
                    (N75)? packet_ram_4__31_ : 
                    (N77)? packet_ram_5__31_ : 
                    (N79)? packet_ram_6__31_ : 
                    (N81)? packet_ram_7__31_ : 1'b0;
  assign T152[30] = (N74)? io_scr_req_bits_data[30] : 
                    (N76)? packet_ram_1__30_ : 
                    (N78)? packet_ram_2__30_ : 
                    (N80)? packet_ram_3__30_ : 
                    (N75)? packet_ram_4__30_ : 
                    (N77)? packet_ram_5__30_ : 
                    (N79)? packet_ram_6__30_ : 
                    (N81)? packet_ram_7__30_ : 1'b0;
  assign T152[29] = (N74)? io_scr_req_bits_data[29] : 
                    (N76)? packet_ram_1__29_ : 
                    (N78)? packet_ram_2__29_ : 
                    (N80)? packet_ram_3__29_ : 
                    (N75)? packet_ram_4__29_ : 
                    (N77)? packet_ram_5__29_ : 
                    (N79)? packet_ram_6__29_ : 
                    (N81)? packet_ram_7__29_ : 1'b0;
  assign T152[28] = (N74)? io_scr_req_bits_data[28] : 
                    (N76)? packet_ram_1__28_ : 
                    (N78)? packet_ram_2__28_ : 
                    (N80)? packet_ram_3__28_ : 
                    (N75)? packet_ram_4__28_ : 
                    (N77)? packet_ram_5__28_ : 
                    (N79)? packet_ram_6__28_ : 
                    (N81)? packet_ram_7__28_ : 1'b0;
  assign T152[27] = (N74)? io_scr_req_bits_data[27] : 
                    (N76)? packet_ram_1__27_ : 
                    (N78)? packet_ram_2__27_ : 
                    (N80)? packet_ram_3__27_ : 
                    (N75)? packet_ram_4__27_ : 
                    (N77)? packet_ram_5__27_ : 
                    (N79)? packet_ram_6__27_ : 
                    (N81)? packet_ram_7__27_ : 1'b0;
  assign T152[26] = (N74)? io_scr_req_bits_data[26] : 
                    (N76)? packet_ram_1__26_ : 
                    (N78)? packet_ram_2__26_ : 
                    (N80)? packet_ram_3__26_ : 
                    (N75)? packet_ram_4__26_ : 
                    (N77)? packet_ram_5__26_ : 
                    (N79)? packet_ram_6__26_ : 
                    (N81)? packet_ram_7__26_ : 1'b0;
  assign T152[25] = (N74)? io_scr_req_bits_data[25] : 
                    (N76)? packet_ram_1__25_ : 
                    (N78)? packet_ram_2__25_ : 
                    (N80)? packet_ram_3__25_ : 
                    (N75)? packet_ram_4__25_ : 
                    (N77)? packet_ram_5__25_ : 
                    (N79)? packet_ram_6__25_ : 
                    (N81)? packet_ram_7__25_ : 1'b0;
  assign T152[24] = (N74)? io_scr_req_bits_data[24] : 
                    (N76)? packet_ram_1__24_ : 
                    (N78)? packet_ram_2__24_ : 
                    (N80)? packet_ram_3__24_ : 
                    (N75)? packet_ram_4__24_ : 
                    (N77)? packet_ram_5__24_ : 
                    (N79)? packet_ram_6__24_ : 
                    (N81)? packet_ram_7__24_ : 1'b0;
  assign T152[23] = (N74)? io_scr_req_bits_data[23] : 
                    (N76)? packet_ram_1__23_ : 
                    (N78)? packet_ram_2__23_ : 
                    (N80)? packet_ram_3__23_ : 
                    (N75)? packet_ram_4__23_ : 
                    (N77)? packet_ram_5__23_ : 
                    (N79)? packet_ram_6__23_ : 
                    (N81)? packet_ram_7__23_ : 1'b0;
  assign T152[22] = (N74)? io_scr_req_bits_data[22] : 
                    (N76)? packet_ram_1__22_ : 
                    (N78)? packet_ram_2__22_ : 
                    (N80)? packet_ram_3__22_ : 
                    (N75)? packet_ram_4__22_ : 
                    (N77)? packet_ram_5__22_ : 
                    (N79)? packet_ram_6__22_ : 
                    (N81)? packet_ram_7__22_ : 1'b0;
  assign T152[21] = (N74)? io_scr_req_bits_data[21] : 
                    (N76)? packet_ram_1__21_ : 
                    (N78)? packet_ram_2__21_ : 
                    (N80)? packet_ram_3__21_ : 
                    (N75)? packet_ram_4__21_ : 
                    (N77)? packet_ram_5__21_ : 
                    (N79)? packet_ram_6__21_ : 
                    (N81)? packet_ram_7__21_ : 1'b0;
  assign T152[20] = (N74)? io_scr_req_bits_data[20] : 
                    (N76)? packet_ram_1__20_ : 
                    (N78)? packet_ram_2__20_ : 
                    (N80)? packet_ram_3__20_ : 
                    (N75)? packet_ram_4__20_ : 
                    (N77)? packet_ram_5__20_ : 
                    (N79)? packet_ram_6__20_ : 
                    (N81)? packet_ram_7__20_ : 1'b0;
  assign T152[19] = (N74)? io_scr_req_bits_data[19] : 
                    (N76)? packet_ram_1__19_ : 
                    (N78)? packet_ram_2__19_ : 
                    (N80)? packet_ram_3__19_ : 
                    (N75)? packet_ram_4__19_ : 
                    (N77)? packet_ram_5__19_ : 
                    (N79)? packet_ram_6__19_ : 
                    (N81)? packet_ram_7__19_ : 1'b0;
  assign T152[18] = (N74)? io_scr_req_bits_data[18] : 
                    (N76)? packet_ram_1__18_ : 
                    (N78)? packet_ram_2__18_ : 
                    (N80)? packet_ram_3__18_ : 
                    (N75)? packet_ram_4__18_ : 
                    (N77)? packet_ram_5__18_ : 
                    (N79)? packet_ram_6__18_ : 
                    (N81)? packet_ram_7__18_ : 1'b0;
  assign T152[17] = (N74)? io_scr_req_bits_data[17] : 
                    (N76)? packet_ram_1__17_ : 
                    (N78)? packet_ram_2__17_ : 
                    (N80)? packet_ram_3__17_ : 
                    (N75)? packet_ram_4__17_ : 
                    (N77)? packet_ram_5__17_ : 
                    (N79)? packet_ram_6__17_ : 
                    (N81)? packet_ram_7__17_ : 1'b0;
  assign T152[16] = (N74)? io_scr_req_bits_data[16] : 
                    (N76)? packet_ram_1__16_ : 
                    (N78)? packet_ram_2__16_ : 
                    (N80)? packet_ram_3__16_ : 
                    (N75)? packet_ram_4__16_ : 
                    (N77)? packet_ram_5__16_ : 
                    (N79)? packet_ram_6__16_ : 
                    (N81)? packet_ram_7__16_ : 1'b0;
  assign T152[15] = (N74)? io_scr_req_bits_data[15] : 
                    (N76)? packet_ram_1__15_ : 
                    (N78)? packet_ram_2__15_ : 
                    (N80)? packet_ram_3__15_ : 
                    (N75)? packet_ram_4__15_ : 
                    (N77)? packet_ram_5__15_ : 
                    (N79)? packet_ram_6__15_ : 
                    (N81)? packet_ram_7__15_ : 1'b0;
  assign T152[14] = (N74)? io_scr_req_bits_data[14] : 
                    (N76)? packet_ram_1__14_ : 
                    (N78)? packet_ram_2__14_ : 
                    (N80)? packet_ram_3__14_ : 
                    (N75)? packet_ram_4__14_ : 
                    (N77)? packet_ram_5__14_ : 
                    (N79)? packet_ram_6__14_ : 
                    (N81)? packet_ram_7__14_ : 1'b0;
  assign T152[13] = (N74)? io_scr_req_bits_data[13] : 
                    (N76)? packet_ram_1__13_ : 
                    (N78)? packet_ram_2__13_ : 
                    (N80)? packet_ram_3__13_ : 
                    (N75)? packet_ram_4__13_ : 
                    (N77)? packet_ram_5__13_ : 
                    (N79)? packet_ram_6__13_ : 
                    (N81)? packet_ram_7__13_ : 1'b0;
  assign T152[12] = (N74)? io_scr_req_bits_data[12] : 
                    (N76)? packet_ram_1__12_ : 
                    (N78)? packet_ram_2__12_ : 
                    (N80)? packet_ram_3__12_ : 
                    (N75)? packet_ram_4__12_ : 
                    (N77)? packet_ram_5__12_ : 
                    (N79)? packet_ram_6__12_ : 
                    (N81)? packet_ram_7__12_ : 1'b0;
  assign T152[11] = (N74)? io_scr_req_bits_data[11] : 
                    (N76)? packet_ram_1__11_ : 
                    (N78)? packet_ram_2__11_ : 
                    (N80)? packet_ram_3__11_ : 
                    (N75)? packet_ram_4__11_ : 
                    (N77)? packet_ram_5__11_ : 
                    (N79)? packet_ram_6__11_ : 
                    (N81)? packet_ram_7__11_ : 1'b0;
  assign T152[10] = (N74)? io_scr_req_bits_data[10] : 
                    (N76)? packet_ram_1__10_ : 
                    (N78)? packet_ram_2__10_ : 
                    (N80)? packet_ram_3__10_ : 
                    (N75)? packet_ram_4__10_ : 
                    (N77)? packet_ram_5__10_ : 
                    (N79)? packet_ram_6__10_ : 
                    (N81)? packet_ram_7__10_ : 1'b0;
  assign T152[9] = (N74)? io_scr_req_bits_data[9] : 
                   (N76)? packet_ram_1__9_ : 
                   (N78)? packet_ram_2__9_ : 
                   (N80)? packet_ram_3__9_ : 
                   (N75)? packet_ram_4__9_ : 
                   (N77)? packet_ram_5__9_ : 
                   (N79)? packet_ram_6__9_ : 
                   (N81)? packet_ram_7__9_ : 1'b0;
  assign T152[8] = (N74)? io_scr_req_bits_data[8] : 
                   (N76)? packet_ram_1__8_ : 
                   (N78)? packet_ram_2__8_ : 
                   (N80)? packet_ram_3__8_ : 
                   (N75)? packet_ram_4__8_ : 
                   (N77)? packet_ram_5__8_ : 
                   (N79)? packet_ram_6__8_ : 
                   (N81)? packet_ram_7__8_ : 1'b0;
  assign T152[7] = (N74)? io_scr_req_bits_data[7] : 
                   (N76)? packet_ram_1__7_ : 
                   (N78)? packet_ram_2__7_ : 
                   (N80)? packet_ram_3__7_ : 
                   (N75)? packet_ram_4__7_ : 
                   (N77)? packet_ram_5__7_ : 
                   (N79)? packet_ram_6__7_ : 
                   (N81)? packet_ram_7__7_ : 1'b0;
  assign T152[6] = (N74)? io_scr_req_bits_data[6] : 
                   (N76)? packet_ram_1__6_ : 
                   (N78)? packet_ram_2__6_ : 
                   (N80)? packet_ram_3__6_ : 
                   (N75)? packet_ram_4__6_ : 
                   (N77)? packet_ram_5__6_ : 
                   (N79)? packet_ram_6__6_ : 
                   (N81)? packet_ram_7__6_ : 1'b0;
  assign T152[5] = (N74)? io_scr_req_bits_data[5] : 
                   (N76)? packet_ram_1__5_ : 
                   (N78)? packet_ram_2__5_ : 
                   (N80)? packet_ram_3__5_ : 
                   (N75)? packet_ram_4__5_ : 
                   (N77)? packet_ram_5__5_ : 
                   (N79)? packet_ram_6__5_ : 
                   (N81)? packet_ram_7__5_ : 1'b0;
  assign T152[4] = (N74)? io_scr_req_bits_data[4] : 
                   (N76)? packet_ram_1__4_ : 
                   (N78)? packet_ram_2__4_ : 
                   (N80)? packet_ram_3__4_ : 
                   (N75)? packet_ram_4__4_ : 
                   (N77)? packet_ram_5__4_ : 
                   (N79)? packet_ram_6__4_ : 
                   (N81)? packet_ram_7__4_ : 1'b0;
  assign T152[3] = (N74)? io_scr_req_bits_data[3] : 
                   (N76)? packet_ram_1__3_ : 
                   (N78)? packet_ram_2__3_ : 
                   (N80)? packet_ram_3__3_ : 
                   (N75)? packet_ram_4__3_ : 
                   (N77)? packet_ram_5__3_ : 
                   (N79)? packet_ram_6__3_ : 
                   (N81)? packet_ram_7__3_ : 1'b0;
  assign T152[2] = (N74)? io_scr_req_bits_data[2] : 
                   (N76)? packet_ram_1__2_ : 
                   (N78)? packet_ram_2__2_ : 
                   (N80)? packet_ram_3__2_ : 
                   (N75)? packet_ram_4__2_ : 
                   (N77)? packet_ram_5__2_ : 
                   (N79)? packet_ram_6__2_ : 
                   (N81)? packet_ram_7__2_ : 1'b0;
  assign T152[1] = (N74)? io_scr_req_bits_data[1] : 
                   (N76)? packet_ram_1__1_ : 
                   (N78)? packet_ram_2__1_ : 
                   (N80)? packet_ram_3__1_ : 
                   (N75)? packet_ram_4__1_ : 
                   (N77)? packet_ram_5__1_ : 
                   (N79)? packet_ram_6__1_ : 
                   (N81)? packet_ram_7__1_ : 1'b0;
  assign T152[0] = (N74)? io_scr_req_bits_data[0] : 
                   (N76)? packet_ram_1__0_ : 
                   (N78)? packet_ram_2__0_ : 
                   (N80)? packet_ram_3__0_ : 
                   (N75)? packet_ram_4__0_ : 
                   (N77)? packet_ram_5__0_ : 
                   (N79)? packet_ram_6__0_ : 
                   (N81)? packet_ram_7__0_ : 1'b0;
  assign T152[127] = (N87)? io_scr_req_bits_data[63] : 
                     (N89)? packet_ram_1__63_ : 
                     (N91)? packet_ram_2__63_ : 
                     (N93)? packet_ram_3__63_ : 
                     (N88)? packet_ram_4__63_ : 
                     (N90)? packet_ram_5__63_ : 
                     (N92)? packet_ram_6__63_ : 
                     (N94)? packet_ram_7__63_ : 1'b0;
  assign T152[126] = (N87)? io_scr_req_bits_data[62] : 
                     (N89)? packet_ram_1__62_ : 
                     (N91)? packet_ram_2__62_ : 
                     (N93)? packet_ram_3__62_ : 
                     (N88)? packet_ram_4__62_ : 
                     (N90)? packet_ram_5__62_ : 
                     (N92)? packet_ram_6__62_ : 
                     (N94)? packet_ram_7__62_ : 1'b0;
  assign T152[125] = (N87)? io_scr_req_bits_data[61] : 
                     (N89)? packet_ram_1__61_ : 
                     (N91)? packet_ram_2__61_ : 
                     (N93)? packet_ram_3__61_ : 
                     (N88)? packet_ram_4__61_ : 
                     (N90)? packet_ram_5__61_ : 
                     (N92)? packet_ram_6__61_ : 
                     (N94)? packet_ram_7__61_ : 1'b0;
  assign T152[124] = (N87)? io_scr_req_bits_data[60] : 
                     (N89)? packet_ram_1__60_ : 
                     (N91)? packet_ram_2__60_ : 
                     (N93)? packet_ram_3__60_ : 
                     (N88)? packet_ram_4__60_ : 
                     (N90)? packet_ram_5__60_ : 
                     (N92)? packet_ram_6__60_ : 
                     (N94)? packet_ram_7__60_ : 1'b0;
  assign T152[123] = (N87)? io_scr_req_bits_data[59] : 
                     (N89)? packet_ram_1__59_ : 
                     (N91)? packet_ram_2__59_ : 
                     (N93)? packet_ram_3__59_ : 
                     (N88)? packet_ram_4__59_ : 
                     (N90)? packet_ram_5__59_ : 
                     (N92)? packet_ram_6__59_ : 
                     (N94)? packet_ram_7__59_ : 1'b0;
  assign T152[122] = (N87)? io_scr_req_bits_data[58] : 
                     (N89)? packet_ram_1__58_ : 
                     (N91)? packet_ram_2__58_ : 
                     (N93)? packet_ram_3__58_ : 
                     (N88)? packet_ram_4__58_ : 
                     (N90)? packet_ram_5__58_ : 
                     (N92)? packet_ram_6__58_ : 
                     (N94)? packet_ram_7__58_ : 1'b0;
  assign T152[121] = (N87)? io_scr_req_bits_data[57] : 
                     (N89)? packet_ram_1__57_ : 
                     (N91)? packet_ram_2__57_ : 
                     (N93)? packet_ram_3__57_ : 
                     (N88)? packet_ram_4__57_ : 
                     (N90)? packet_ram_5__57_ : 
                     (N92)? packet_ram_6__57_ : 
                     (N94)? packet_ram_7__57_ : 1'b0;
  assign T152[120] = (N87)? io_scr_req_bits_data[56] : 
                     (N89)? packet_ram_1__56_ : 
                     (N91)? packet_ram_2__56_ : 
                     (N93)? packet_ram_3__56_ : 
                     (N88)? packet_ram_4__56_ : 
                     (N90)? packet_ram_5__56_ : 
                     (N92)? packet_ram_6__56_ : 
                     (N94)? packet_ram_7__56_ : 1'b0;
  assign T152[119] = (N87)? io_scr_req_bits_data[55] : 
                     (N89)? packet_ram_1__55_ : 
                     (N91)? packet_ram_2__55_ : 
                     (N93)? packet_ram_3__55_ : 
                     (N88)? packet_ram_4__55_ : 
                     (N90)? packet_ram_5__55_ : 
                     (N92)? packet_ram_6__55_ : 
                     (N94)? packet_ram_7__55_ : 1'b0;
  assign T152[118] = (N87)? io_scr_req_bits_data[54] : 
                     (N89)? packet_ram_1__54_ : 
                     (N91)? packet_ram_2__54_ : 
                     (N93)? packet_ram_3__54_ : 
                     (N88)? packet_ram_4__54_ : 
                     (N90)? packet_ram_5__54_ : 
                     (N92)? packet_ram_6__54_ : 
                     (N94)? packet_ram_7__54_ : 1'b0;
  assign T152[117] = (N87)? io_scr_req_bits_data[53] : 
                     (N89)? packet_ram_1__53_ : 
                     (N91)? packet_ram_2__53_ : 
                     (N93)? packet_ram_3__53_ : 
                     (N88)? packet_ram_4__53_ : 
                     (N90)? packet_ram_5__53_ : 
                     (N92)? packet_ram_6__53_ : 
                     (N94)? packet_ram_7__53_ : 1'b0;
  assign T152[116] = (N87)? io_scr_req_bits_data[52] : 
                     (N89)? packet_ram_1__52_ : 
                     (N91)? packet_ram_2__52_ : 
                     (N93)? packet_ram_3__52_ : 
                     (N88)? packet_ram_4__52_ : 
                     (N90)? packet_ram_5__52_ : 
                     (N92)? packet_ram_6__52_ : 
                     (N94)? packet_ram_7__52_ : 1'b0;
  assign T152[115] = (N87)? io_scr_req_bits_data[51] : 
                     (N89)? packet_ram_1__51_ : 
                     (N91)? packet_ram_2__51_ : 
                     (N93)? packet_ram_3__51_ : 
                     (N88)? packet_ram_4__51_ : 
                     (N90)? packet_ram_5__51_ : 
                     (N92)? packet_ram_6__51_ : 
                     (N94)? packet_ram_7__51_ : 1'b0;
  assign T152[114] = (N87)? io_scr_req_bits_data[50] : 
                     (N89)? packet_ram_1__50_ : 
                     (N91)? packet_ram_2__50_ : 
                     (N93)? packet_ram_3__50_ : 
                     (N88)? packet_ram_4__50_ : 
                     (N90)? packet_ram_5__50_ : 
                     (N92)? packet_ram_6__50_ : 
                     (N94)? packet_ram_7__50_ : 1'b0;
  assign T152[113] = (N87)? io_scr_req_bits_data[49] : 
                     (N89)? packet_ram_1__49_ : 
                     (N91)? packet_ram_2__49_ : 
                     (N93)? packet_ram_3__49_ : 
                     (N88)? packet_ram_4__49_ : 
                     (N90)? packet_ram_5__49_ : 
                     (N92)? packet_ram_6__49_ : 
                     (N94)? packet_ram_7__49_ : 1'b0;
  assign T152[112] = (N87)? io_scr_req_bits_data[48] : 
                     (N89)? packet_ram_1__48_ : 
                     (N91)? packet_ram_2__48_ : 
                     (N93)? packet_ram_3__48_ : 
                     (N88)? packet_ram_4__48_ : 
                     (N90)? packet_ram_5__48_ : 
                     (N92)? packet_ram_6__48_ : 
                     (N94)? packet_ram_7__48_ : 1'b0;
  assign T152[111] = (N87)? io_scr_req_bits_data[47] : 
                     (N89)? packet_ram_1__47_ : 
                     (N91)? packet_ram_2__47_ : 
                     (N93)? packet_ram_3__47_ : 
                     (N88)? packet_ram_4__47_ : 
                     (N90)? packet_ram_5__47_ : 
                     (N92)? packet_ram_6__47_ : 
                     (N94)? packet_ram_7__47_ : 1'b0;
  assign T152[110] = (N87)? io_scr_req_bits_data[46] : 
                     (N89)? packet_ram_1__46_ : 
                     (N91)? packet_ram_2__46_ : 
                     (N93)? packet_ram_3__46_ : 
                     (N88)? packet_ram_4__46_ : 
                     (N90)? packet_ram_5__46_ : 
                     (N92)? packet_ram_6__46_ : 
                     (N94)? packet_ram_7__46_ : 1'b0;
  assign T152[109] = (N87)? io_scr_req_bits_data[45] : 
                     (N89)? packet_ram_1__45_ : 
                     (N91)? packet_ram_2__45_ : 
                     (N93)? packet_ram_3__45_ : 
                     (N88)? packet_ram_4__45_ : 
                     (N90)? packet_ram_5__45_ : 
                     (N92)? packet_ram_6__45_ : 
                     (N94)? packet_ram_7__45_ : 1'b0;
  assign T152[108] = (N87)? io_scr_req_bits_data[44] : 
                     (N89)? packet_ram_1__44_ : 
                     (N91)? packet_ram_2__44_ : 
                     (N93)? packet_ram_3__44_ : 
                     (N88)? packet_ram_4__44_ : 
                     (N90)? packet_ram_5__44_ : 
                     (N92)? packet_ram_6__44_ : 
                     (N94)? packet_ram_7__44_ : 1'b0;
  assign T152[107] = (N87)? io_scr_req_bits_data[43] : 
                     (N89)? packet_ram_1__43_ : 
                     (N91)? packet_ram_2__43_ : 
                     (N93)? packet_ram_3__43_ : 
                     (N88)? packet_ram_4__43_ : 
                     (N90)? packet_ram_5__43_ : 
                     (N92)? packet_ram_6__43_ : 
                     (N94)? packet_ram_7__43_ : 1'b0;
  assign T152[106] = (N87)? io_scr_req_bits_data[42] : 
                     (N89)? packet_ram_1__42_ : 
                     (N91)? packet_ram_2__42_ : 
                     (N93)? packet_ram_3__42_ : 
                     (N88)? packet_ram_4__42_ : 
                     (N90)? packet_ram_5__42_ : 
                     (N92)? packet_ram_6__42_ : 
                     (N94)? packet_ram_7__42_ : 1'b0;
  assign T152[105] = (N87)? io_scr_req_bits_data[41] : 
                     (N89)? packet_ram_1__41_ : 
                     (N91)? packet_ram_2__41_ : 
                     (N93)? packet_ram_3__41_ : 
                     (N88)? packet_ram_4__41_ : 
                     (N90)? packet_ram_5__41_ : 
                     (N92)? packet_ram_6__41_ : 
                     (N94)? packet_ram_7__41_ : 1'b0;
  assign T152[104] = (N87)? io_scr_req_bits_data[40] : 
                     (N89)? packet_ram_1__40_ : 
                     (N91)? packet_ram_2__40_ : 
                     (N93)? packet_ram_3__40_ : 
                     (N88)? packet_ram_4__40_ : 
                     (N90)? packet_ram_5__40_ : 
                     (N92)? packet_ram_6__40_ : 
                     (N94)? packet_ram_7__40_ : 1'b0;
  assign T152[103] = (N87)? io_scr_req_bits_data[39] : 
                     (N89)? packet_ram_1__39_ : 
                     (N91)? packet_ram_2__39_ : 
                     (N93)? packet_ram_3__39_ : 
                     (N88)? packet_ram_4__39_ : 
                     (N90)? packet_ram_5__39_ : 
                     (N92)? packet_ram_6__39_ : 
                     (N94)? packet_ram_7__39_ : 1'b0;
  assign T152[102] = (N87)? io_scr_req_bits_data[38] : 
                     (N89)? packet_ram_1__38_ : 
                     (N91)? packet_ram_2__38_ : 
                     (N93)? packet_ram_3__38_ : 
                     (N88)? packet_ram_4__38_ : 
                     (N90)? packet_ram_5__38_ : 
                     (N92)? packet_ram_6__38_ : 
                     (N94)? packet_ram_7__38_ : 1'b0;
  assign T152[101] = (N87)? io_scr_req_bits_data[37] : 
                     (N89)? packet_ram_1__37_ : 
                     (N91)? packet_ram_2__37_ : 
                     (N93)? packet_ram_3__37_ : 
                     (N88)? packet_ram_4__37_ : 
                     (N90)? packet_ram_5__37_ : 
                     (N92)? packet_ram_6__37_ : 
                     (N94)? packet_ram_7__37_ : 1'b0;
  assign T152[100] = (N87)? io_scr_req_bits_data[36] : 
                     (N89)? packet_ram_1__36_ : 
                     (N91)? packet_ram_2__36_ : 
                     (N93)? packet_ram_3__36_ : 
                     (N88)? packet_ram_4__36_ : 
                     (N90)? packet_ram_5__36_ : 
                     (N92)? packet_ram_6__36_ : 
                     (N94)? packet_ram_7__36_ : 1'b0;
  assign T152[99] = (N87)? io_scr_req_bits_data[35] : 
                    (N89)? packet_ram_1__35_ : 
                    (N91)? packet_ram_2__35_ : 
                    (N93)? packet_ram_3__35_ : 
                    (N88)? packet_ram_4__35_ : 
                    (N90)? packet_ram_5__35_ : 
                    (N92)? packet_ram_6__35_ : 
                    (N94)? packet_ram_7__35_ : 1'b0;
  assign T152[98] = (N87)? io_scr_req_bits_data[34] : 
                    (N89)? packet_ram_1__34_ : 
                    (N91)? packet_ram_2__34_ : 
                    (N93)? packet_ram_3__34_ : 
                    (N88)? packet_ram_4__34_ : 
                    (N90)? packet_ram_5__34_ : 
                    (N92)? packet_ram_6__34_ : 
                    (N94)? packet_ram_7__34_ : 1'b0;
  assign T152[97] = (N87)? io_scr_req_bits_data[33] : 
                    (N89)? packet_ram_1__33_ : 
                    (N91)? packet_ram_2__33_ : 
                    (N93)? packet_ram_3__33_ : 
                    (N88)? packet_ram_4__33_ : 
                    (N90)? packet_ram_5__33_ : 
                    (N92)? packet_ram_6__33_ : 
                    (N94)? packet_ram_7__33_ : 1'b0;
  assign T152[96] = (N87)? io_scr_req_bits_data[32] : 
                    (N89)? packet_ram_1__32_ : 
                    (N91)? packet_ram_2__32_ : 
                    (N93)? packet_ram_3__32_ : 
                    (N88)? packet_ram_4__32_ : 
                    (N90)? packet_ram_5__32_ : 
                    (N92)? packet_ram_6__32_ : 
                    (N94)? packet_ram_7__32_ : 1'b0;
  assign T152[95] = (N87)? io_scr_req_bits_data[31] : 
                    (N89)? packet_ram_1__31_ : 
                    (N91)? packet_ram_2__31_ : 
                    (N93)? packet_ram_3__31_ : 
                    (N88)? packet_ram_4__31_ : 
                    (N90)? packet_ram_5__31_ : 
                    (N92)? packet_ram_6__31_ : 
                    (N94)? packet_ram_7__31_ : 1'b0;
  assign T152[94] = (N87)? io_scr_req_bits_data[30] : 
                    (N89)? packet_ram_1__30_ : 
                    (N91)? packet_ram_2__30_ : 
                    (N93)? packet_ram_3__30_ : 
                    (N88)? packet_ram_4__30_ : 
                    (N90)? packet_ram_5__30_ : 
                    (N92)? packet_ram_6__30_ : 
                    (N94)? packet_ram_7__30_ : 1'b0;
  assign T152[93] = (N87)? io_scr_req_bits_data[29] : 
                    (N89)? packet_ram_1__29_ : 
                    (N91)? packet_ram_2__29_ : 
                    (N93)? packet_ram_3__29_ : 
                    (N88)? packet_ram_4__29_ : 
                    (N90)? packet_ram_5__29_ : 
                    (N92)? packet_ram_6__29_ : 
                    (N94)? packet_ram_7__29_ : 1'b0;
  assign T152[92] = (N87)? io_scr_req_bits_data[28] : 
                    (N89)? packet_ram_1__28_ : 
                    (N91)? packet_ram_2__28_ : 
                    (N93)? packet_ram_3__28_ : 
                    (N88)? packet_ram_4__28_ : 
                    (N90)? packet_ram_5__28_ : 
                    (N92)? packet_ram_6__28_ : 
                    (N94)? packet_ram_7__28_ : 1'b0;
  assign T152[91] = (N87)? io_scr_req_bits_data[27] : 
                    (N89)? packet_ram_1__27_ : 
                    (N91)? packet_ram_2__27_ : 
                    (N93)? packet_ram_3__27_ : 
                    (N88)? packet_ram_4__27_ : 
                    (N90)? packet_ram_5__27_ : 
                    (N92)? packet_ram_6__27_ : 
                    (N94)? packet_ram_7__27_ : 1'b0;
  assign T152[90] = (N87)? io_scr_req_bits_data[26] : 
                    (N89)? packet_ram_1__26_ : 
                    (N91)? packet_ram_2__26_ : 
                    (N93)? packet_ram_3__26_ : 
                    (N88)? packet_ram_4__26_ : 
                    (N90)? packet_ram_5__26_ : 
                    (N92)? packet_ram_6__26_ : 
                    (N94)? packet_ram_7__26_ : 1'b0;
  assign T152[89] = (N87)? io_scr_req_bits_data[25] : 
                    (N89)? packet_ram_1__25_ : 
                    (N91)? packet_ram_2__25_ : 
                    (N93)? packet_ram_3__25_ : 
                    (N88)? packet_ram_4__25_ : 
                    (N90)? packet_ram_5__25_ : 
                    (N92)? packet_ram_6__25_ : 
                    (N94)? packet_ram_7__25_ : 1'b0;
  assign T152[88] = (N87)? io_scr_req_bits_data[24] : 
                    (N89)? packet_ram_1__24_ : 
                    (N91)? packet_ram_2__24_ : 
                    (N93)? packet_ram_3__24_ : 
                    (N88)? packet_ram_4__24_ : 
                    (N90)? packet_ram_5__24_ : 
                    (N92)? packet_ram_6__24_ : 
                    (N94)? packet_ram_7__24_ : 1'b0;
  assign T152[87] = (N87)? io_scr_req_bits_data[23] : 
                    (N89)? packet_ram_1__23_ : 
                    (N91)? packet_ram_2__23_ : 
                    (N93)? packet_ram_3__23_ : 
                    (N88)? packet_ram_4__23_ : 
                    (N90)? packet_ram_5__23_ : 
                    (N92)? packet_ram_6__23_ : 
                    (N94)? packet_ram_7__23_ : 1'b0;
  assign T152[86] = (N87)? io_scr_req_bits_data[22] : 
                    (N89)? packet_ram_1__22_ : 
                    (N91)? packet_ram_2__22_ : 
                    (N93)? packet_ram_3__22_ : 
                    (N88)? packet_ram_4__22_ : 
                    (N90)? packet_ram_5__22_ : 
                    (N92)? packet_ram_6__22_ : 
                    (N94)? packet_ram_7__22_ : 1'b0;
  assign T152[85] = (N87)? io_scr_req_bits_data[21] : 
                    (N89)? packet_ram_1__21_ : 
                    (N91)? packet_ram_2__21_ : 
                    (N93)? packet_ram_3__21_ : 
                    (N88)? packet_ram_4__21_ : 
                    (N90)? packet_ram_5__21_ : 
                    (N92)? packet_ram_6__21_ : 
                    (N94)? packet_ram_7__21_ : 1'b0;
  assign T152[84] = (N87)? io_scr_req_bits_data[20] : 
                    (N89)? packet_ram_1__20_ : 
                    (N91)? packet_ram_2__20_ : 
                    (N93)? packet_ram_3__20_ : 
                    (N88)? packet_ram_4__20_ : 
                    (N90)? packet_ram_5__20_ : 
                    (N92)? packet_ram_6__20_ : 
                    (N94)? packet_ram_7__20_ : 1'b0;
  assign T152[83] = (N87)? io_scr_req_bits_data[19] : 
                    (N89)? packet_ram_1__19_ : 
                    (N91)? packet_ram_2__19_ : 
                    (N93)? packet_ram_3__19_ : 
                    (N88)? packet_ram_4__19_ : 
                    (N90)? packet_ram_5__19_ : 
                    (N92)? packet_ram_6__19_ : 
                    (N94)? packet_ram_7__19_ : 1'b0;
  assign T152[82] = (N87)? io_scr_req_bits_data[18] : 
                    (N89)? packet_ram_1__18_ : 
                    (N91)? packet_ram_2__18_ : 
                    (N93)? packet_ram_3__18_ : 
                    (N88)? packet_ram_4__18_ : 
                    (N90)? packet_ram_5__18_ : 
                    (N92)? packet_ram_6__18_ : 
                    (N94)? packet_ram_7__18_ : 1'b0;
  assign T152[81] = (N87)? io_scr_req_bits_data[17] : 
                    (N89)? packet_ram_1__17_ : 
                    (N91)? packet_ram_2__17_ : 
                    (N93)? packet_ram_3__17_ : 
                    (N88)? packet_ram_4__17_ : 
                    (N90)? packet_ram_5__17_ : 
                    (N92)? packet_ram_6__17_ : 
                    (N94)? packet_ram_7__17_ : 1'b0;
  assign T152[80] = (N87)? io_scr_req_bits_data[16] : 
                    (N89)? packet_ram_1__16_ : 
                    (N91)? packet_ram_2__16_ : 
                    (N93)? packet_ram_3__16_ : 
                    (N88)? packet_ram_4__16_ : 
                    (N90)? packet_ram_5__16_ : 
                    (N92)? packet_ram_6__16_ : 
                    (N94)? packet_ram_7__16_ : 1'b0;
  assign T152[79] = (N87)? io_scr_req_bits_data[15] : 
                    (N89)? packet_ram_1__15_ : 
                    (N91)? packet_ram_2__15_ : 
                    (N93)? packet_ram_3__15_ : 
                    (N88)? packet_ram_4__15_ : 
                    (N90)? packet_ram_5__15_ : 
                    (N92)? packet_ram_6__15_ : 
                    (N94)? packet_ram_7__15_ : 1'b0;
  assign T152[78] = (N87)? io_scr_req_bits_data[14] : 
                    (N89)? packet_ram_1__14_ : 
                    (N91)? packet_ram_2__14_ : 
                    (N93)? packet_ram_3__14_ : 
                    (N88)? packet_ram_4__14_ : 
                    (N90)? packet_ram_5__14_ : 
                    (N92)? packet_ram_6__14_ : 
                    (N94)? packet_ram_7__14_ : 1'b0;
  assign T152[77] = (N87)? io_scr_req_bits_data[13] : 
                    (N89)? packet_ram_1__13_ : 
                    (N91)? packet_ram_2__13_ : 
                    (N93)? packet_ram_3__13_ : 
                    (N88)? packet_ram_4__13_ : 
                    (N90)? packet_ram_5__13_ : 
                    (N92)? packet_ram_6__13_ : 
                    (N94)? packet_ram_7__13_ : 1'b0;
  assign T152[76] = (N87)? io_scr_req_bits_data[12] : 
                    (N89)? packet_ram_1__12_ : 
                    (N91)? packet_ram_2__12_ : 
                    (N93)? packet_ram_3__12_ : 
                    (N88)? packet_ram_4__12_ : 
                    (N90)? packet_ram_5__12_ : 
                    (N92)? packet_ram_6__12_ : 
                    (N94)? packet_ram_7__12_ : 1'b0;
  assign T152[75] = (N87)? io_scr_req_bits_data[11] : 
                    (N89)? packet_ram_1__11_ : 
                    (N91)? packet_ram_2__11_ : 
                    (N93)? packet_ram_3__11_ : 
                    (N88)? packet_ram_4__11_ : 
                    (N90)? packet_ram_5__11_ : 
                    (N92)? packet_ram_6__11_ : 
                    (N94)? packet_ram_7__11_ : 1'b0;
  assign T152[74] = (N87)? io_scr_req_bits_data[10] : 
                    (N89)? packet_ram_1__10_ : 
                    (N91)? packet_ram_2__10_ : 
                    (N93)? packet_ram_3__10_ : 
                    (N88)? packet_ram_4__10_ : 
                    (N90)? packet_ram_5__10_ : 
                    (N92)? packet_ram_6__10_ : 
                    (N94)? packet_ram_7__10_ : 1'b0;
  assign T152[73] = (N87)? io_scr_req_bits_data[9] : 
                    (N89)? packet_ram_1__9_ : 
                    (N91)? packet_ram_2__9_ : 
                    (N93)? packet_ram_3__9_ : 
                    (N88)? packet_ram_4__9_ : 
                    (N90)? packet_ram_5__9_ : 
                    (N92)? packet_ram_6__9_ : 
                    (N94)? packet_ram_7__9_ : 1'b0;
  assign T152[72] = (N87)? io_scr_req_bits_data[8] : 
                    (N89)? packet_ram_1__8_ : 
                    (N91)? packet_ram_2__8_ : 
                    (N93)? packet_ram_3__8_ : 
                    (N88)? packet_ram_4__8_ : 
                    (N90)? packet_ram_5__8_ : 
                    (N92)? packet_ram_6__8_ : 
                    (N94)? packet_ram_7__8_ : 1'b0;
  assign T152[71] = (N87)? io_scr_req_bits_data[7] : 
                    (N89)? packet_ram_1__7_ : 
                    (N91)? packet_ram_2__7_ : 
                    (N93)? packet_ram_3__7_ : 
                    (N88)? packet_ram_4__7_ : 
                    (N90)? packet_ram_5__7_ : 
                    (N92)? packet_ram_6__7_ : 
                    (N94)? packet_ram_7__7_ : 1'b0;
  assign T152[70] = (N87)? io_scr_req_bits_data[6] : 
                    (N89)? packet_ram_1__6_ : 
                    (N91)? packet_ram_2__6_ : 
                    (N93)? packet_ram_3__6_ : 
                    (N88)? packet_ram_4__6_ : 
                    (N90)? packet_ram_5__6_ : 
                    (N92)? packet_ram_6__6_ : 
                    (N94)? packet_ram_7__6_ : 1'b0;
  assign T152[69] = (N87)? io_scr_req_bits_data[5] : 
                    (N89)? packet_ram_1__5_ : 
                    (N91)? packet_ram_2__5_ : 
                    (N93)? packet_ram_3__5_ : 
                    (N88)? packet_ram_4__5_ : 
                    (N90)? packet_ram_5__5_ : 
                    (N92)? packet_ram_6__5_ : 
                    (N94)? packet_ram_7__5_ : 1'b0;
  assign T152[68] = (N87)? io_scr_req_bits_data[4] : 
                    (N89)? packet_ram_1__4_ : 
                    (N91)? packet_ram_2__4_ : 
                    (N93)? packet_ram_3__4_ : 
                    (N88)? packet_ram_4__4_ : 
                    (N90)? packet_ram_5__4_ : 
                    (N92)? packet_ram_6__4_ : 
                    (N94)? packet_ram_7__4_ : 1'b0;
  assign T152[67] = (N87)? io_scr_req_bits_data[3] : 
                    (N89)? packet_ram_1__3_ : 
                    (N91)? packet_ram_2__3_ : 
                    (N93)? packet_ram_3__3_ : 
                    (N88)? packet_ram_4__3_ : 
                    (N90)? packet_ram_5__3_ : 
                    (N92)? packet_ram_6__3_ : 
                    (N94)? packet_ram_7__3_ : 1'b0;
  assign T152[66] = (N87)? io_scr_req_bits_data[2] : 
                    (N89)? packet_ram_1__2_ : 
                    (N91)? packet_ram_2__2_ : 
                    (N93)? packet_ram_3__2_ : 
                    (N88)? packet_ram_4__2_ : 
                    (N90)? packet_ram_5__2_ : 
                    (N92)? packet_ram_6__2_ : 
                    (N94)? packet_ram_7__2_ : 1'b0;
  assign T152[65] = (N87)? io_scr_req_bits_data[1] : 
                    (N89)? packet_ram_1__1_ : 
                    (N91)? packet_ram_2__1_ : 
                    (N93)? packet_ram_3__1_ : 
                    (N88)? packet_ram_4__1_ : 
                    (N90)? packet_ram_5__1_ : 
                    (N92)? packet_ram_6__1_ : 
                    (N94)? packet_ram_7__1_ : 1'b0;
  assign T152[64] = (N87)? io_scr_req_bits_data[0] : 
                    (N89)? packet_ram_1__0_ : 
                    (N91)? packet_ram_2__0_ : 
                    (N93)? packet_ram_3__0_ : 
                    (N88)? packet_ram_4__0_ : 
                    (N90)? packet_ram_5__0_ : 
                    (N92)? packet_ram_6__0_ : 
                    (N94)? packet_ram_7__0_ : 1'b0;
  assign { SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2, SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4, SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6, SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11, SV2V_UNCONNECTED_12, SV2V_UNCONNECTED_13, SV2V_UNCONNECTED_14, SV2V_UNCONNECTED_15, SV2V_UNCONNECTED_16, SV2V_UNCONNECTED_17, SV2V_UNCONNECTED_18, SV2V_UNCONNECTED_19, SV2V_UNCONNECTED_20, SV2V_UNCONNECTED_21, SV2V_UNCONNECTED_22, SV2V_UNCONNECTED_23, SV2V_UNCONNECTED_24, SV2V_UNCONNECTED_25, SV2V_UNCONNECTED_26, SV2V_UNCONNECTED_27, SV2V_UNCONNECTED_28, SV2V_UNCONNECTED_29, SV2V_UNCONNECTED_30, SV2V_UNCONNECTED_31, SV2V_UNCONNECTED_32, SV2V_UNCONNECTED_33, SV2V_UNCONNECTED_34, SV2V_UNCONNECTED_35, SV2V_UNCONNECTED_36, SV2V_UNCONNECTED_37, SV2V_UNCONNECTED_38, SV2V_UNCONNECTED_39, SV2V_UNCONNECTED_40, SV2V_UNCONNECTED_41, SV2V_UNCONNECTED_42, SV2V_UNCONNECTED_43, SV2V_UNCONNECTED_44, SV2V_UNCONNECTED_45, SV2V_UNCONNECTED_46, SV2V_UNCONNECTED_47, SV2V_UNCONNECTED_48, io_host_out_bits } = tx_data >> { tx_subword_count, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign T196[63] = (N103)? io_scr_req_bits_data[63] : 
                    (N105)? packet_ram_1__63_ : 
                    (N107)? packet_ram_2__63_ : 
                    (N109)? packet_ram_3__63_ : 
                    (N104)? packet_ram_4__63_ : 
                    (N106)? packet_ram_5__63_ : 
                    (N108)? packet_ram_6__63_ : 
                    (N110)? packet_ram_7__63_ : 1'b0;
  assign T196[62] = (N103)? io_scr_req_bits_data[62] : 
                    (N105)? packet_ram_1__62_ : 
                    (N107)? packet_ram_2__62_ : 
                    (N109)? packet_ram_3__62_ : 
                    (N104)? packet_ram_4__62_ : 
                    (N106)? packet_ram_5__62_ : 
                    (N108)? packet_ram_6__62_ : 
                    (N110)? packet_ram_7__62_ : 1'b0;
  assign T196[61] = (N103)? io_scr_req_bits_data[61] : 
                    (N105)? packet_ram_1__61_ : 
                    (N107)? packet_ram_2__61_ : 
                    (N109)? packet_ram_3__61_ : 
                    (N104)? packet_ram_4__61_ : 
                    (N106)? packet_ram_5__61_ : 
                    (N108)? packet_ram_6__61_ : 
                    (N110)? packet_ram_7__61_ : 1'b0;
  assign T196[60] = (N103)? io_scr_req_bits_data[60] : 
                    (N105)? packet_ram_1__60_ : 
                    (N107)? packet_ram_2__60_ : 
                    (N109)? packet_ram_3__60_ : 
                    (N104)? packet_ram_4__60_ : 
                    (N106)? packet_ram_5__60_ : 
                    (N108)? packet_ram_6__60_ : 
                    (N110)? packet_ram_7__60_ : 1'b0;
  assign T196[59] = (N103)? io_scr_req_bits_data[59] : 
                    (N105)? packet_ram_1__59_ : 
                    (N107)? packet_ram_2__59_ : 
                    (N109)? packet_ram_3__59_ : 
                    (N104)? packet_ram_4__59_ : 
                    (N106)? packet_ram_5__59_ : 
                    (N108)? packet_ram_6__59_ : 
                    (N110)? packet_ram_7__59_ : 1'b0;
  assign T196[58] = (N103)? io_scr_req_bits_data[58] : 
                    (N105)? packet_ram_1__58_ : 
                    (N107)? packet_ram_2__58_ : 
                    (N109)? packet_ram_3__58_ : 
                    (N104)? packet_ram_4__58_ : 
                    (N106)? packet_ram_5__58_ : 
                    (N108)? packet_ram_6__58_ : 
                    (N110)? packet_ram_7__58_ : 1'b0;
  assign T196[57] = (N103)? io_scr_req_bits_data[57] : 
                    (N105)? packet_ram_1__57_ : 
                    (N107)? packet_ram_2__57_ : 
                    (N109)? packet_ram_3__57_ : 
                    (N104)? packet_ram_4__57_ : 
                    (N106)? packet_ram_5__57_ : 
                    (N108)? packet_ram_6__57_ : 
                    (N110)? packet_ram_7__57_ : 1'b0;
  assign T196[56] = (N103)? io_scr_req_bits_data[56] : 
                    (N105)? packet_ram_1__56_ : 
                    (N107)? packet_ram_2__56_ : 
                    (N109)? packet_ram_3__56_ : 
                    (N104)? packet_ram_4__56_ : 
                    (N106)? packet_ram_5__56_ : 
                    (N108)? packet_ram_6__56_ : 
                    (N110)? packet_ram_7__56_ : 1'b0;
  assign T196[55] = (N103)? io_scr_req_bits_data[55] : 
                    (N105)? packet_ram_1__55_ : 
                    (N107)? packet_ram_2__55_ : 
                    (N109)? packet_ram_3__55_ : 
                    (N104)? packet_ram_4__55_ : 
                    (N106)? packet_ram_5__55_ : 
                    (N108)? packet_ram_6__55_ : 
                    (N110)? packet_ram_7__55_ : 1'b0;
  assign T196[54] = (N103)? io_scr_req_bits_data[54] : 
                    (N105)? packet_ram_1__54_ : 
                    (N107)? packet_ram_2__54_ : 
                    (N109)? packet_ram_3__54_ : 
                    (N104)? packet_ram_4__54_ : 
                    (N106)? packet_ram_5__54_ : 
                    (N108)? packet_ram_6__54_ : 
                    (N110)? packet_ram_7__54_ : 1'b0;
  assign T196[53] = (N103)? io_scr_req_bits_data[53] : 
                    (N105)? packet_ram_1__53_ : 
                    (N107)? packet_ram_2__53_ : 
                    (N109)? packet_ram_3__53_ : 
                    (N104)? packet_ram_4__53_ : 
                    (N106)? packet_ram_5__53_ : 
                    (N108)? packet_ram_6__53_ : 
                    (N110)? packet_ram_7__53_ : 1'b0;
  assign T196[52] = (N103)? io_scr_req_bits_data[52] : 
                    (N105)? packet_ram_1__52_ : 
                    (N107)? packet_ram_2__52_ : 
                    (N109)? packet_ram_3__52_ : 
                    (N104)? packet_ram_4__52_ : 
                    (N106)? packet_ram_5__52_ : 
                    (N108)? packet_ram_6__52_ : 
                    (N110)? packet_ram_7__52_ : 1'b0;
  assign T196[51] = (N103)? io_scr_req_bits_data[51] : 
                    (N105)? packet_ram_1__51_ : 
                    (N107)? packet_ram_2__51_ : 
                    (N109)? packet_ram_3__51_ : 
                    (N104)? packet_ram_4__51_ : 
                    (N106)? packet_ram_5__51_ : 
                    (N108)? packet_ram_6__51_ : 
                    (N110)? packet_ram_7__51_ : 1'b0;
  assign T196[50] = (N103)? io_scr_req_bits_data[50] : 
                    (N105)? packet_ram_1__50_ : 
                    (N107)? packet_ram_2__50_ : 
                    (N109)? packet_ram_3__50_ : 
                    (N104)? packet_ram_4__50_ : 
                    (N106)? packet_ram_5__50_ : 
                    (N108)? packet_ram_6__50_ : 
                    (N110)? packet_ram_7__50_ : 1'b0;
  assign T196[49] = (N103)? io_scr_req_bits_data[49] : 
                    (N105)? packet_ram_1__49_ : 
                    (N107)? packet_ram_2__49_ : 
                    (N109)? packet_ram_3__49_ : 
                    (N104)? packet_ram_4__49_ : 
                    (N106)? packet_ram_5__49_ : 
                    (N108)? packet_ram_6__49_ : 
                    (N110)? packet_ram_7__49_ : 1'b0;
  assign T196[48] = (N103)? io_scr_req_bits_data[48] : 
                    (N105)? packet_ram_1__48_ : 
                    (N107)? packet_ram_2__48_ : 
                    (N109)? packet_ram_3__48_ : 
                    (N104)? packet_ram_4__48_ : 
                    (N106)? packet_ram_5__48_ : 
                    (N108)? packet_ram_6__48_ : 
                    (N110)? packet_ram_7__48_ : 1'b0;
  assign T196[47] = (N103)? io_scr_req_bits_data[47] : 
                    (N105)? packet_ram_1__47_ : 
                    (N107)? packet_ram_2__47_ : 
                    (N109)? packet_ram_3__47_ : 
                    (N104)? packet_ram_4__47_ : 
                    (N106)? packet_ram_5__47_ : 
                    (N108)? packet_ram_6__47_ : 
                    (N110)? packet_ram_7__47_ : 1'b0;
  assign T196[46] = (N103)? io_scr_req_bits_data[46] : 
                    (N105)? packet_ram_1__46_ : 
                    (N107)? packet_ram_2__46_ : 
                    (N109)? packet_ram_3__46_ : 
                    (N104)? packet_ram_4__46_ : 
                    (N106)? packet_ram_5__46_ : 
                    (N108)? packet_ram_6__46_ : 
                    (N110)? packet_ram_7__46_ : 1'b0;
  assign T196[45] = (N103)? io_scr_req_bits_data[45] : 
                    (N105)? packet_ram_1__45_ : 
                    (N107)? packet_ram_2__45_ : 
                    (N109)? packet_ram_3__45_ : 
                    (N104)? packet_ram_4__45_ : 
                    (N106)? packet_ram_5__45_ : 
                    (N108)? packet_ram_6__45_ : 
                    (N110)? packet_ram_7__45_ : 1'b0;
  assign T196[44] = (N103)? io_scr_req_bits_data[44] : 
                    (N105)? packet_ram_1__44_ : 
                    (N107)? packet_ram_2__44_ : 
                    (N109)? packet_ram_3__44_ : 
                    (N104)? packet_ram_4__44_ : 
                    (N106)? packet_ram_5__44_ : 
                    (N108)? packet_ram_6__44_ : 
                    (N110)? packet_ram_7__44_ : 1'b0;
  assign T196[43] = (N103)? io_scr_req_bits_data[43] : 
                    (N105)? packet_ram_1__43_ : 
                    (N107)? packet_ram_2__43_ : 
                    (N109)? packet_ram_3__43_ : 
                    (N104)? packet_ram_4__43_ : 
                    (N106)? packet_ram_5__43_ : 
                    (N108)? packet_ram_6__43_ : 
                    (N110)? packet_ram_7__43_ : 1'b0;
  assign T196[42] = (N103)? io_scr_req_bits_data[42] : 
                    (N105)? packet_ram_1__42_ : 
                    (N107)? packet_ram_2__42_ : 
                    (N109)? packet_ram_3__42_ : 
                    (N104)? packet_ram_4__42_ : 
                    (N106)? packet_ram_5__42_ : 
                    (N108)? packet_ram_6__42_ : 
                    (N110)? packet_ram_7__42_ : 1'b0;
  assign T196[41] = (N103)? io_scr_req_bits_data[41] : 
                    (N105)? packet_ram_1__41_ : 
                    (N107)? packet_ram_2__41_ : 
                    (N109)? packet_ram_3__41_ : 
                    (N104)? packet_ram_4__41_ : 
                    (N106)? packet_ram_5__41_ : 
                    (N108)? packet_ram_6__41_ : 
                    (N110)? packet_ram_7__41_ : 1'b0;
  assign T196[40] = (N103)? io_scr_req_bits_data[40] : 
                    (N105)? packet_ram_1__40_ : 
                    (N107)? packet_ram_2__40_ : 
                    (N109)? packet_ram_3__40_ : 
                    (N104)? packet_ram_4__40_ : 
                    (N106)? packet_ram_5__40_ : 
                    (N108)? packet_ram_6__40_ : 
                    (N110)? packet_ram_7__40_ : 1'b0;
  assign T196[39] = (N103)? io_scr_req_bits_data[39] : 
                    (N105)? packet_ram_1__39_ : 
                    (N107)? packet_ram_2__39_ : 
                    (N109)? packet_ram_3__39_ : 
                    (N104)? packet_ram_4__39_ : 
                    (N106)? packet_ram_5__39_ : 
                    (N108)? packet_ram_6__39_ : 
                    (N110)? packet_ram_7__39_ : 1'b0;
  assign T196[38] = (N103)? io_scr_req_bits_data[38] : 
                    (N105)? packet_ram_1__38_ : 
                    (N107)? packet_ram_2__38_ : 
                    (N109)? packet_ram_3__38_ : 
                    (N104)? packet_ram_4__38_ : 
                    (N106)? packet_ram_5__38_ : 
                    (N108)? packet_ram_6__38_ : 
                    (N110)? packet_ram_7__38_ : 1'b0;
  assign T196[37] = (N103)? io_scr_req_bits_data[37] : 
                    (N105)? packet_ram_1__37_ : 
                    (N107)? packet_ram_2__37_ : 
                    (N109)? packet_ram_3__37_ : 
                    (N104)? packet_ram_4__37_ : 
                    (N106)? packet_ram_5__37_ : 
                    (N108)? packet_ram_6__37_ : 
                    (N110)? packet_ram_7__37_ : 1'b0;
  assign T196[36] = (N103)? io_scr_req_bits_data[36] : 
                    (N105)? packet_ram_1__36_ : 
                    (N107)? packet_ram_2__36_ : 
                    (N109)? packet_ram_3__36_ : 
                    (N104)? packet_ram_4__36_ : 
                    (N106)? packet_ram_5__36_ : 
                    (N108)? packet_ram_6__36_ : 
                    (N110)? packet_ram_7__36_ : 1'b0;
  assign T196[35] = (N103)? io_scr_req_bits_data[35] : 
                    (N105)? packet_ram_1__35_ : 
                    (N107)? packet_ram_2__35_ : 
                    (N109)? packet_ram_3__35_ : 
                    (N104)? packet_ram_4__35_ : 
                    (N106)? packet_ram_5__35_ : 
                    (N108)? packet_ram_6__35_ : 
                    (N110)? packet_ram_7__35_ : 1'b0;
  assign T196[34] = (N103)? io_scr_req_bits_data[34] : 
                    (N105)? packet_ram_1__34_ : 
                    (N107)? packet_ram_2__34_ : 
                    (N109)? packet_ram_3__34_ : 
                    (N104)? packet_ram_4__34_ : 
                    (N106)? packet_ram_5__34_ : 
                    (N108)? packet_ram_6__34_ : 
                    (N110)? packet_ram_7__34_ : 1'b0;
  assign T196[33] = (N103)? io_scr_req_bits_data[33] : 
                    (N105)? packet_ram_1__33_ : 
                    (N107)? packet_ram_2__33_ : 
                    (N109)? packet_ram_3__33_ : 
                    (N104)? packet_ram_4__33_ : 
                    (N106)? packet_ram_5__33_ : 
                    (N108)? packet_ram_6__33_ : 
                    (N110)? packet_ram_7__33_ : 1'b0;
  assign T196[32] = (N103)? io_scr_req_bits_data[32] : 
                    (N105)? packet_ram_1__32_ : 
                    (N107)? packet_ram_2__32_ : 
                    (N109)? packet_ram_3__32_ : 
                    (N104)? packet_ram_4__32_ : 
                    (N106)? packet_ram_5__32_ : 
                    (N108)? packet_ram_6__32_ : 
                    (N110)? packet_ram_7__32_ : 1'b0;
  assign T196[31] = (N103)? io_scr_req_bits_data[31] : 
                    (N105)? packet_ram_1__31_ : 
                    (N107)? packet_ram_2__31_ : 
                    (N109)? packet_ram_3__31_ : 
                    (N104)? packet_ram_4__31_ : 
                    (N106)? packet_ram_5__31_ : 
                    (N108)? packet_ram_6__31_ : 
                    (N110)? packet_ram_7__31_ : 1'b0;
  assign T196[30] = (N103)? io_scr_req_bits_data[30] : 
                    (N105)? packet_ram_1__30_ : 
                    (N107)? packet_ram_2__30_ : 
                    (N109)? packet_ram_3__30_ : 
                    (N104)? packet_ram_4__30_ : 
                    (N106)? packet_ram_5__30_ : 
                    (N108)? packet_ram_6__30_ : 
                    (N110)? packet_ram_7__30_ : 1'b0;
  assign T196[29] = (N103)? io_scr_req_bits_data[29] : 
                    (N105)? packet_ram_1__29_ : 
                    (N107)? packet_ram_2__29_ : 
                    (N109)? packet_ram_3__29_ : 
                    (N104)? packet_ram_4__29_ : 
                    (N106)? packet_ram_5__29_ : 
                    (N108)? packet_ram_6__29_ : 
                    (N110)? packet_ram_7__29_ : 1'b0;
  assign T196[28] = (N103)? io_scr_req_bits_data[28] : 
                    (N105)? packet_ram_1__28_ : 
                    (N107)? packet_ram_2__28_ : 
                    (N109)? packet_ram_3__28_ : 
                    (N104)? packet_ram_4__28_ : 
                    (N106)? packet_ram_5__28_ : 
                    (N108)? packet_ram_6__28_ : 
                    (N110)? packet_ram_7__28_ : 1'b0;
  assign T196[27] = (N103)? io_scr_req_bits_data[27] : 
                    (N105)? packet_ram_1__27_ : 
                    (N107)? packet_ram_2__27_ : 
                    (N109)? packet_ram_3__27_ : 
                    (N104)? packet_ram_4__27_ : 
                    (N106)? packet_ram_5__27_ : 
                    (N108)? packet_ram_6__27_ : 
                    (N110)? packet_ram_7__27_ : 1'b0;
  assign T196[26] = (N103)? io_scr_req_bits_data[26] : 
                    (N105)? packet_ram_1__26_ : 
                    (N107)? packet_ram_2__26_ : 
                    (N109)? packet_ram_3__26_ : 
                    (N104)? packet_ram_4__26_ : 
                    (N106)? packet_ram_5__26_ : 
                    (N108)? packet_ram_6__26_ : 
                    (N110)? packet_ram_7__26_ : 1'b0;
  assign T196[25] = (N103)? io_scr_req_bits_data[25] : 
                    (N105)? packet_ram_1__25_ : 
                    (N107)? packet_ram_2__25_ : 
                    (N109)? packet_ram_3__25_ : 
                    (N104)? packet_ram_4__25_ : 
                    (N106)? packet_ram_5__25_ : 
                    (N108)? packet_ram_6__25_ : 
                    (N110)? packet_ram_7__25_ : 1'b0;
  assign T196[24] = (N103)? io_scr_req_bits_data[24] : 
                    (N105)? packet_ram_1__24_ : 
                    (N107)? packet_ram_2__24_ : 
                    (N109)? packet_ram_3__24_ : 
                    (N104)? packet_ram_4__24_ : 
                    (N106)? packet_ram_5__24_ : 
                    (N108)? packet_ram_6__24_ : 
                    (N110)? packet_ram_7__24_ : 1'b0;
  assign T196[23] = (N103)? io_scr_req_bits_data[23] : 
                    (N105)? packet_ram_1__23_ : 
                    (N107)? packet_ram_2__23_ : 
                    (N109)? packet_ram_3__23_ : 
                    (N104)? packet_ram_4__23_ : 
                    (N106)? packet_ram_5__23_ : 
                    (N108)? packet_ram_6__23_ : 
                    (N110)? packet_ram_7__23_ : 1'b0;
  assign T196[22] = (N103)? io_scr_req_bits_data[22] : 
                    (N105)? packet_ram_1__22_ : 
                    (N107)? packet_ram_2__22_ : 
                    (N109)? packet_ram_3__22_ : 
                    (N104)? packet_ram_4__22_ : 
                    (N106)? packet_ram_5__22_ : 
                    (N108)? packet_ram_6__22_ : 
                    (N110)? packet_ram_7__22_ : 1'b0;
  assign T196[21] = (N103)? io_scr_req_bits_data[21] : 
                    (N105)? packet_ram_1__21_ : 
                    (N107)? packet_ram_2__21_ : 
                    (N109)? packet_ram_3__21_ : 
                    (N104)? packet_ram_4__21_ : 
                    (N106)? packet_ram_5__21_ : 
                    (N108)? packet_ram_6__21_ : 
                    (N110)? packet_ram_7__21_ : 1'b0;
  assign T196[20] = (N103)? io_scr_req_bits_data[20] : 
                    (N105)? packet_ram_1__20_ : 
                    (N107)? packet_ram_2__20_ : 
                    (N109)? packet_ram_3__20_ : 
                    (N104)? packet_ram_4__20_ : 
                    (N106)? packet_ram_5__20_ : 
                    (N108)? packet_ram_6__20_ : 
                    (N110)? packet_ram_7__20_ : 1'b0;
  assign T196[19] = (N103)? io_scr_req_bits_data[19] : 
                    (N105)? packet_ram_1__19_ : 
                    (N107)? packet_ram_2__19_ : 
                    (N109)? packet_ram_3__19_ : 
                    (N104)? packet_ram_4__19_ : 
                    (N106)? packet_ram_5__19_ : 
                    (N108)? packet_ram_6__19_ : 
                    (N110)? packet_ram_7__19_ : 1'b0;
  assign T196[18] = (N103)? io_scr_req_bits_data[18] : 
                    (N105)? packet_ram_1__18_ : 
                    (N107)? packet_ram_2__18_ : 
                    (N109)? packet_ram_3__18_ : 
                    (N104)? packet_ram_4__18_ : 
                    (N106)? packet_ram_5__18_ : 
                    (N108)? packet_ram_6__18_ : 
                    (N110)? packet_ram_7__18_ : 1'b0;
  assign T196[17] = (N103)? io_scr_req_bits_data[17] : 
                    (N105)? packet_ram_1__17_ : 
                    (N107)? packet_ram_2__17_ : 
                    (N109)? packet_ram_3__17_ : 
                    (N104)? packet_ram_4__17_ : 
                    (N106)? packet_ram_5__17_ : 
                    (N108)? packet_ram_6__17_ : 
                    (N110)? packet_ram_7__17_ : 1'b0;
  assign T196[16] = (N103)? io_scr_req_bits_data[16] : 
                    (N105)? packet_ram_1__16_ : 
                    (N107)? packet_ram_2__16_ : 
                    (N109)? packet_ram_3__16_ : 
                    (N104)? packet_ram_4__16_ : 
                    (N106)? packet_ram_5__16_ : 
                    (N108)? packet_ram_6__16_ : 
                    (N110)? packet_ram_7__16_ : 1'b0;
  assign T196[15] = (N103)? io_scr_req_bits_data[15] : 
                    (N105)? packet_ram_1__15_ : 
                    (N107)? packet_ram_2__15_ : 
                    (N109)? packet_ram_3__15_ : 
                    (N104)? packet_ram_4__15_ : 
                    (N106)? packet_ram_5__15_ : 
                    (N108)? packet_ram_6__15_ : 
                    (N110)? packet_ram_7__15_ : 1'b0;
  assign T196[14] = (N103)? io_scr_req_bits_data[14] : 
                    (N105)? packet_ram_1__14_ : 
                    (N107)? packet_ram_2__14_ : 
                    (N109)? packet_ram_3__14_ : 
                    (N104)? packet_ram_4__14_ : 
                    (N106)? packet_ram_5__14_ : 
                    (N108)? packet_ram_6__14_ : 
                    (N110)? packet_ram_7__14_ : 1'b0;
  assign T196[13] = (N103)? io_scr_req_bits_data[13] : 
                    (N105)? packet_ram_1__13_ : 
                    (N107)? packet_ram_2__13_ : 
                    (N109)? packet_ram_3__13_ : 
                    (N104)? packet_ram_4__13_ : 
                    (N106)? packet_ram_5__13_ : 
                    (N108)? packet_ram_6__13_ : 
                    (N110)? packet_ram_7__13_ : 1'b0;
  assign T196[12] = (N103)? io_scr_req_bits_data[12] : 
                    (N105)? packet_ram_1__12_ : 
                    (N107)? packet_ram_2__12_ : 
                    (N109)? packet_ram_3__12_ : 
                    (N104)? packet_ram_4__12_ : 
                    (N106)? packet_ram_5__12_ : 
                    (N108)? packet_ram_6__12_ : 
                    (N110)? packet_ram_7__12_ : 1'b0;
  assign T196[11] = (N103)? io_scr_req_bits_data[11] : 
                    (N105)? packet_ram_1__11_ : 
                    (N107)? packet_ram_2__11_ : 
                    (N109)? packet_ram_3__11_ : 
                    (N104)? packet_ram_4__11_ : 
                    (N106)? packet_ram_5__11_ : 
                    (N108)? packet_ram_6__11_ : 
                    (N110)? packet_ram_7__11_ : 1'b0;
  assign T196[10] = (N103)? io_scr_req_bits_data[10] : 
                    (N105)? packet_ram_1__10_ : 
                    (N107)? packet_ram_2__10_ : 
                    (N109)? packet_ram_3__10_ : 
                    (N104)? packet_ram_4__10_ : 
                    (N106)? packet_ram_5__10_ : 
                    (N108)? packet_ram_6__10_ : 
                    (N110)? packet_ram_7__10_ : 1'b0;
  assign T196[9] = (N103)? io_scr_req_bits_data[9] : 
                   (N105)? packet_ram_1__9_ : 
                   (N107)? packet_ram_2__9_ : 
                   (N109)? packet_ram_3__9_ : 
                   (N104)? packet_ram_4__9_ : 
                   (N106)? packet_ram_5__9_ : 
                   (N108)? packet_ram_6__9_ : 
                   (N110)? packet_ram_7__9_ : 1'b0;
  assign T196[8] = (N103)? io_scr_req_bits_data[8] : 
                   (N105)? packet_ram_1__8_ : 
                   (N107)? packet_ram_2__8_ : 
                   (N109)? packet_ram_3__8_ : 
                   (N104)? packet_ram_4__8_ : 
                   (N106)? packet_ram_5__8_ : 
                   (N108)? packet_ram_6__8_ : 
                   (N110)? packet_ram_7__8_ : 1'b0;
  assign T196[7] = (N103)? io_scr_req_bits_data[7] : 
                   (N105)? packet_ram_1__7_ : 
                   (N107)? packet_ram_2__7_ : 
                   (N109)? packet_ram_3__7_ : 
                   (N104)? packet_ram_4__7_ : 
                   (N106)? packet_ram_5__7_ : 
                   (N108)? packet_ram_6__7_ : 
                   (N110)? packet_ram_7__7_ : 1'b0;
  assign T196[6] = (N103)? io_scr_req_bits_data[6] : 
                   (N105)? packet_ram_1__6_ : 
                   (N107)? packet_ram_2__6_ : 
                   (N109)? packet_ram_3__6_ : 
                   (N104)? packet_ram_4__6_ : 
                   (N106)? packet_ram_5__6_ : 
                   (N108)? packet_ram_6__6_ : 
                   (N110)? packet_ram_7__6_ : 1'b0;
  assign T196[5] = (N103)? io_scr_req_bits_data[5] : 
                   (N105)? packet_ram_1__5_ : 
                   (N107)? packet_ram_2__5_ : 
                   (N109)? packet_ram_3__5_ : 
                   (N104)? packet_ram_4__5_ : 
                   (N106)? packet_ram_5__5_ : 
                   (N108)? packet_ram_6__5_ : 
                   (N110)? packet_ram_7__5_ : 1'b0;
  assign T196[4] = (N103)? io_scr_req_bits_data[4] : 
                   (N105)? packet_ram_1__4_ : 
                   (N107)? packet_ram_2__4_ : 
                   (N109)? packet_ram_3__4_ : 
                   (N104)? packet_ram_4__4_ : 
                   (N106)? packet_ram_5__4_ : 
                   (N108)? packet_ram_6__4_ : 
                   (N110)? packet_ram_7__4_ : 1'b0;
  assign T196[3] = (N103)? io_scr_req_bits_data[3] : 
                   (N105)? packet_ram_1__3_ : 
                   (N107)? packet_ram_2__3_ : 
                   (N109)? packet_ram_3__3_ : 
                   (N104)? packet_ram_4__3_ : 
                   (N106)? packet_ram_5__3_ : 
                   (N108)? packet_ram_6__3_ : 
                   (N110)? packet_ram_7__3_ : 1'b0;
  assign T196[2] = (N103)? io_scr_req_bits_data[2] : 
                   (N105)? packet_ram_1__2_ : 
                   (N107)? packet_ram_2__2_ : 
                   (N109)? packet_ram_3__2_ : 
                   (N104)? packet_ram_4__2_ : 
                   (N106)? packet_ram_5__2_ : 
                   (N108)? packet_ram_6__2_ : 
                   (N110)? packet_ram_7__2_ : 1'b0;
  assign T196[1] = (N103)? io_scr_req_bits_data[1] : 
                   (N105)? packet_ram_1__1_ : 
                   (N107)? packet_ram_2__1_ : 
                   (N109)? packet_ram_3__1_ : 
                   (N104)? packet_ram_4__1_ : 
                   (N106)? packet_ram_5__1_ : 
                   (N108)? packet_ram_6__1_ : 
                   (N110)? packet_ram_7__1_ : 1'b0;
  assign T196[0] = (N103)? io_scr_req_bits_data[0] : 
                   (N105)? packet_ram_1__0_ : 
                   (N107)? packet_ram_2__0_ : 
                   (N109)? packet_ram_3__0_ : 
                   (N104)? packet_ram_4__0_ : 
                   (N106)? packet_ram_5__0_ : 
                   (N108)? packet_ram_6__0_ : 
                   (N110)? packet_ram_7__0_ : 1'b0;

  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__63_ <= N2381;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__62_ <= N2380;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__61_ <= N2379;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__60_ <= N2378;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__59_ <= N2377;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__58_ <= N2376;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__57_ <= N2375;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__56_ <= N2374;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__55_ <= N2373;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__54_ <= N2372;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__53_ <= N2371;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__52_ <= N2370;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__51_ <= N2369;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__50_ <= N2368;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__49_ <= N2367;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__48_ <= N2366;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__47_ <= N2365;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__46_ <= N2364;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__45_ <= N2363;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__44_ <= N2362;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__43_ <= N2361;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__42_ <= N2360;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__41_ <= N2359;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__40_ <= N2358;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__39_ <= N2357;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__38_ <= N2356;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__37_ <= N2355;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__36_ <= N2354;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__35_ <= N2353;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__34_ <= N2352;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__33_ <= N2351;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__32_ <= N2350;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__31_ <= N2349;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__30_ <= N2348;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__29_ <= N2347;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__28_ <= N2346;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__27_ <= N2345;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__26_ <= N2344;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__25_ <= N2343;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__24_ <= N2342;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__23_ <= N2341;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__22_ <= N2340;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__21_ <= N2339;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__20_ <= N2338;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__19_ <= N2337;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__18_ <= N2336;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__17_ <= N2335;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__16_ <= N2334;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__15_ <= N2333;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__14_ <= N2332;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__13_ <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__12_ <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__11_ <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__10_ <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__9_ <= N2327;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__8_ <= N2326;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__7_ <= N2325;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__6_ <= N2324;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__5_ <= N2323;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__4_ <= N2322;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__3_ <= N2321;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__2_ <= N2320;
    end 
  end


  always @(posedge clk) begin
    if(N2318) begin
      packet_ram_7__1_ <= N2319;
    end 
  end


  always @(posedge clk) begin
    if(N2316) begin
      packet_ram_7__0_ <= N2317;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__63_ <= N2315;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__62_ <= N2314;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__61_ <= N2313;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__60_ <= N2312;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__59_ <= N2311;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__58_ <= N2310;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__57_ <= N2309;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__56_ <= N2308;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__55_ <= N2307;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__54_ <= N2306;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__53_ <= N2305;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__52_ <= N2304;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__51_ <= N2303;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__50_ <= N2302;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__49_ <= N2301;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__48_ <= N2300;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__47_ <= N2299;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__46_ <= N2298;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__45_ <= N2297;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__44_ <= N2296;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__43_ <= N2295;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__42_ <= N2294;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__41_ <= N2293;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__40_ <= N2292;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__39_ <= N2291;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__38_ <= N2290;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__37_ <= N2289;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__36_ <= N2288;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__35_ <= N2287;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__34_ <= N2286;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__33_ <= N2285;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__32_ <= N2284;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__31_ <= N2283;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__30_ <= N2282;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__29_ <= N2281;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__28_ <= N2280;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__27_ <= N2279;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__26_ <= N2278;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__25_ <= N2277;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__24_ <= N2276;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__23_ <= N2275;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__22_ <= N2274;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__21_ <= N2273;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__20_ <= N2272;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__19_ <= N2271;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__18_ <= N2270;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__17_ <= N2269;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__16_ <= N2268;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      packet_ram_6__15_ <= N2267;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__14_ <= N2265;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__13_ <= N2264;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__12_ <= N2263;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__11_ <= N2262;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__10_ <= N2261;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__9_ <= N2260;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__8_ <= N2259;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__7_ <= N2258;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__6_ <= N2257;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__5_ <= N2256;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__4_ <= N2255;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__3_ <= N2254;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__2_ <= N2253;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__1_ <= N2252;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      packet_ram_6__0_ <= N2251;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__63_ <= N2249;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__62_ <= N2248;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__61_ <= N2247;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__60_ <= N2246;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__59_ <= N2245;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__58_ <= N2244;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__57_ <= N2243;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__56_ <= N2242;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__55_ <= N2241;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__54_ <= N2240;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__53_ <= N2239;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__52_ <= N2238;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__51_ <= N2237;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__50_ <= N2236;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__49_ <= N2235;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__48_ <= N2234;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__47_ <= N2233;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__46_ <= N2232;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__45_ <= N2231;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__44_ <= N2230;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__43_ <= N2229;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__42_ <= N2228;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__41_ <= N2227;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__40_ <= N2226;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__39_ <= N2225;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__38_ <= N2224;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__37_ <= N2223;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__36_ <= N2222;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__35_ <= N2221;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__34_ <= N2220;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__33_ <= N2219;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__32_ <= N2218;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__31_ <= N2217;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__30_ <= N2216;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__29_ <= N2215;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__28_ <= N2214;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__27_ <= N2213;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__26_ <= N2212;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__25_ <= N2211;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__24_ <= N2210;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__23_ <= N2209;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__22_ <= N2208;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__21_ <= N2207;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__20_ <= N2206;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__19_ <= N2205;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__18_ <= N2204;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__17_ <= N2203;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__16_ <= N2202;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__15_ <= N2201;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__14_ <= N2200;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__13_ <= N2199;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__12_ <= N2198;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__11_ <= N2197;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__10_ <= N2196;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__9_ <= N2195;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__8_ <= N2194;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__7_ <= N2193;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__6_ <= N2192;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__5_ <= N2191;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__4_ <= N2190;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__3_ <= N2189;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__2_ <= N2188;
    end 
  end


  always @(posedge clk) begin
    if(N2186) begin
      packet_ram_5__1_ <= N2187;
    end 
  end


  always @(posedge clk) begin
    if(N2184) begin
      packet_ram_5__0_ <= N2185;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__63_ <= N2183;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__62_ <= N2182;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__61_ <= N2181;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__60_ <= N2180;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__59_ <= N2179;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__58_ <= N2178;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__57_ <= N2177;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__56_ <= N2176;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__55_ <= N2175;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__54_ <= N2174;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__53_ <= N2173;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__52_ <= N2172;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__51_ <= N2171;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__50_ <= N2170;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__49_ <= N2169;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__48_ <= N2168;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__47_ <= N2167;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__46_ <= N2166;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__45_ <= N2165;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__44_ <= N2164;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__43_ <= N2163;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__42_ <= N2162;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__41_ <= N2161;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__40_ <= N2160;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__39_ <= N2159;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__38_ <= N2158;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__37_ <= N2157;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__36_ <= N2156;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__35_ <= N2155;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__34_ <= N2154;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__33_ <= N2153;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__32_ <= N2152;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__31_ <= N2151;
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      packet_ram_4__30_ <= N2150;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__29_ <= N2148;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__28_ <= N2147;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__27_ <= N2146;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__26_ <= N2145;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__25_ <= N2144;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__24_ <= N2143;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__23_ <= N2142;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__22_ <= N2141;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__21_ <= N2140;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__20_ <= N2139;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__19_ <= N2138;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__18_ <= N2137;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__17_ <= N2136;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__16_ <= N2135;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__15_ <= N2134;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__14_ <= N2133;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__13_ <= N2132;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__12_ <= N2131;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__11_ <= N2130;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__10_ <= N2129;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__9_ <= N2128;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__8_ <= N2127;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__7_ <= N2126;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__6_ <= N2125;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__5_ <= N2124;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__4_ <= N2123;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__3_ <= N2122;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__2_ <= N2121;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__1_ <= N2120;
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      packet_ram_4__0_ <= N2119;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__63_ <= N2117;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__62_ <= N2116;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__61_ <= N2115;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__60_ <= N2114;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__59_ <= N2113;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__58_ <= N2112;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__57_ <= N2111;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__56_ <= N2110;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__55_ <= N2109;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__54_ <= N2108;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__53_ <= N2107;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__52_ <= N2106;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__51_ <= N2105;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__50_ <= N2104;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__49_ <= N2103;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__48_ <= N2102;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__47_ <= N2101;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__46_ <= N2100;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__45_ <= N2099;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__44_ <= N2098;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__43_ <= N2097;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__42_ <= N2096;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__41_ <= N2095;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__40_ <= N2094;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__39_ <= N2093;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__38_ <= N2092;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__37_ <= N2091;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__36_ <= N2090;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__35_ <= N2089;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__34_ <= N2088;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__33_ <= N2087;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__32_ <= N2086;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__31_ <= N2085;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__30_ <= N2084;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__29_ <= N2083;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__28_ <= N2082;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__27_ <= N2081;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__26_ <= N2080;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__25_ <= N2079;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__24_ <= N2078;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__23_ <= N2077;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__22_ <= N2076;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__21_ <= N2075;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__20_ <= N2074;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__19_ <= N2073;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__18_ <= N2072;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__17_ <= N2071;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__16_ <= N2070;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__15_ <= N2069;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__14_ <= N2068;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__13_ <= N2067;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__12_ <= N2066;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__11_ <= N2065;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__10_ <= N2064;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__9_ <= N2063;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__8_ <= N2062;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__7_ <= N2061;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__6_ <= N2060;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__5_ <= N2059;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__4_ <= N2058;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__3_ <= N2057;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__2_ <= N2056;
    end 
  end


  always @(posedge clk) begin
    if(N2054) begin
      packet_ram_3__1_ <= N2055;
    end 
  end


  always @(posedge clk) begin
    if(N2052) begin
      packet_ram_3__0_ <= N2053;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__63_ <= N2051;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__62_ <= N2050;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__61_ <= N2049;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__60_ <= N2048;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__59_ <= N2047;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__58_ <= N2046;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__57_ <= N2045;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__56_ <= N2044;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__55_ <= N2043;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__54_ <= N2042;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__53_ <= N2041;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__52_ <= N2040;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__51_ <= N2039;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__50_ <= N2038;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__49_ <= N2037;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__48_ <= N2036;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__47_ <= N2035;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__46_ <= N2034;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      packet_ram_2__45_ <= N2033;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__44_ <= N2031;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__43_ <= N2030;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__42_ <= N2029;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__41_ <= N2028;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__40_ <= N2027;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__39_ <= N2026;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__38_ <= N2025;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__37_ <= N2024;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__36_ <= N2023;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__35_ <= N2022;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__34_ <= N2021;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__33_ <= N2020;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__32_ <= N2019;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__31_ <= N2018;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__30_ <= N2017;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__29_ <= N2016;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__28_ <= N2015;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__27_ <= N2014;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__26_ <= N2013;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__25_ <= N2012;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__24_ <= N2011;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__23_ <= N2010;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__22_ <= N2009;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__21_ <= N2008;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__20_ <= N2007;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__19_ <= N2006;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__18_ <= N2005;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__17_ <= N2004;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__16_ <= N2003;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__15_ <= N2002;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__14_ <= N2001;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__13_ <= N2000;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__12_ <= N1999;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__11_ <= N1998;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__10_ <= N1997;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__9_ <= N1996;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__8_ <= N1995;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__7_ <= N1994;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__6_ <= N1993;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__5_ <= N1992;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__4_ <= N1991;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__3_ <= N1990;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__2_ <= N1989;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__1_ <= N1988;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      packet_ram_2__0_ <= N1987;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__63_ <= N1985;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__62_ <= N1984;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__61_ <= N1983;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__60_ <= N1982;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__59_ <= N1981;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__58_ <= N1980;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__57_ <= N1979;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__56_ <= N1978;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__55_ <= N1977;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__54_ <= N1976;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__53_ <= N1975;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__52_ <= N1974;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__51_ <= N1973;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__50_ <= N1972;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__49_ <= N1971;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__48_ <= N1970;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__47_ <= N1969;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__46_ <= N1968;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__45_ <= N1967;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__44_ <= N1966;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__43_ <= N1965;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__42_ <= N1964;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__41_ <= N1963;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__40_ <= N1962;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__39_ <= N1961;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__38_ <= N1960;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__37_ <= N1959;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__36_ <= N1958;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__35_ <= N1957;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__34_ <= N1956;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__33_ <= N1955;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__32_ <= N1954;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__31_ <= N1953;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__30_ <= N1952;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__29_ <= N1951;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__28_ <= N1950;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__27_ <= N1949;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__26_ <= N1948;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__25_ <= N1947;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__24_ <= N1946;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__23_ <= N1945;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__22_ <= N1944;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__21_ <= N1943;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__20_ <= N1942;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__19_ <= N1941;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__18_ <= N1940;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__17_ <= N1939;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__16_ <= N1938;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__15_ <= N1937;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__14_ <= N1936;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__13_ <= N1935;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__12_ <= N1934;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__11_ <= N1933;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__10_ <= N1932;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__9_ <= N1931;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__8_ <= N1930;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__7_ <= N1929;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__6_ <= N1928;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__5_ <= N1927;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__4_ <= N1926;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__3_ <= N1925;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__2_ <= N1924;
    end 
  end


  always @(posedge clk) begin
    if(N1922) begin
      packet_ram_1__1_ <= N1923;
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      packet_ram_1__0_ <= N1921;
    end 
  end


  always @(posedge clk) begin
    if(N1856) begin
      io_scr_req_bits_data[63] <= N1919;
    end 
  end


  always @(posedge clk) begin
    if(N1856) begin
      io_scr_req_bits_data[62] <= N1918;
    end 
  end


  always @(posedge clk) begin
    if(N1856) begin
      io_scr_req_bits_data[61] <= N1917;
    end 
  end


  always @(posedge clk) begin
    if(N1856) begin
      io_scr_req_bits_data[60] <= N1916;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[59] <= N1915;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[58] <= N1914;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[57] <= N1913;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[56] <= N1912;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[55] <= N1911;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[54] <= N1910;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[53] <= N1909;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[52] <= N1908;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[51] <= N1907;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[50] <= N1906;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[49] <= N1905;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[48] <= N1904;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[47] <= N1903;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[46] <= N1902;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[45] <= N1901;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[44] <= N1900;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[43] <= N1899;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[42] <= N1898;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[41] <= N1897;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[40] <= N1896;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[39] <= N1895;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[38] <= N1894;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[37] <= N1893;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[36] <= N1892;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[35] <= N1891;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[34] <= N1890;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[33] <= N1889;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[32] <= N1888;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[31] <= N1887;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[30] <= N1886;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[29] <= N1885;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[28] <= N1884;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[27] <= N1883;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[26] <= N1882;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[25] <= N1881;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[24] <= N1880;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[23] <= N1879;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[22] <= N1878;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[21] <= N1877;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[20] <= N1876;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[19] <= N1875;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[18] <= N1874;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[17] <= N1873;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[16] <= N1872;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[15] <= N1871;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[14] <= N1870;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[13] <= N1869;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[12] <= N1868;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[11] <= N1867;
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      io_scr_req_bits_data[10] <= N1866;
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      io_scr_req_bits_data[9] <= N1865;
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      io_scr_req_bits_data[8] <= N1864;
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      io_scr_req_bits_data[7] <= N1863;
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      io_scr_req_bits_data[6] <= N1862;
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      io_scr_req_bits_data[5] <= N1861;
    end 
  end


  always @(posedge clk) begin
    if(N1858) begin
      io_scr_req_bits_data[4] <= N1859;
    end 
  end


  always @(posedge clk) begin
    if(N1856) begin
      io_scr_req_bits_data[3] <= N1857;
    end 
  end


  always @(posedge clk) begin
    if(N1854) begin
      io_scr_req_bits_data[2] <= N1855;
    end 
  end


  always @(posedge clk) begin
    if(N1852) begin
      io_scr_req_bits_data[1] <= N1853;
    end 
  end


  always @(posedge clk) begin
    if(N1850) begin
      io_scr_req_bits_data[0] <= N1851;
    end 
  end


  always @(posedge clk) begin
    if(N136) begin
      state[2] <= N139;
    end 
  end


  always @(posedge clk) begin
    if(N136) begin
      state[1] <= N138;
    end 
  end


  always @(posedge clk) begin
    if(N136) begin
      state[0] <= N137;
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      cmd[3] <= rx_shifter_in_3;
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      cmd[2] <= rx_shifter_in_2;
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      cmd[1] <= rx_shifter_in_1;
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      cmd[0] <= rx_shifter_in_0;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[12] <= N158;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[11] <= N157;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[10] <= N156;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[9] <= N155;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[8] <= N154;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[7] <= N153;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[6] <= N152;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[5] <= N151;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[4] <= N150;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[3] <= N149;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[2] <= N148;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[1] <= N147;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      rx_word_count[0] <= N146;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      T77[1] <= N145;
    end 
  end


  always @(posedge clk) begin
    if(N143) begin
      T77[0] <= N144;
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[11] <= T29[11];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[10] <= T29[10];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[9] <= T29[9];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[8] <= T29[8];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[7] <= T29[7];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[6] <= T29[6];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[5] <= T29[5];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[4] <= T29[4];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T214[3] <= T29[3];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T53[2] <= T29[2];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T53[1] <= T29[1];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      T53[0] <= T29[0];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[47] <= io_host_in_bits[15];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[46] <= io_host_in_bits[14];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[45] <= io_host_in_bits[13];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[44] <= io_host_in_bits[12];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[43] <= io_host_in_bits[11];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[42] <= io_host_in_bits[10];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[41] <= io_host_in_bits[9];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[40] <= io_host_in_bits[8];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[39] <= io_host_in_bits[7];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[38] <= io_host_in_bits[6];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[37] <= io_host_in_bits[5];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[36] <= io_host_in_bits[4];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[35] <= io_host_in_bits[3];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[34] <= io_host_in_bits[2];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[33] <= io_host_in_bits[1];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[32] <= io_host_in_bits[0];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[31] <= rx_shifter_in[47];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[30] <= rx_shifter_in[46];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[29] <= rx_shifter_in[45];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[28] <= rx_shifter_in[44];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[27] <= rx_shifter_in[43];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[26] <= rx_shifter_in[42];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[25] <= rx_shifter_in[41];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[24] <= rx_shifter_in[40];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[23] <= rx_shifter_in[39];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[22] <= rx_shifter_in[38];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[21] <= rx_shifter_in[37];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[20] <= rx_shifter_in[36];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[19] <= rx_shifter_in[35];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[18] <= rx_shifter_in[34];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[17] <= rx_shifter_in[33];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in[16] <= rx_shifter_in[32];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[11] <= rx_shifter_in[31];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[10] <= rx_shifter_in[30];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[9] <= rx_shifter_in[29];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[8] <= rx_shifter_in[28];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[7] <= rx_shifter_in[27];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[6] <= rx_shifter_in[26];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[5] <= rx_shifter_in[25];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[4] <= rx_shifter_in[24];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[3] <= rx_shifter_in[23];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[2] <= rx_shifter_in[22];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[1] <= rx_shifter_in[21];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      T29[0] <= rx_shifter_in[20];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in_3 <= rx_shifter_in[19];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in_2 <= rx_shifter_in[18];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in_1 <= rx_shifter_in[17];
    end 
  end


  always @(posedge clk) begin
    if(T61) begin
      rx_shifter_in_0 <= rx_shifter_in[16];
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[36] <= N202;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[35] <= N201;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[34] <= N200;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[33] <= N199;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[32] <= N198;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[31] <= N197;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[30] <= N196;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[29] <= N195;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[28] <= N194;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[27] <= N193;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      init_addr[26] <= N192;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[25] <= N191;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[24] <= N190;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[23] <= N189;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[22] <= N188;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[21] <= N187;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[20] <= N186;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[19] <= N185;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[18] <= N184;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[17] <= N183;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[16] <= N182;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[15] <= N181;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[14] <= N180;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[13] <= N179;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[12] <= N178;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[11] <= N177;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[10] <= N176;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_mem_acquire_bits_addr_block[9] <= N175;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_cpu_0_csr_req_bits_addr[11] <= N174;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_cpu_0_csr_req_bits_addr[10] <= N173;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_cpu_0_csr_req_bits_addr[9] <= N172;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_cpu_0_csr_req_bits_addr[8] <= N171;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_cpu_0_csr_req_bits_addr[7] <= N170;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_cpu_0_csr_req_bits_addr[6] <= N169;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_scr_req_bits_addr[5] <= N168;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_scr_req_bits_addr[4] <= N167;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_scr_req_bits_addr[3] <= N166;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_scr_req_bits_addr[2] <= N165;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_scr_req_bits_addr[1] <= N164;
    end 
  end


  always @(posedge clk) begin
    if(N162) begin
      io_scr_req_bits_addr[0] <= N163;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[12] <= N221;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[11] <= N220;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[10] <= N219;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[9] <= N218;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[8] <= N217;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[7] <= N216;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[6] <= N215;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[5] <= N214;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[4] <= N213;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[3] <= N212;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[2] <= N211;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[1] <= N210;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_word_count[0] <= N209;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_subword_count[1] <= N208;
    end 
  end


  always @(posedge clk) begin
    if(N206) begin
      tx_subword_count[0] <= N207;
    end 
  end


  always @(posedge clk) begin
    if(N224) begin
      T154[2] <= N226;
    end 
  end


  always @(posedge clk) begin
    if(N224) begin
      T154[1] <= N225;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[8] <= N239;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[7] <= N238;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[6] <= N237;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[5] <= N236;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[4] <= N235;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[3] <= N234;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[2] <= N233;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[1] <= N232;
    end 
  end


  always @(posedge clk) begin
    if(N230) begin
      pos[0] <= N231;
    end 
  end


  always @(posedge clk) begin
    if(N2384) begin
      io_cpu_0_reset <= N2385;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[63] <= N2453;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[62] <= N2452;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[61] <= N2451;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[60] <= N2450;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[59] <= N2449;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[58] <= N2448;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[57] <= N2447;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[56] <= N2446;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[55] <= N2445;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[54] <= N2444;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[53] <= N2443;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[52] <= N2442;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[51] <= N2441;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[50] <= N2440;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[49] <= N2439;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[48] <= N2438;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[47] <= N2437;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[46] <= N2436;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[45] <= N2435;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[44] <= N2434;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[43] <= N2433;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[42] <= N2432;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[41] <= N2431;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[40] <= N2430;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[39] <= N2429;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[38] <= N2428;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[37] <= N2427;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[36] <= N2426;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[35] <= N2425;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[34] <= N2424;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[33] <= N2423;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[32] <= N2422;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[31] <= N2421;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[30] <= N2420;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[29] <= N2419;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[28] <= N2418;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[27] <= N2417;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[26] <= N2416;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[25] <= N2415;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[24] <= N2414;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[23] <= N2413;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[22] <= N2412;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[21] <= N2411;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[20] <= N2410;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[19] <= N2409;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[18] <= N2408;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[17] <= N2407;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[16] <= N2406;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[15] <= N2405;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[14] <= N2404;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[13] <= N2403;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[12] <= N2402;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[11] <= N2401;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[10] <= N2400;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[9] <= N2399;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[8] <= N2398;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[7] <= N2397;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[6] <= N2396;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[5] <= N2395;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[4] <= N2394;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[3] <= N2393;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[2] <= N2392;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[1] <= N2391;
    end 
  end


  always @(posedge clk) begin
    if(N2389) begin
      csrReadData[0] <= N2390;
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[23] <= rx_shifter_in[23];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[22] <= rx_shifter_in[22];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[21] <= rx_shifter_in[21];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[20] <= rx_shifter_in[20];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[19] <= rx_shifter_in[19];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[18] <= rx_shifter_in[18];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[17] <= rx_shifter_in[17];
    end 
  end


  always @(posedge clk) begin
    if(T21) begin
      tx_header[16] <= rx_shifter_in[16];
    end 
  end

  assign N2504 = ~cmd[1];
  assign N2505 = ~cmd[0];
  assign N2506 = cmd[2] | cmd[3];
  assign N2507 = N2504 | N2506;
  assign N2508 = N2505 | N2507;
  assign io_cpu_0_csr_req_bits_rw = ~N2508;
  assign N2510 = cmd[2] | cmd[3];
  assign N2511 = N2504 | N2510;
  assign N2512 = N2505 | N2511;
  assign io_scr_req_bits_rw = ~N2512;
  assign N2514 = ~state[1];
  assign N2515 = ~state[0];
  assign N2516 = N2514 | state[2];
  assign N2517 = N2515 | N2516;
  assign N2518 = ~N2517;
  assign N2519 = ~state[2];
  assign N2520 = state[1] | N2519;
  assign N2521 = state[0] | N2520;
  assign N2522 = ~N2521;
  assign N2523 = cmd[2] | cmd[3];
  assign N2524 = cmd[1] | N2523;
  assign N2525 = N2505 | N2524;
  assign N2526 = ~N2525;
  assign N2527 = tx_word_count[11] | tx_word_count[12];
  assign N2528 = tx_word_count[10] | N2527;
  assign N2529 = tx_word_count[9] | N2528;
  assign N2530 = tx_word_count[8] | N2529;
  assign N2531 = tx_word_count[7] | N2530;
  assign N2532 = tx_word_count[6] | N2531;
  assign N2533 = tx_word_count[5] | N2532;
  assign N2534 = tx_word_count[4] | N2533;
  assign N2535 = tx_word_count[3] | N2534;
  assign N2536 = tx_word_count[2] | N2535;
  assign N2537 = tx_word_count[1] | N2536;
  assign N2538 = tx_word_count[0] | N2537;
  assign N2539 = ~N2538;
  assign N2540 = rx_cmd[2] | rx_cmd[3];
  assign N2541 = rx_cmd[1] | N2540;
  assign N2542 = rx_cmd[0] | N2541;
  assign N2543 = ~N2542;
  assign N2544 = cmd[2] | cmd[3];
  assign N2545 = N2504 | N2544;
  assign N2546 = cmd[0] | N2545;
  assign N2547 = ~N2546;
  assign N2548 = cmd[2] | cmd[3];
  assign N2549 = N2504 | N2548;
  assign N2550 = N2505 | N2549;
  assign N2551 = ~N2550;
  assign N2552 = state[1] | state[2];
  assign N2553 = state[0] | N2552;
  assign N2554 = ~N2553;
  assign N2555 = cmd[2] | cmd[3];
  assign N2556 = cmd[1] | N2555;
  assign N2557 = cmd[0] | N2556;
  assign N2558 = ~N2557;
  assign N2559 = pos[7] | pos[8];
  assign N2560 = pos[6] | N2559;
  assign N2561 = pos[5] | N2560;
  assign N2562 = pos[4] | N2561;
  assign N2563 = pos[3] | N2562;
  assign N2564 = pos[2] | N2563;
  assign N2565 = pos[1] | N2564;
  assign N2566 = pos[0] | N2565;
  assign N2567 = cmd[2] | cmd[3];
  assign N2568 = cmd[1] | N2567;
  assign N2569 = cmd[0] | N2568;
  assign N2570 = ~N2569;
  assign N2571 = ~pos[0];
  assign N2572 = pos[7] | pos[8];
  assign N2573 = pos[6] | N2572;
  assign N2574 = pos[5] | N2573;
  assign N2575 = pos[4] | N2574;
  assign N2576 = pos[3] | N2575;
  assign N2577 = pos[2] | N2576;
  assign N2578 = pos[1] | N2577;
  assign N2579 = N2571 | N2578;
  assign N2580 = ~N2579;
  assign N2581 = cmd[2] | cmd[3];
  assign N2582 = cmd[1] | N2581;
  assign N2583 = cmd[0] | N2582;
  assign N2584 = ~N2583;
  assign N2585 = pos[7] | pos[8];
  assign N2586 = pos[6] | N2585;
  assign N2587 = pos[5] | N2586;
  assign N2588 = pos[4] | N2587;
  assign N2589 = pos[3] | N2588;
  assign N2590 = pos[2] | N2589;
  assign N2591 = pos[1] | N2590;
  assign N2592 = N2571 | N2591;
  assign N2593 = ~N2592;
  assign N2594 = ~rx_cmd[0];
  assign N2595 = rx_cmd[2] | rx_cmd[3];
  assign N2596 = rx_cmd[1] | N2595;
  assign N2597 = N2594 | N2596;
  assign N2598 = ~N2597;
  assign N2599 = state[1] & state[2];
  assign io_host_out_valid = state[0] & N2599;
  assign N2601 = ~T77[1];
  assign N2602 = ~T77[0];
  assign N2603 = rx_word_count[11] | rx_word_count[12];
  assign N2604 = rx_word_count[10] | N2603;
  assign N2605 = rx_word_count[9] | N2604;
  assign N2606 = rx_word_count[8] | N2605;
  assign N2607 = rx_word_count[7] | N2606;
  assign N2608 = rx_word_count[6] | N2607;
  assign N2609 = rx_word_count[5] | N2608;
  assign N2610 = rx_word_count[4] | N2609;
  assign N2611 = rx_word_count[3] | N2610;
  assign N2612 = rx_word_count[2] | N2611;
  assign N2613 = rx_word_count[1] | N2612;
  assign N2614 = rx_word_count[0] | N2613;
  assign N2615 = N2601 | N2614;
  assign N2616 = N2602 | N2615;
  assign N2617 = ~N2616;
  assign N2618 = cmd[2] | cmd[3];
  assign N2619 = N2504 | N2618;
  assign N2620 = N2505 | N2619;
  assign N2621 = ~N2620;
  assign N2622 = state[1] | N2519;
  assign N2623 = state[0] | N2622;
  assign N2624 = ~N2623;
  assign N2625 = state[1] | state[2];
  assign N2626 = state[0] | N2625;
  assign io_host_in_ready = ~N2626;
  assign N2628 = ~rx_cmd[1];
  assign N2629 = rx_cmd[2] | rx_cmd[3];
  assign N2630 = N2628 | N2629;
  assign N2631 = rx_cmd[0] | N2630;
  assign N2632 = ~N2631;
  assign N2633 = rx_cmd[2] | rx_cmd[3];
  assign N2634 = N2628 | N2633;
  assign N2635 = N2594 | N2634;
  assign N2636 = ~N2635;
  assign N2637 = N2514 | state[2];
  assign N2638 = N2515 | N2637;
  assign N2639 = ~N2638;
  assign N2640 = T77[0] & T77[1];
  assign N2641 = ~rx_shifter_in_0;
  assign N2642 = rx_shifter_in_2 | rx_shifter_in_3;
  assign N2643 = rx_shifter_in_1 | N2642;
  assign N2644 = N2641 | N2643;
  assign N2645 = ~rx_shifter_in_1;
  assign N2646 = rx_shifter_in_2 | rx_shifter_in_3;
  assign N2647 = N2645 | N2646;
  assign N2648 = N2641 | N2647;
  assign N2649 = rx_word_count[1] | rx_word_count[2];
  assign N2650 = rx_word_count[0] | N2649;
  assign N2651 = ~N2650;
  assign N2652 = N2514 | N2519;
  assign N2653 = state[0] | N2652;
  assign N2654 = ~N2653;
  assign N2655 = state[1] | N2519;
  assign N2656 = N2515 | N2655;
  assign N2657 = ~N2656;
  assign N2658 = state[1] | N2519;
  assign N2659 = N2515 | N2658;
  assign N2660 = ~N2659;
  assign N2661 = rx_word_count[11] | rx_word_count[12];
  assign N2662 = rx_word_count[10] | N2661;
  assign N2663 = rx_word_count[9] | N2662;
  assign N2664 = rx_word_count[8] | N2663;
  assign N2665 = rx_word_count[7] | N2664;
  assign N2666 = rx_word_count[6] | N2665;
  assign N2667 = rx_word_count[5] | N2666;
  assign N2668 = rx_word_count[4] | N2667;
  assign N2669 = rx_word_count[3] | N2668;
  assign N2670 = rx_word_count[2] | N2669;
  assign N2671 = rx_word_count[1] | N2670;
  assign N2672 = rx_word_count[0] | N2671;
  assign N2673 = ~N2672;
  assign N2674 = state[1] | N2519;
  assign N2675 = N2515 | N2674;
  assign N2676 = ~N2675;
  assign N2677 = state[1] & state[2];
  assign N2678 = state[0] & N2677;
  assign N2679 = T154[1] & T154[2];
  assign N2680 = rx_word_count[11] | rx_word_count[12];
  assign N2681 = rx_word_count[10] | N2680;
  assign N2682 = rx_word_count[9] | N2681;
  assign N2683 = rx_word_count[8] | N2682;
  assign N2684 = rx_word_count[7] | N2683;
  assign N2685 = rx_word_count[6] | N2684;
  assign N2686 = rx_word_count[5] | N2685;
  assign N2687 = rx_word_count[4] | N2686;
  assign N2688 = rx_word_count[3] | N2687;
  assign N2689 = rx_word_count[2] | N2688;
  assign N2690 = rx_word_count[1] | N2689;
  assign N2691 = rx_word_count[0] | N2690;
  assign N2692 = ~N2691;
  assign N2693 = ~io_cpu_0_csr_req_bits_addr[10];
  assign N2694 = ~io_cpu_0_csr_req_bits_addr[9];
  assign N2695 = ~io_cpu_0_csr_req_bits_addr[8];
  assign N2696 = ~io_cpu_0_csr_req_bits_addr[7];
  assign N2697 = ~io_scr_req_bits_addr[1];
  assign N2698 = N2693 | io_cpu_0_csr_req_bits_addr[11];
  assign N2699 = N2694 | N2698;
  assign N2700 = N2695 | N2699;
  assign N2701 = N2696 | N2700;
  assign N2702 = io_cpu_0_csr_req_bits_addr[6] | N2701;
  assign N2703 = io_scr_req_bits_addr[5] | N2702;
  assign N2704 = io_scr_req_bits_addr[4] | N2703;
  assign N2705 = io_scr_req_bits_addr[3] | N2704;
  assign N2706 = io_scr_req_bits_addr[2] | N2705;
  assign N2707 = N2697 | N2706;
  assign N2708 = io_scr_req_bits_addr[0] | N2707;
  assign N2709 = ~N2708;
  assign N2710 = N2693 | io_cpu_0_csr_req_bits_addr[11];
  assign N2711 = N2694 | N2710;
  assign N2712 = N2695 | N2711;
  assign N2713 = N2696 | N2712;
  assign N2714 = io_cpu_0_csr_req_bits_addr[6] | N2713;
  assign N2715 = io_scr_req_bits_addr[5] | N2714;
  assign N2716 = io_scr_req_bits_addr[4] | N2715;
  assign N2717 = io_scr_req_bits_addr[3] | N2716;
  assign N2718 = io_scr_req_bits_addr[2] | N2717;
  assign N2719 = N2697 | N2718;
  assign N2720 = io_scr_req_bits_addr[0] | N2719;
  assign N2721 = tx_subword_count[0] & tx_subword_count[1];
  assign N2722 = state[1] | N2519;
  assign N2723 = state[0] | N2722;
  assign N2724 = ~N2723;
  assign N2725 = state[1] | N2519;
  assign N2726 = N2515 | N2725;
  assign N2727 = ~N2726;
  assign N2728 = N2514 | state[2];
  assign N2729 = state[0] | N2728;
  assign N2730 = ~N2729;
  assign N2731 = state[1] | state[2];
  assign N2732 = N2515 | N2731;
  assign N2733 = ~N2732;
  assign N2734 = state[1] | state[2];
  assign N2735 = N2515 | N2734;
  assign N2736 = ~N2735;
  assign N2737 = io_mem_acquire_bits_addr_block[17] | io_mem_acquire_bits_addr_block[18];
  assign N2738 = ~N2737;
  assign N2739 = N2514 | state[2];
  assign N2740 = state[0] | N2739;
  assign N2741 = ~N2740;
  assign N2742 = state[1] | state[2];
  assign N2743 = N2515 | N2742;
  assign N2744 = ~N2743;
  assign N2745 = io_mem_acquire_bits_addr_block[17] & io_mem_acquire_bits_addr_block[18];
  assign N2746 = cmd[2] | cmd[3];
  assign N2747 = N2504 | N2746;
  assign N2748 = N2505 | N2747;
  assign N2749 = ~N2748;
  assign N2750 = cmd[2] | cmd[3];
  assign N2751 = cmd[1] | N2750;
  assign N2752 = cmd[0] | N2751;
  assign N2753 = ~N2752;
  assign N2754 = cmd[2] | cmd[3];
  assign N2755 = N2504 | N2754;
  assign N2756 = cmd[0] | N2755;
  assign N2757 = ~N2756;
  assign N2758 = T53[1] | T53[2];
  assign N2759 = T53[0] | N2758;
  assign N2760 = io_scr_req_bits_addr[1] | io_scr_req_bits_addr[2];
  assign N2761 = io_scr_req_bits_addr[0] | N2760;
  assign N2762 = ~T53[0];
  assign N2763 = T214[10] | T214[11];
  assign N2764 = T214[9] | N2763;
  assign N2765 = T214[8] | N2764;
  assign N2766 = T214[7] | N2765;
  assign N2767 = T214[6] | N2766;
  assign N2768 = T214[5] | N2767;
  assign N2769 = T214[4] | N2768;
  assign N2770 = T214[3] | N2769;
  assign N2771 = T53[2] | N2770;
  assign N2772 = T53[1] | N2771;
  assign N2773 = N2762 | N2772;
  assign N2774 = cmd[2] | cmd[3];
  assign N2775 = cmd[1] | N2774;
  assign N2776 = cmd[0] | N2775;
  assign N2777 = ~N2776;
  assign N2778 = cmd[2] | cmd[3];
  assign N2779 = cmd[1] | N2778;
  assign N2780 = N2505 | N2779;
  assign N2781 = ~N2780;
  assign N2782 = cmd[2] | cmd[3];
  assign N2783 = N2504 | N2782;
  assign N2784 = cmd[0] | N2783;
  assign N2785 = ~N2784;
  assign N2786 = cmd[2] | cmd[3];
  assign N2787 = N2504 | N2786;
  assign N2788 = N2505 | N2787;
  assign N2789 = ~N2788;
  assign T142 = rx_word_count[2:0] - 1'b1;
  assign T25 = { rx_word_count, T77 } + 1'b1;
  assign T50 = { init_addr, io_mem_acquire_bits_addr_block[25:9], io_cpu_0_csr_req_bits_addr[11:6], io_scr_req_bits_addr } + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign T51 = { init_addr, io_mem_acquire_bits_addr_block[25:9], io_cpu_0_csr_req_bits_addr[11:6], io_scr_req_bits_addr } + { 1'b1, 1'b0, 1'b0, 1'b0 };
  assign packet_ram_raddr = tx_word_count[2:0] - 1'b1;
  assign T59 = { tx_word_count, tx_subword_count } + 1'b1;
  assign T82 = T154 + 1'b1;
  assign T98 = pos - 1'b1;
  assign T99 = pos - 1'b1;
  assign N115 = io_mem_grant_bits_addr_beat[0] & io_mem_grant_bits_addr_beat[1];
  assign N114 = N0 & io_mem_grant_bits_addr_beat[1];
  assign N0 = ~io_mem_grant_bits_addr_beat[0];
  assign N113 = io_mem_grant_bits_addr_beat[0] & N1;
  assign N1 = ~io_mem_grant_bits_addr_beat[1];
  assign N112 = N2 & N3;
  assign N2 = ~io_mem_grant_bits_addr_beat[0];
  assign N3 = ~io_mem_grant_bits_addr_beat[1];
  assign N702 = io_mem_grant_bits_addr_beat[0] & io_mem_grant_bits_addr_beat[1];
  assign N570 = N4 & io_mem_grant_bits_addr_beat[1];
  assign N4 = ~io_mem_grant_bits_addr_beat[0];
  assign N438 = io_mem_grant_bits_addr_beat[0] & N5;
  assign N5 = ~io_mem_grant_bits_addr_beat[1];
  assign N306 = N6 & N7;
  assign N6 = ~io_mem_grant_bits_addr_beat[0];
  assign N7 = ~io_mem_grant_bits_addr_beat[1];
  assign N2790 = T142[0] & T142[1];
  assign N1309 = N2790 & T142[2];
  assign N2791 = N8 & T142[1];
  assign N8 = ~T142[0];
  assign N1308 = N2791 & T142[2];
  assign N2792 = T142[0] & N9;
  assign N9 = ~T142[1];
  assign N1307 = N2792 & T142[2];
  assign N2793 = N10 & N11;
  assign N10 = ~T142[0];
  assign N11 = ~T142[1];
  assign N1306 = N2793 & T142[2];
  assign N2794 = T142[0] & T142[1];
  assign N1305 = N2794 & N12;
  assign N12 = ~T142[2];
  assign N2795 = N13 & T142[1];
  assign N13 = ~T142[0];
  assign N1304 = N2795 & N14;
  assign N14 = ~T142[2];
  assign N2796 = T142[0] & N15;
  assign N15 = ~T142[1];
  assign N1303 = N2796 & N16;
  assign N16 = ~T142[2];
  assign N2797 = N17 & N18;
  assign N17 = ~T142[0];
  assign N18 = ~T142[1];
  assign N1302 = N2797 & N19;
  assign N19 = ~T142[2];
  assign T15 = (N20)? { 1'b0, 1'b1, 1'b1 } : 
               (N21)? T16 : 1'b0;
  assign N20 = N2543;
  assign N21 = N2542;
  assign T16[2:1] = (N22)? { 1'b1, 1'b0 } : 
                    (N23)? { T17[2:2], T17[2:2] } : 1'b0;
  assign N22 = N2598;
  assign N23 = T16[0];
  assign rx_cmd = (N24)? { rx_shifter_in_3, rx_shifter_in_2, rx_shifter_in_1, rx_shifter_in_0 } : 
                  (N25)? cmd : 1'b0;
  assign N24 = N2692;
  assign N25 = N2691;
  assign T212 = (N26)? { T214, T53 } : 
                (N27)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = T32;
  assign N27 = N64;
  assign nack = (N28)? bad_mem_packet : 
                (N29)? T39 : 1'b0;
  assign N28 = T54;
  assign N29 = N65;
  assign T39 = (N30)? N2773 : 
               (N31)? 1'b1 : 1'b0;
  assign N30 = T41;
  assign N31 = N66;
  assign T67 = (N32)? T72 : 
               (N33)? T68 : 1'b0;
  assign N32 = N2673;
  assign N33 = N2672;
  assign io_mem_acquire_bits_data = (N34)? T152 : 
                                    (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34 = N2526;
  assign N35 = N2525;
  assign io_mem_acquire_bits_addr_beat = (N36)? T154 : 
                                         (N35)? { 1'b0, 1'b0 } : 1'b0;
  assign N36 = io_mem_acquire_bits_a_type[1];
  assign tx_data = (N37)? { init_addr, io_mem_acquire_bits_addr_block[25:9], io_cpu_0_csr_req_bits_addr[11:6], io_scr_req_bits_addr, tx_header, T212, 1'b0, 1'b1, 1'b0, tx_header_0 } : 
                   (N38)? T195 : 1'b0;
  assign N37 = N2539;
  assign N38 = N2538;
  assign T195 = (N39)? csrReadData : 
                (N40)? T196 : 1'b0;
  assign N39 = T200;
  assign N40 = N95;
  assign { N123, N122, N121, N120, N119, N118, N117, N116 } = (N41)? { N115, N115, N114, N114, N113, N113, N112, N112 } : 
                                                              (N42)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = T2;
  assign N42 = N111;
  assign N136 = (N43)? 1'b1 : 
                (N2454)? 1'b1 : 
                (N2457)? 1'b1 : 
                (N2460)? 1'b1 : 
                (N2463)? 1'b1 : 
                (N2466)? 1'b1 : 
                (N2469)? 1'b1 : 
                (N2472)? 1'b1 : 
                (N2475)? 1'b1 : 
                (N2478)? 1'b1 : 
                (N2481)? 1'b1 : 
                (N2484)? 1'b1 : 
                (N135)? 1'b0 : 1'b0;
  assign N43 = reset;
  assign { N139, N138, N137 } = (N43)? { 1'b0, 1'b0, 1'b0 } : 
                                (N2454)? { 1'b1, 1'b1, 1'b1 } : 
                                (N2457)? { 1'b0, 1'b1, 1'b0 } : 
                                (N2460)? { 1'b1, 1'b1, 1'b1 } : 
                                (N2463)? { 1'b1, 1'b1, 1'b1 } : 
                                (N2466)? { 1'b0, 1'b1, 1'b0 } : 
                                (N2469)? { 1'b0, T109[1:1], T109[1:1] } : 
                                (N2472)? { T103[2:2], T103[2:2], T103[2:2] } : 
                                (N2475)? { T91[2:2], T91[2:2], T91[2:2] } : 
                                (N2478)? { 1'b1, 1'b0, 1'b1 } : 
                                (N2481)? { 1'b1, 1'b1, 1'b0 } : 
                                (N2484)? T15 : 1'b0;
  assign N143 = (N43)? 1'b1 : 
                (N2485)? 1'b1 : 
                (N2488)? 1'b1 : 
                (N142)? 1'b0 : 1'b0;
  assign { N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144 } = (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                        (N2485)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                        (N2488)? T25 : 1'b0;
  assign N162 = (N44)? 1'b1 : 
                (N2489)? 1'b1 : 
                (N2491)? 1'b1 : 
                (N161)? 1'b0 : 1'b0;
  assign N44 = T107;
  assign { N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163 } = (N44)? T51 : 
                                                                                                                                                                                                                                                              (N2489)? T50 : 
                                                                                                                                                                                                                                                              (N2491)? { io_host_in_bits, rx_shifter_in[47:24] } : 1'b0;
  assign N206 = (N43)? 1'b1 : 
                (N2492)? 1'b1 : 
                (N2494)? 1'b1 : 
                (N205)? 1'b0 : 1'b0;
  assign { N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207 } = (N43)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                        (N2492)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                        (N2494)? T59 : 1'b0;
  assign N224 = (N43)? 1'b1 : 
                (N2496)? 1'b1 : 
                (N223)? 1'b0 : 1'b0;
  assign { N226, N225 } = (N43)? { 1'b0, 1'b0 } : 
                          (N2496)? T82 : 1'b0;
  assign N230 = (N44)? 1'b1 : 
                (N2497)? 1'b1 : 
                (N2499)? 1'b1 : 
                (N229)? 1'b0 : 1'b0;
  assign { N239, N238, N237, N236, N235, N234, N233, N232, N231 } = (N44)? T99 : 
                                                                    (N2497)? T98 : 
                                                                    (N2499)? T29[11:3] : 1'b0;
  assign { N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242 } = (N45)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N241)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign N45 = N306;
  assign { N371, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307 } = (N46)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N67)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign N46 = 1'b0;
  assign { N372, N370 } = (N46)? { 1'b1, 1'b1 } : 
                          (N67)? { N116, N117 } : 1'b0;
  assign { N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } = (N47)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N373)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign N47 = N438;
  assign { N503, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439 } = (N46)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N67)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign { N504, N502 } = (N46)? { 1'b1, 1'b1 } : 
                          (N67)? { N118, N119 } : 1'b0;
  assign { N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506 } = (N48)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N505)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign N48 = N570;
  assign { N635, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571 } = (N46)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N67)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign { N636, N634 } = (N46)? { 1'b1, 1'b1 } : 
                          (N67)? { N120, N121 } : 1'b0;
  assign { N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638 } = (N49)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N637)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign N49 = N702;
  assign { N767, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703 } = (N46)? { io_mem_grant_bits_data[0:0], io_mem_grant_bits_data[1:1], io_mem_grant_bits_data[2:2], io_mem_grant_bits_data[3:3], io_mem_grant_bits_data[4:4], io_mem_grant_bits_data[5:5], io_mem_grant_bits_data[6:6], io_mem_grant_bits_data[7:7], io_mem_grant_bits_data[8:8], io_mem_grant_bits_data[9:9], io_mem_grant_bits_data[10:10], io_mem_grant_bits_data[11:11], io_mem_grant_bits_data[12:12], io_mem_grant_bits_data[13:13], io_mem_grant_bits_data[14:14], io_mem_grant_bits_data[15:15], io_mem_grant_bits_data[16:16], io_mem_grant_bits_data[17:17], io_mem_grant_bits_data[18:18], io_mem_grant_bits_data[19:19], io_mem_grant_bits_data[20:20], io_mem_grant_bits_data[21:21], io_mem_grant_bits_data[22:22], io_mem_grant_bits_data[23:23], io_mem_grant_bits_data[24:24], io_mem_grant_bits_data[25:25], io_mem_grant_bits_data[26:26], io_mem_grant_bits_data[27:27], io_mem_grant_bits_data[28:28], io_mem_grant_bits_data[29:29], io_mem_grant_bits_data[30:30], io_mem_grant_bits_data[31:31], io_mem_grant_bits_data[32:32], io_mem_grant_bits_data[33:33], io_mem_grant_bits_data[34:34], io_mem_grant_bits_data[35:35], io_mem_grant_bits_data[36:36], io_mem_grant_bits_data[37:37], io_mem_grant_bits_data[38:38], io_mem_grant_bits_data[39:39], io_mem_grant_bits_data[40:40], io_mem_grant_bits_data[41:41], io_mem_grant_bits_data[42:42], io_mem_grant_bits_data[43:43], io_mem_grant_bits_data[44:44], io_mem_grant_bits_data[45:45], io_mem_grant_bits_data[46:46], io_mem_grant_bits_data[47:47], io_mem_grant_bits_data[48:48], io_mem_grant_bits_data[49:49], io_mem_grant_bits_data[50:50], io_mem_grant_bits_data[51:51], io_mem_grant_bits_data[52:52], io_mem_grant_bits_data[53:53], io_mem_grant_bits_data[54:54], io_mem_grant_bits_data[55:55], io_mem_grant_bits_data[56:56], io_mem_grant_bits_data[57:57], io_mem_grant_bits_data[58:58], io_mem_grant_bits_data[59:59], io_mem_grant_bits_data[60:60], io_mem_grant_bits_data[61:61], io_mem_grant_bits_data[62:62], io_mem_grant_bits_data[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N67)? { io_mem_grant_bits_data[64:64], io_mem_grant_bits_data[65:65], io_mem_grant_bits_data[66:66], io_mem_grant_bits_data[67:67], io_mem_grant_bits_data[68:68], io_mem_grant_bits_data[69:69], io_mem_grant_bits_data[70:70], io_mem_grant_bits_data[71:71], io_mem_grant_bits_data[72:72], io_mem_grant_bits_data[73:73], io_mem_grant_bits_data[74:74], io_mem_grant_bits_data[75:75], io_mem_grant_bits_data[76:76], io_mem_grant_bits_data[77:77], io_mem_grant_bits_data[78:78], io_mem_grant_bits_data[79:79], io_mem_grant_bits_data[80:80], io_mem_grant_bits_data[81:81], io_mem_grant_bits_data[82:82], io_mem_grant_bits_data[83:83], io_mem_grant_bits_data[84:84], io_mem_grant_bits_data[85:85], io_mem_grant_bits_data[86:86], io_mem_grant_bits_data[87:87], io_mem_grant_bits_data[88:88], io_mem_grant_bits_data[89:89], io_mem_grant_bits_data[90:90], io_mem_grant_bits_data[91:91], io_mem_grant_bits_data[92:92], io_mem_grant_bits_data[93:93], io_mem_grant_bits_data[94:94], io_mem_grant_bits_data[95:95], io_mem_grant_bits_data[96:96], io_mem_grant_bits_data[97:97], io_mem_grant_bits_data[98:98], io_mem_grant_bits_data[99:99], io_mem_grant_bits_data[100:100], io_mem_grant_bits_data[101:101], io_mem_grant_bits_data[102:102], io_mem_grant_bits_data[103:103], io_mem_grant_bits_data[104:104], io_mem_grant_bits_data[105:105], io_mem_grant_bits_data[106:106], io_mem_grant_bits_data[107:107], io_mem_grant_bits_data[108:108], io_mem_grant_bits_data[109:109], io_mem_grant_bits_data[110:110], io_mem_grant_bits_data[111:111], io_mem_grant_bits_data[112:112], io_mem_grant_bits_data[113:113], io_mem_grant_bits_data[114:114], io_mem_grant_bits_data[115:115], io_mem_grant_bits_data[116:116], io_mem_grant_bits_data[117:117], io_mem_grant_bits_data[118:118], io_mem_grant_bits_data[119:119], io_mem_grant_bits_data[120:120], io_mem_grant_bits_data[121:121], io_mem_grant_bits_data[122:122], io_mem_grant_bits_data[123:123], io_mem_grant_bits_data[124:124], io_mem_grant_bits_data[125:125], io_mem_grant_bits_data[126:126], io_mem_grant_bits_data[127:127] } : 1'b0;
  assign { N768, N766 } = (N46)? { 1'b1, 1'b1 } : 
                          (N67)? { N122, N123 } : 1'b0;
  assign { N1237, N1235, N1185, N1169, N1105, N1103, N1068, N1037, N973, N971, N951, N905, N841, N839, N779, N777, N775, N773, N771, N769 } = (N50)? { N766, N768, N702, N702, N634, N636, N570, N570, N502, N504, N438, N438, N370, N372, N306, N306, N306, N306, N306, N306 } : 
                                                                                                                                              (N51)? { N123, N122, 1'b0, 1'b0, N121, N120, 1'b0, 1'b0, N119, N118, 1'b0, 1'b0, N117, N116, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N50 = T137;
  assign N51 = N240;
  assign { N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1236, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1104, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N972, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N840, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N778, N776, N774, N772, N770 } = (N50)? { N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N767, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N635, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N503, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N371, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (N51)? { io_mem_grant_bits_data[127:64], io_mem_grant_bits_data[127:64], io_mem_grant_bits_data[127:64], io_mem_grant_bits_data[127:64], io_mem_grant_bits_data[127:64], io_mem_grant_bits_data[127:64], io_mem_grant_bits_data[127:64], io_mem_grant_bits_data[127:64] } : 1'b0;
  assign { N1379, N1377, N1375, N1373, N1371, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311 } = (N52)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1310)? { N770, N772, N774, N776, N778, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838 } : 1'b0;
  assign N52 = N1302;
  assign { N1380, N1378, N1376, N1374, N1372, N1370 } = (N52)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                        (N1310)? { N769, N771, N773, N775, N777, N779 } : 1'b0;
  assign { N1446, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382 } = (N53)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1381)? { N840, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904 } : 1'b0;
  assign N53 = N1303;
  assign { N1447, N1445 } = (N53)? { 1'b1, 1'b1 } : 
                            (N1381)? { N839, N841 } : 1'b0;
  assign { N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449 } = (N54)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1448)? { N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970 } : 1'b0;
  assign N54 = N1304;
  assign { N1514, N1468 } = (N54)? { 1'b1, 1'b1 } : 
                            (N1448)? { N905, N951 } : 1'b0;
  assign { N1580, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516 } = (N55)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1515)? { N972, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036 } : 1'b0;
  assign N55 = N1305;
  assign { N1581, N1579 } = (N55)? { 1'b1, 1'b1 } : 
                            (N1515)? { N971, N973 } : 1'b0;
  assign { N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583 } = (N56)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1582)? { N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102 } : 1'b0;
  assign N56 = N1306;
  assign { N1648, N1617 } = (N56)? { 1'b1, 1'b1 } : 
                            (N1582)? { N1037, N1068 } : 1'b0;
  assign { N1714, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650 } = (N57)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1649)? { N1104, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168 } : 1'b0;
  assign N57 = N1307;
  assign { N1715, N1713 } = (N57)? { 1'b1, 1'b1 } : 
                            (N1649)? { N1103, N1105 } : 1'b0;
  assign { N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717 } = (N58)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1716)? { N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234 } : 1'b0;
  assign N58 = N1308;
  assign { N1782, N1766 } = (N58)? { 1'b1, 1'b1 } : 
                            (N1716)? { N1169, N1185 } : 1'b0;
  assign { N1848, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784 } = (N59)? { rx_shifter_in_0, rx_shifter_in_1, rx_shifter_in_2, rx_shifter_in_3, T29[0:0], T29[1:1], T29[2:2], T29[3:3], T29[4:4], T29[5:5], T29[6:6], T29[7:7], T29[8:8], T29[9:9], T29[10:10], T29[11:11], rx_shifter_in[16:16], rx_shifter_in[17:17], rx_shifter_in[18:18], rx_shifter_in[19:19], rx_shifter_in[20:20], rx_shifter_in[21:21], rx_shifter_in[22:22], rx_shifter_in[23:23], rx_shifter_in[24:24], rx_shifter_in[25:25], rx_shifter_in[26:26], rx_shifter_in[27:27], rx_shifter_in[28:28], rx_shifter_in[29:29], rx_shifter_in[30:30], rx_shifter_in[31:31], rx_shifter_in[32:32], rx_shifter_in[33:33], rx_shifter_in[34:34], rx_shifter_in[35:35], rx_shifter_in[36:36], rx_shifter_in[37:37], rx_shifter_in[38:38], rx_shifter_in[39:39], rx_shifter_in[40:40], rx_shifter_in[41:41], rx_shifter_in[42:42], rx_shifter_in[43:43], rx_shifter_in[44:44], rx_shifter_in[45:45], rx_shifter_in[46:46], rx_shifter_in[47:47], io_host_in_bits[0:0], io_host_in_bits[1:1], io_host_in_bits[2:2], io_host_in_bits[3:3], io_host_in_bits[4:4], io_host_in_bits[5:5], io_host_in_bits[6:6], io_host_in_bits[7:7], io_host_in_bits[8:8], io_host_in_bits[9:9], io_host_in_bits[10:10], io_host_in_bits[11:11], io_host_in_bits[12:12], io_host_in_bits[13:13], io_host_in_bits[14:14], io_host_in_bits[15:15] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1783)? { N1236, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300 } : 1'b0;
  assign N59 = N1309;
  assign { N1849, N1847 } = (N59)? { 1'b1, 1'b1 } : 
                            (N1783)? { N1235, N1237 } : 1'b0;
  assign { N2318, N2316, N2266, N2250, N2186, N2184, N2149, N2118, N2054, N2052, N2032, N1986, N1922, N1920, N1860, N1858, N1856, N1854, N1852, N1850 } = (N60)? { N1847, N1849, N1766, N1782, N1713, N1715, N1617, N1648, N1579, N1581, N1468, N1514, N1445, N1447, N1370, N1372, N1374, N1376, N1378, N1380 } : 
                                                                                                                                                          (N61)? { N1237, N1235, N1185, N1169, N1105, N1103, N1068, N1037, N973, N971, N951, N905, N841, N839, N779, N777, N775, N773, N771, N769 } : 1'b0;
  assign N60 = T141;
  assign N61 = N1301;
  assign { N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2317, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2185, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2053, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1921, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1859, N1857, N1855, N1853, N1851 } = (N60)? { N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804, N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823, N1824, N1825, N1826, N1827, N1828, N1829, N1830, N1831, N1832, N1833, N1834, N1835, N1836, N1837, N1838, N1839, N1840, N1841, N1842, N1843, N1844, N1845, N1846, N1848, N1717, N1718, N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1765, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1650, N1651, N1652, N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1664, N1665, N1666, N1667, N1668, N1669, N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1714, N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616, N1618, N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578, N1580, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466, N1467, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1446, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1371, N1373, N1375, N1377, N1379 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N61)? { N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1236, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1104, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N972, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N840, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N778, N776, N774, N772, N770 } : 1'b0;
  assign N2384 = (N43)? 1'b1 : 
                 (N2500)? 1'b1 : 
                 (N2383)? 1'b0 : 1'b0;
  assign N2385 = (N43)? 1'b1 : 
                 (N2500)? io_scr_req_bits_data[0] : 1'b0;
  assign N2389 = (N62)? 1'b1 : 
                 (N2501)? 1'b1 : 
                 (N2503)? 1'b1 : 
                 (N2388)? 1'b0 : 1'b0;
  assign N62 = T132;
  assign { N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390 } = (N62)? io_scr_resp_bits : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2501)? io_cpu_0_csr_resp_bits : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2503)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, io_cpu_0_reset } : 1'b0;
  assign T2 = N2657 & io_mem_grant_valid;
  assign T16[0] = N2597;
  assign N63 = ~T18;
  assign T17[2] = N63;
  assign T18 = N2632 | N2636;
  assign T21 = T61 & N2617;
  assign T26 = T113 & T27;
  assign N64 = ~T32;
  assign T32 = T38 & T33;
  assign T33 = T35 | N2749;
  assign T35 = N2753 | N2757;
  assign T38 = ~nack;
  assign N65 = ~T54;
  assign N66 = ~T41;
  assign T41 = N2785 | N2789;
  assign bad_mem_packet = N2759 | N2761;
  assign T54 = N2777 | N2781;
  assign T60 = io_host_out_valid & io_host_out_ready;
  assign T61 = io_host_in_valid & io_host_in_ready;
  assign T66 = N2554 & rx_done;
  assign rx_done = rx_word_done & T67;
  assign T68 = T71 | N2651;
  assign T72 = N2644 & N2648;
  assign rx_word_done = io_host_in_valid & N2640;
  assign T79 = N2624 & cnt_done;
  assign cnt_done = T83 & N2679;
  assign T83 = T86 | T84;
  assign T84 = N2727 & io_mem_grant_valid;
  assign T86 = N2724 & io_mem_acquire_ready;
  assign T89 = N2639 & io_mem_acquire_ready;
  assign T91[2] = T92;
  assign T92 = N2584 | N2593;
  assign T101 = N2654 & io_mem_grant_valid;
  assign T103[2] = T104;
  assign T104 = N2570 | N2580;
  assign T107 = N2676 & cnt_done;
  assign T109[1] = T110;
  assign T110 = N2558 & N2566;
  assign T113 = N2678 & tx_done;
  assign tx_done = T120 & T114;
  assign T114 = T119 | T115;
  assign T115 = T118 & T116;
  assign T120 = io_host_out_ready & N2721;
  assign T123 = io_cpu_0_csr_req_ready & io_cpu_0_csr_req_valid;
  assign T124 = T126 & N2709;
  assign T126 = N2733 & N2738;
  assign T129 = N2730 & io_cpu_0_csr_resp_valid;
  assign T131 = io_scr_req_ready & io_scr_req_valid;
  assign T132 = N2741 & io_scr_resp_valid;
  assign T137 = N2660 & io_mem_grant_valid;
  assign T141 = rx_word_done & io_host_in_ready;
  assign io_scr_req_valid = N2744 & N2745;
  assign N67 = ~1'b0;
  assign N68 = ~T154[1];
  assign N69 = N67 & N68;
  assign N70 = N67 & T154[1];
  assign N71 = 1'b0 & N68;
  assign N72 = 1'b0 & T154[1];
  assign N73 = ~T154[2];
  assign N74 = N69 & N73;
  assign N75 = N69 & T154[2];
  assign N76 = N71 & N73;
  assign N77 = N71 & T154[2];
  assign N78 = N70 & N73;
  assign N79 = N70 & T154[2];
  assign N80 = N72 & N73;
  assign N81 = N72 & T154[2];
  assign N82 = ~1'b1;
  assign N83 = N82 & N68;
  assign N84 = N82 & T154[1];
  assign N85 = 1'b1 & N68;
  assign N86 = 1'b1 & T154[1];
  assign N87 = N83 & N73;
  assign N88 = N83 & T154[2];
  assign N89 = N85 & N73;
  assign N90 = N85 & T154[2];
  assign N91 = N84 & N73;
  assign N92 = N84 & T154[2];
  assign N93 = N86 & N73;
  assign N94 = N86 & T154[2];
  assign io_mem_acquire_bits_a_type[1] = N2526;
  assign io_mem_acquire_valid = N2518 | N2522;
  assign io_cpu_0_csr_req_valid = T185 & N2720;
  assign T185 = N2736 & N2738;
  assign T190 = T124 & N2621;
  assign N95 = ~T200;
  assign N96 = ~packet_ram_raddr[0];
  assign N97 = ~packet_ram_raddr[1];
  assign N98 = N96 & N97;
  assign N99 = N96 & packet_ram_raddr[1];
  assign N100 = packet_ram_raddr[0] & N97;
  assign N101 = packet_ram_raddr[0] & packet_ram_raddr[1];
  assign N102 = ~packet_ram_raddr[2];
  assign N103 = N98 & N102;
  assign N104 = N98 & packet_ram_raddr[2];
  assign N105 = N100 & N102;
  assign N106 = N100 & packet_ram_raddr[2];
  assign N107 = N99 & N102;
  assign N108 = N99 & packet_ram_raddr[2];
  assign N109 = N101 & N102;
  assign N110 = N101 & packet_ram_raddr[2];
  assign T200 = N2547 | N2551;
  assign tx_header_0 = nack;
  assign N111 = ~T2;
  assign N124 = T132 | reset;
  assign N125 = T131 | N124;
  assign N126 = T129 | N125;
  assign N127 = T124 | N126;
  assign N128 = T123 | N127;
  assign N129 = T113 | N128;
  assign N130 = T107 | N129;
  assign N131 = T101 | N130;
  assign N132 = T89 | N131;
  assign N133 = T79 | N132;
  assign N134 = T66 | N133;
  assign N135 = ~N134;
  assign N140 = T26 | reset;
  assign N141 = T61 | N140;
  assign N142 = ~N141;
  assign N159 = T101 | T107;
  assign N160 = T21 | N159;
  assign N161 = ~N160;
  assign N203 = T26 | reset;
  assign N204 = T60 | N203;
  assign N205 = ~N204;
  assign N222 = T83 | reset;
  assign N223 = ~N222;
  assign N227 = T101 | T107;
  assign N228 = T21 | N227;
  assign N229 = ~N228;
  assign N240 = ~T137;
  assign N241 = ~N306;
  assign N373 = ~N438;
  assign N505 = ~N570;
  assign N637 = ~N702;
  assign N1301 = ~T141;
  assign N1310 = ~N1302;
  assign N1381 = ~N1303;
  assign N1448 = ~N1304;
  assign N1515 = ~N1305;
  assign N1582 = ~N1306;
  assign N1649 = ~N1307;
  assign N1716 = ~N1308;
  assign N1783 = ~N1309;
  assign N2382 = T190 | reset;
  assign N2383 = ~N2382;
  assign N2386 = T129 | T132;
  assign N2387 = T124 | N2386;
  assign N2388 = ~N2387;
  assign N2454 = T132 & N2495;
  assign N2455 = ~T132;
  assign N2456 = N2495 & N2455;
  assign N2457 = T131 & N2456;
  assign N2458 = ~T131;
  assign N2459 = N2456 & N2458;
  assign N2460 = T129 & N2459;
  assign N2461 = ~T129;
  assign N2462 = N2459 & N2461;
  assign N2463 = T124 & N2462;
  assign N2464 = ~T124;
  assign N2465 = N2462 & N2464;
  assign N2466 = T123 & N2465;
  assign N2467 = ~T123;
  assign N2468 = N2465 & N2467;
  assign N2469 = T113 & N2468;
  assign N2470 = ~T113;
  assign N2471 = N2468 & N2470;
  assign N2472 = T107 & N2471;
  assign N2473 = ~T107;
  assign N2474 = N2471 & N2473;
  assign N2475 = T101 & N2474;
  assign N2476 = ~T101;
  assign N2477 = N2474 & N2476;
  assign N2478 = T89 & N2477;
  assign N2479 = ~T89;
  assign N2480 = N2477 & N2479;
  assign N2481 = T79 & N2480;
  assign N2482 = ~T79;
  assign N2483 = N2480 & N2482;
  assign N2484 = T66 & N2483;
  assign N2485 = T26 & N2495;
  assign N2486 = ~T26;
  assign N2487 = N2495 & N2486;
  assign N2488 = T61 & N2487;
  assign N2489 = T101 & N2473;
  assign N2490 = N2473 & N2476;
  assign N2491 = T21 & N2490;
  assign N2492 = T26 & N2495;
  assign N2493 = N2495 & N2486;
  assign N2494 = T60 & N2493;
  assign N2495 = ~reset;
  assign N2496 = T83 & N2495;
  assign N2497 = T101 & N2473;
  assign N2498 = N2473 & N2476;
  assign N2499 = T21 & N2498;
  assign N2500 = T190 & N2495;
  assign N2501 = T129 & N2455;
  assign N2502 = N2455 & N2461;
  assign N2503 = T124 & N2502;

endmodule