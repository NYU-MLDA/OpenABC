module bsg_mem_1r1w_synth_width_p73_els_p128_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [6:0] w_addr_i;
  input [72:0] w_data_i;
  input [6:0] r_addr_i;
  output [72:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [72:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566;
  reg [9343:0] mem;
  assign r_data_o[72] = (N145)? mem[72] : 
                        (N147)? mem[145] : 
                        (N149)? mem[218] : 
                        (N151)? mem[291] : 
                        (N153)? mem[364] : 
                        (N155)? mem[437] : 
                        (N157)? mem[510] : 
                        (N159)? mem[583] : 
                        (N161)? mem[656] : 
                        (N163)? mem[729] : 
                        (N165)? mem[802] : 
                        (N167)? mem[875] : 
                        (N169)? mem[948] : 
                        (N171)? mem[1021] : 
                        (N173)? mem[1094] : 
                        (N175)? mem[1167] : 
                        (N177)? mem[1240] : 
                        (N179)? mem[1313] : 
                        (N181)? mem[1386] : 
                        (N183)? mem[1459] : 
                        (N185)? mem[1532] : 
                        (N187)? mem[1605] : 
                        (N189)? mem[1678] : 
                        (N191)? mem[1751] : 
                        (N193)? mem[1824] : 
                        (N195)? mem[1897] : 
                        (N197)? mem[1970] : 
                        (N199)? mem[2043] : 
                        (N201)? mem[2116] : 
                        (N203)? mem[2189] : 
                        (N205)? mem[2262] : 
                        (N207)? mem[2335] : 
                        (N209)? mem[2408] : 
                        (N211)? mem[2481] : 
                        (N213)? mem[2554] : 
                        (N215)? mem[2627] : 
                        (N217)? mem[2700] : 
                        (N219)? mem[2773] : 
                        (N221)? mem[2846] : 
                        (N223)? mem[2919] : 
                        (N225)? mem[2992] : 
                        (N227)? mem[3065] : 
                        (N229)? mem[3138] : 
                        (N231)? mem[3211] : 
                        (N233)? mem[3284] : 
                        (N235)? mem[3357] : 
                        (N237)? mem[3430] : 
                        (N239)? mem[3503] : 
                        (N241)? mem[3576] : 
                        (N243)? mem[3649] : 
                        (N245)? mem[3722] : 
                        (N247)? mem[3795] : 
                        (N249)? mem[3868] : 
                        (N251)? mem[3941] : 
                        (N253)? mem[4014] : 
                        (N255)? mem[4087] : 
                        (N257)? mem[4160] : 
                        (N259)? mem[4233] : 
                        (N261)? mem[4306] : 
                        (N263)? mem[4379] : 
                        (N265)? mem[4452] : 
                        (N267)? mem[4525] : 
                        (N269)? mem[4598] : 
                        (N271)? mem[4671] : 
                        (N146)? mem[4744] : 
                        (N148)? mem[4817] : 
                        (N150)? mem[4890] : 
                        (N152)? mem[4963] : 
                        (N154)? mem[5036] : 
                        (N156)? mem[5109] : 
                        (N158)? mem[5182] : 
                        (N160)? mem[5255] : 
                        (N162)? mem[5328] : 
                        (N164)? mem[5401] : 
                        (N166)? mem[5474] : 
                        (N168)? mem[5547] : 
                        (N170)? mem[5620] : 
                        (N172)? mem[5693] : 
                        (N174)? mem[5766] : 
                        (N176)? mem[5839] : 
                        (N178)? mem[5912] : 
                        (N180)? mem[5985] : 
                        (N182)? mem[6058] : 
                        (N184)? mem[6131] : 
                        (N186)? mem[6204] : 
                        (N188)? mem[6277] : 
                        (N190)? mem[6350] : 
                        (N192)? mem[6423] : 
                        (N194)? mem[6496] : 
                        (N196)? mem[6569] : 
                        (N198)? mem[6642] : 
                        (N200)? mem[6715] : 
                        (N202)? mem[6788] : 
                        (N204)? mem[6861] : 
                        (N206)? mem[6934] : 
                        (N208)? mem[7007] : 
                        (N210)? mem[7080] : 
                        (N212)? mem[7153] : 
                        (N214)? mem[7226] : 
                        (N216)? mem[7299] : 
                        (N218)? mem[7372] : 
                        (N220)? mem[7445] : 
                        (N222)? mem[7518] : 
                        (N224)? mem[7591] : 
                        (N226)? mem[7664] : 
                        (N228)? mem[7737] : 
                        (N230)? mem[7810] : 
                        (N232)? mem[7883] : 
                        (N234)? mem[7956] : 
                        (N236)? mem[8029] : 
                        (N238)? mem[8102] : 
                        (N240)? mem[8175] : 
                        (N242)? mem[8248] : 
                        (N244)? mem[8321] : 
                        (N246)? mem[8394] : 
                        (N248)? mem[8467] : 
                        (N250)? mem[8540] : 
                        (N252)? mem[8613] : 
                        (N254)? mem[8686] : 
                        (N256)? mem[8759] : 
                        (N258)? mem[8832] : 
                        (N260)? mem[8905] : 
                        (N262)? mem[8978] : 
                        (N264)? mem[9051] : 
                        (N266)? mem[9124] : 
                        (N268)? mem[9197] : 
                        (N270)? mem[9270] : 
                        (N272)? mem[9343] : 1'b0;
  assign r_data_o[71] = (N145)? mem[71] : 
                        (N147)? mem[144] : 
                        (N149)? mem[217] : 
                        (N151)? mem[290] : 
                        (N153)? mem[363] : 
                        (N155)? mem[436] : 
                        (N157)? mem[509] : 
                        (N159)? mem[582] : 
                        (N161)? mem[655] : 
                        (N163)? mem[728] : 
                        (N165)? mem[801] : 
                        (N167)? mem[874] : 
                        (N169)? mem[947] : 
                        (N171)? mem[1020] : 
                        (N173)? mem[1093] : 
                        (N175)? mem[1166] : 
                        (N177)? mem[1239] : 
                        (N179)? mem[1312] : 
                        (N181)? mem[1385] : 
                        (N183)? mem[1458] : 
                        (N185)? mem[1531] : 
                        (N187)? mem[1604] : 
                        (N189)? mem[1677] : 
                        (N191)? mem[1750] : 
                        (N193)? mem[1823] : 
                        (N195)? mem[1896] : 
                        (N197)? mem[1969] : 
                        (N199)? mem[2042] : 
                        (N201)? mem[2115] : 
                        (N203)? mem[2188] : 
                        (N205)? mem[2261] : 
                        (N207)? mem[2334] : 
                        (N209)? mem[2407] : 
                        (N211)? mem[2480] : 
                        (N213)? mem[2553] : 
                        (N215)? mem[2626] : 
                        (N217)? mem[2699] : 
                        (N219)? mem[2772] : 
                        (N221)? mem[2845] : 
                        (N223)? mem[2918] : 
                        (N225)? mem[2991] : 
                        (N227)? mem[3064] : 
                        (N229)? mem[3137] : 
                        (N231)? mem[3210] : 
                        (N233)? mem[3283] : 
                        (N235)? mem[3356] : 
                        (N237)? mem[3429] : 
                        (N239)? mem[3502] : 
                        (N241)? mem[3575] : 
                        (N243)? mem[3648] : 
                        (N245)? mem[3721] : 
                        (N247)? mem[3794] : 
                        (N249)? mem[3867] : 
                        (N251)? mem[3940] : 
                        (N253)? mem[4013] : 
                        (N255)? mem[4086] : 
                        (N257)? mem[4159] : 
                        (N259)? mem[4232] : 
                        (N261)? mem[4305] : 
                        (N263)? mem[4378] : 
                        (N265)? mem[4451] : 
                        (N267)? mem[4524] : 
                        (N269)? mem[4597] : 
                        (N271)? mem[4670] : 
                        (N146)? mem[4743] : 
                        (N148)? mem[4816] : 
                        (N150)? mem[4889] : 
                        (N152)? mem[4962] : 
                        (N154)? mem[5035] : 
                        (N156)? mem[5108] : 
                        (N158)? mem[5181] : 
                        (N160)? mem[5254] : 
                        (N162)? mem[5327] : 
                        (N164)? mem[5400] : 
                        (N166)? mem[5473] : 
                        (N168)? mem[5546] : 
                        (N170)? mem[5619] : 
                        (N172)? mem[5692] : 
                        (N174)? mem[5765] : 
                        (N176)? mem[5838] : 
                        (N178)? mem[5911] : 
                        (N180)? mem[5984] : 
                        (N182)? mem[6057] : 
                        (N184)? mem[6130] : 
                        (N186)? mem[6203] : 
                        (N188)? mem[6276] : 
                        (N190)? mem[6349] : 
                        (N192)? mem[6422] : 
                        (N194)? mem[6495] : 
                        (N196)? mem[6568] : 
                        (N198)? mem[6641] : 
                        (N200)? mem[6714] : 
                        (N202)? mem[6787] : 
                        (N204)? mem[6860] : 
                        (N206)? mem[6933] : 
                        (N208)? mem[7006] : 
                        (N210)? mem[7079] : 
                        (N212)? mem[7152] : 
                        (N214)? mem[7225] : 
                        (N216)? mem[7298] : 
                        (N218)? mem[7371] : 
                        (N220)? mem[7444] : 
                        (N222)? mem[7517] : 
                        (N224)? mem[7590] : 
                        (N226)? mem[7663] : 
                        (N228)? mem[7736] : 
                        (N230)? mem[7809] : 
                        (N232)? mem[7882] : 
                        (N234)? mem[7955] : 
                        (N236)? mem[8028] : 
                        (N238)? mem[8101] : 
                        (N240)? mem[8174] : 
                        (N242)? mem[8247] : 
                        (N244)? mem[8320] : 
                        (N246)? mem[8393] : 
                        (N248)? mem[8466] : 
                        (N250)? mem[8539] : 
                        (N252)? mem[8612] : 
                        (N254)? mem[8685] : 
                        (N256)? mem[8758] : 
                        (N258)? mem[8831] : 
                        (N260)? mem[8904] : 
                        (N262)? mem[8977] : 
                        (N264)? mem[9050] : 
                        (N266)? mem[9123] : 
                        (N268)? mem[9196] : 
                        (N270)? mem[9269] : 
                        (N272)? mem[9342] : 1'b0;
  assign r_data_o[70] = (N145)? mem[70] : 
                        (N147)? mem[143] : 
                        (N149)? mem[216] : 
                        (N151)? mem[289] : 
                        (N153)? mem[362] : 
                        (N155)? mem[435] : 
                        (N157)? mem[508] : 
                        (N159)? mem[581] : 
                        (N161)? mem[654] : 
                        (N163)? mem[727] : 
                        (N165)? mem[800] : 
                        (N167)? mem[873] : 
                        (N169)? mem[946] : 
                        (N171)? mem[1019] : 
                        (N173)? mem[1092] : 
                        (N175)? mem[1165] : 
                        (N177)? mem[1238] : 
                        (N179)? mem[1311] : 
                        (N181)? mem[1384] : 
                        (N183)? mem[1457] : 
                        (N185)? mem[1530] : 
                        (N187)? mem[1603] : 
                        (N189)? mem[1676] : 
                        (N191)? mem[1749] : 
                        (N193)? mem[1822] : 
                        (N195)? mem[1895] : 
                        (N197)? mem[1968] : 
                        (N199)? mem[2041] : 
                        (N201)? mem[2114] : 
                        (N203)? mem[2187] : 
                        (N205)? mem[2260] : 
                        (N207)? mem[2333] : 
                        (N209)? mem[2406] : 
                        (N211)? mem[2479] : 
                        (N213)? mem[2552] : 
                        (N215)? mem[2625] : 
                        (N217)? mem[2698] : 
                        (N219)? mem[2771] : 
                        (N221)? mem[2844] : 
                        (N223)? mem[2917] : 
                        (N225)? mem[2990] : 
                        (N227)? mem[3063] : 
                        (N229)? mem[3136] : 
                        (N231)? mem[3209] : 
                        (N233)? mem[3282] : 
                        (N235)? mem[3355] : 
                        (N237)? mem[3428] : 
                        (N239)? mem[3501] : 
                        (N241)? mem[3574] : 
                        (N243)? mem[3647] : 
                        (N245)? mem[3720] : 
                        (N247)? mem[3793] : 
                        (N249)? mem[3866] : 
                        (N251)? mem[3939] : 
                        (N253)? mem[4012] : 
                        (N255)? mem[4085] : 
                        (N257)? mem[4158] : 
                        (N259)? mem[4231] : 
                        (N261)? mem[4304] : 
                        (N263)? mem[4377] : 
                        (N265)? mem[4450] : 
                        (N267)? mem[4523] : 
                        (N269)? mem[4596] : 
                        (N271)? mem[4669] : 
                        (N146)? mem[4742] : 
                        (N148)? mem[4815] : 
                        (N150)? mem[4888] : 
                        (N152)? mem[4961] : 
                        (N154)? mem[5034] : 
                        (N156)? mem[5107] : 
                        (N158)? mem[5180] : 
                        (N160)? mem[5253] : 
                        (N162)? mem[5326] : 
                        (N164)? mem[5399] : 
                        (N166)? mem[5472] : 
                        (N168)? mem[5545] : 
                        (N170)? mem[5618] : 
                        (N172)? mem[5691] : 
                        (N174)? mem[5764] : 
                        (N176)? mem[5837] : 
                        (N178)? mem[5910] : 
                        (N180)? mem[5983] : 
                        (N182)? mem[6056] : 
                        (N184)? mem[6129] : 
                        (N186)? mem[6202] : 
                        (N188)? mem[6275] : 
                        (N190)? mem[6348] : 
                        (N192)? mem[6421] : 
                        (N194)? mem[6494] : 
                        (N196)? mem[6567] : 
                        (N198)? mem[6640] : 
                        (N200)? mem[6713] : 
                        (N202)? mem[6786] : 
                        (N204)? mem[6859] : 
                        (N206)? mem[6932] : 
                        (N208)? mem[7005] : 
                        (N210)? mem[7078] : 
                        (N212)? mem[7151] : 
                        (N214)? mem[7224] : 
                        (N216)? mem[7297] : 
                        (N218)? mem[7370] : 
                        (N220)? mem[7443] : 
                        (N222)? mem[7516] : 
                        (N224)? mem[7589] : 
                        (N226)? mem[7662] : 
                        (N228)? mem[7735] : 
                        (N230)? mem[7808] : 
                        (N232)? mem[7881] : 
                        (N234)? mem[7954] : 
                        (N236)? mem[8027] : 
                        (N238)? mem[8100] : 
                        (N240)? mem[8173] : 
                        (N242)? mem[8246] : 
                        (N244)? mem[8319] : 
                        (N246)? mem[8392] : 
                        (N248)? mem[8465] : 
                        (N250)? mem[8538] : 
                        (N252)? mem[8611] : 
                        (N254)? mem[8684] : 
                        (N256)? mem[8757] : 
                        (N258)? mem[8830] : 
                        (N260)? mem[8903] : 
                        (N262)? mem[8976] : 
                        (N264)? mem[9049] : 
                        (N266)? mem[9122] : 
                        (N268)? mem[9195] : 
                        (N270)? mem[9268] : 
                        (N272)? mem[9341] : 1'b0;
  assign r_data_o[69] = (N145)? mem[69] : 
                        (N147)? mem[142] : 
                        (N149)? mem[215] : 
                        (N151)? mem[288] : 
                        (N153)? mem[361] : 
                        (N155)? mem[434] : 
                        (N157)? mem[507] : 
                        (N159)? mem[580] : 
                        (N161)? mem[653] : 
                        (N163)? mem[726] : 
                        (N165)? mem[799] : 
                        (N167)? mem[872] : 
                        (N169)? mem[945] : 
                        (N171)? mem[1018] : 
                        (N173)? mem[1091] : 
                        (N175)? mem[1164] : 
                        (N177)? mem[1237] : 
                        (N179)? mem[1310] : 
                        (N181)? mem[1383] : 
                        (N183)? mem[1456] : 
                        (N185)? mem[1529] : 
                        (N187)? mem[1602] : 
                        (N189)? mem[1675] : 
                        (N191)? mem[1748] : 
                        (N193)? mem[1821] : 
                        (N195)? mem[1894] : 
                        (N197)? mem[1967] : 
                        (N199)? mem[2040] : 
                        (N201)? mem[2113] : 
                        (N203)? mem[2186] : 
                        (N205)? mem[2259] : 
                        (N207)? mem[2332] : 
                        (N209)? mem[2405] : 
                        (N211)? mem[2478] : 
                        (N213)? mem[2551] : 
                        (N215)? mem[2624] : 
                        (N217)? mem[2697] : 
                        (N219)? mem[2770] : 
                        (N221)? mem[2843] : 
                        (N223)? mem[2916] : 
                        (N225)? mem[2989] : 
                        (N227)? mem[3062] : 
                        (N229)? mem[3135] : 
                        (N231)? mem[3208] : 
                        (N233)? mem[3281] : 
                        (N235)? mem[3354] : 
                        (N237)? mem[3427] : 
                        (N239)? mem[3500] : 
                        (N241)? mem[3573] : 
                        (N243)? mem[3646] : 
                        (N245)? mem[3719] : 
                        (N247)? mem[3792] : 
                        (N249)? mem[3865] : 
                        (N251)? mem[3938] : 
                        (N253)? mem[4011] : 
                        (N255)? mem[4084] : 
                        (N257)? mem[4157] : 
                        (N259)? mem[4230] : 
                        (N261)? mem[4303] : 
                        (N263)? mem[4376] : 
                        (N265)? mem[4449] : 
                        (N267)? mem[4522] : 
                        (N269)? mem[4595] : 
                        (N271)? mem[4668] : 
                        (N146)? mem[4741] : 
                        (N148)? mem[4814] : 
                        (N150)? mem[4887] : 
                        (N152)? mem[4960] : 
                        (N154)? mem[5033] : 
                        (N156)? mem[5106] : 
                        (N158)? mem[5179] : 
                        (N160)? mem[5252] : 
                        (N162)? mem[5325] : 
                        (N164)? mem[5398] : 
                        (N166)? mem[5471] : 
                        (N168)? mem[5544] : 
                        (N170)? mem[5617] : 
                        (N172)? mem[5690] : 
                        (N174)? mem[5763] : 
                        (N176)? mem[5836] : 
                        (N178)? mem[5909] : 
                        (N180)? mem[5982] : 
                        (N182)? mem[6055] : 
                        (N184)? mem[6128] : 
                        (N186)? mem[6201] : 
                        (N188)? mem[6274] : 
                        (N190)? mem[6347] : 
                        (N192)? mem[6420] : 
                        (N194)? mem[6493] : 
                        (N196)? mem[6566] : 
                        (N198)? mem[6639] : 
                        (N200)? mem[6712] : 
                        (N202)? mem[6785] : 
                        (N204)? mem[6858] : 
                        (N206)? mem[6931] : 
                        (N208)? mem[7004] : 
                        (N210)? mem[7077] : 
                        (N212)? mem[7150] : 
                        (N214)? mem[7223] : 
                        (N216)? mem[7296] : 
                        (N218)? mem[7369] : 
                        (N220)? mem[7442] : 
                        (N222)? mem[7515] : 
                        (N224)? mem[7588] : 
                        (N226)? mem[7661] : 
                        (N228)? mem[7734] : 
                        (N230)? mem[7807] : 
                        (N232)? mem[7880] : 
                        (N234)? mem[7953] : 
                        (N236)? mem[8026] : 
                        (N238)? mem[8099] : 
                        (N240)? mem[8172] : 
                        (N242)? mem[8245] : 
                        (N244)? mem[8318] : 
                        (N246)? mem[8391] : 
                        (N248)? mem[8464] : 
                        (N250)? mem[8537] : 
                        (N252)? mem[8610] : 
                        (N254)? mem[8683] : 
                        (N256)? mem[8756] : 
                        (N258)? mem[8829] : 
                        (N260)? mem[8902] : 
                        (N262)? mem[8975] : 
                        (N264)? mem[9048] : 
                        (N266)? mem[9121] : 
                        (N268)? mem[9194] : 
                        (N270)? mem[9267] : 
                        (N272)? mem[9340] : 1'b0;
  assign r_data_o[68] = (N145)? mem[68] : 
                        (N147)? mem[141] : 
                        (N149)? mem[214] : 
                        (N151)? mem[287] : 
                        (N153)? mem[360] : 
                        (N155)? mem[433] : 
                        (N157)? mem[506] : 
                        (N159)? mem[579] : 
                        (N161)? mem[652] : 
                        (N163)? mem[725] : 
                        (N165)? mem[798] : 
                        (N167)? mem[871] : 
                        (N169)? mem[944] : 
                        (N171)? mem[1017] : 
                        (N173)? mem[1090] : 
                        (N175)? mem[1163] : 
                        (N177)? mem[1236] : 
                        (N179)? mem[1309] : 
                        (N181)? mem[1382] : 
                        (N183)? mem[1455] : 
                        (N185)? mem[1528] : 
                        (N187)? mem[1601] : 
                        (N189)? mem[1674] : 
                        (N191)? mem[1747] : 
                        (N193)? mem[1820] : 
                        (N195)? mem[1893] : 
                        (N197)? mem[1966] : 
                        (N199)? mem[2039] : 
                        (N201)? mem[2112] : 
                        (N203)? mem[2185] : 
                        (N205)? mem[2258] : 
                        (N207)? mem[2331] : 
                        (N209)? mem[2404] : 
                        (N211)? mem[2477] : 
                        (N213)? mem[2550] : 
                        (N215)? mem[2623] : 
                        (N217)? mem[2696] : 
                        (N219)? mem[2769] : 
                        (N221)? mem[2842] : 
                        (N223)? mem[2915] : 
                        (N225)? mem[2988] : 
                        (N227)? mem[3061] : 
                        (N229)? mem[3134] : 
                        (N231)? mem[3207] : 
                        (N233)? mem[3280] : 
                        (N235)? mem[3353] : 
                        (N237)? mem[3426] : 
                        (N239)? mem[3499] : 
                        (N241)? mem[3572] : 
                        (N243)? mem[3645] : 
                        (N245)? mem[3718] : 
                        (N247)? mem[3791] : 
                        (N249)? mem[3864] : 
                        (N251)? mem[3937] : 
                        (N253)? mem[4010] : 
                        (N255)? mem[4083] : 
                        (N257)? mem[4156] : 
                        (N259)? mem[4229] : 
                        (N261)? mem[4302] : 
                        (N263)? mem[4375] : 
                        (N265)? mem[4448] : 
                        (N267)? mem[4521] : 
                        (N269)? mem[4594] : 
                        (N271)? mem[4667] : 
                        (N146)? mem[4740] : 
                        (N148)? mem[4813] : 
                        (N150)? mem[4886] : 
                        (N152)? mem[4959] : 
                        (N154)? mem[5032] : 
                        (N156)? mem[5105] : 
                        (N158)? mem[5178] : 
                        (N160)? mem[5251] : 
                        (N162)? mem[5324] : 
                        (N164)? mem[5397] : 
                        (N166)? mem[5470] : 
                        (N168)? mem[5543] : 
                        (N170)? mem[5616] : 
                        (N172)? mem[5689] : 
                        (N174)? mem[5762] : 
                        (N176)? mem[5835] : 
                        (N178)? mem[5908] : 
                        (N180)? mem[5981] : 
                        (N182)? mem[6054] : 
                        (N184)? mem[6127] : 
                        (N186)? mem[6200] : 
                        (N188)? mem[6273] : 
                        (N190)? mem[6346] : 
                        (N192)? mem[6419] : 
                        (N194)? mem[6492] : 
                        (N196)? mem[6565] : 
                        (N198)? mem[6638] : 
                        (N200)? mem[6711] : 
                        (N202)? mem[6784] : 
                        (N204)? mem[6857] : 
                        (N206)? mem[6930] : 
                        (N208)? mem[7003] : 
                        (N210)? mem[7076] : 
                        (N212)? mem[7149] : 
                        (N214)? mem[7222] : 
                        (N216)? mem[7295] : 
                        (N218)? mem[7368] : 
                        (N220)? mem[7441] : 
                        (N222)? mem[7514] : 
                        (N224)? mem[7587] : 
                        (N226)? mem[7660] : 
                        (N228)? mem[7733] : 
                        (N230)? mem[7806] : 
                        (N232)? mem[7879] : 
                        (N234)? mem[7952] : 
                        (N236)? mem[8025] : 
                        (N238)? mem[8098] : 
                        (N240)? mem[8171] : 
                        (N242)? mem[8244] : 
                        (N244)? mem[8317] : 
                        (N246)? mem[8390] : 
                        (N248)? mem[8463] : 
                        (N250)? mem[8536] : 
                        (N252)? mem[8609] : 
                        (N254)? mem[8682] : 
                        (N256)? mem[8755] : 
                        (N258)? mem[8828] : 
                        (N260)? mem[8901] : 
                        (N262)? mem[8974] : 
                        (N264)? mem[9047] : 
                        (N266)? mem[9120] : 
                        (N268)? mem[9193] : 
                        (N270)? mem[9266] : 
                        (N272)? mem[9339] : 1'b0;
  assign r_data_o[67] = (N145)? mem[67] : 
                        (N147)? mem[140] : 
                        (N149)? mem[213] : 
                        (N151)? mem[286] : 
                        (N153)? mem[359] : 
                        (N155)? mem[432] : 
                        (N157)? mem[505] : 
                        (N159)? mem[578] : 
                        (N161)? mem[651] : 
                        (N163)? mem[724] : 
                        (N165)? mem[797] : 
                        (N167)? mem[870] : 
                        (N169)? mem[943] : 
                        (N171)? mem[1016] : 
                        (N173)? mem[1089] : 
                        (N175)? mem[1162] : 
                        (N177)? mem[1235] : 
                        (N179)? mem[1308] : 
                        (N181)? mem[1381] : 
                        (N183)? mem[1454] : 
                        (N185)? mem[1527] : 
                        (N187)? mem[1600] : 
                        (N189)? mem[1673] : 
                        (N191)? mem[1746] : 
                        (N193)? mem[1819] : 
                        (N195)? mem[1892] : 
                        (N197)? mem[1965] : 
                        (N199)? mem[2038] : 
                        (N201)? mem[2111] : 
                        (N203)? mem[2184] : 
                        (N205)? mem[2257] : 
                        (N207)? mem[2330] : 
                        (N209)? mem[2403] : 
                        (N211)? mem[2476] : 
                        (N213)? mem[2549] : 
                        (N215)? mem[2622] : 
                        (N217)? mem[2695] : 
                        (N219)? mem[2768] : 
                        (N221)? mem[2841] : 
                        (N223)? mem[2914] : 
                        (N225)? mem[2987] : 
                        (N227)? mem[3060] : 
                        (N229)? mem[3133] : 
                        (N231)? mem[3206] : 
                        (N233)? mem[3279] : 
                        (N235)? mem[3352] : 
                        (N237)? mem[3425] : 
                        (N239)? mem[3498] : 
                        (N241)? mem[3571] : 
                        (N243)? mem[3644] : 
                        (N245)? mem[3717] : 
                        (N247)? mem[3790] : 
                        (N249)? mem[3863] : 
                        (N251)? mem[3936] : 
                        (N253)? mem[4009] : 
                        (N255)? mem[4082] : 
                        (N257)? mem[4155] : 
                        (N259)? mem[4228] : 
                        (N261)? mem[4301] : 
                        (N263)? mem[4374] : 
                        (N265)? mem[4447] : 
                        (N267)? mem[4520] : 
                        (N269)? mem[4593] : 
                        (N271)? mem[4666] : 
                        (N146)? mem[4739] : 
                        (N148)? mem[4812] : 
                        (N150)? mem[4885] : 
                        (N152)? mem[4958] : 
                        (N154)? mem[5031] : 
                        (N156)? mem[5104] : 
                        (N158)? mem[5177] : 
                        (N160)? mem[5250] : 
                        (N162)? mem[5323] : 
                        (N164)? mem[5396] : 
                        (N166)? mem[5469] : 
                        (N168)? mem[5542] : 
                        (N170)? mem[5615] : 
                        (N172)? mem[5688] : 
                        (N174)? mem[5761] : 
                        (N176)? mem[5834] : 
                        (N178)? mem[5907] : 
                        (N180)? mem[5980] : 
                        (N182)? mem[6053] : 
                        (N184)? mem[6126] : 
                        (N186)? mem[6199] : 
                        (N188)? mem[6272] : 
                        (N190)? mem[6345] : 
                        (N192)? mem[6418] : 
                        (N194)? mem[6491] : 
                        (N196)? mem[6564] : 
                        (N198)? mem[6637] : 
                        (N200)? mem[6710] : 
                        (N202)? mem[6783] : 
                        (N204)? mem[6856] : 
                        (N206)? mem[6929] : 
                        (N208)? mem[7002] : 
                        (N210)? mem[7075] : 
                        (N212)? mem[7148] : 
                        (N214)? mem[7221] : 
                        (N216)? mem[7294] : 
                        (N218)? mem[7367] : 
                        (N220)? mem[7440] : 
                        (N222)? mem[7513] : 
                        (N224)? mem[7586] : 
                        (N226)? mem[7659] : 
                        (N228)? mem[7732] : 
                        (N230)? mem[7805] : 
                        (N232)? mem[7878] : 
                        (N234)? mem[7951] : 
                        (N236)? mem[8024] : 
                        (N238)? mem[8097] : 
                        (N240)? mem[8170] : 
                        (N242)? mem[8243] : 
                        (N244)? mem[8316] : 
                        (N246)? mem[8389] : 
                        (N248)? mem[8462] : 
                        (N250)? mem[8535] : 
                        (N252)? mem[8608] : 
                        (N254)? mem[8681] : 
                        (N256)? mem[8754] : 
                        (N258)? mem[8827] : 
                        (N260)? mem[8900] : 
                        (N262)? mem[8973] : 
                        (N264)? mem[9046] : 
                        (N266)? mem[9119] : 
                        (N268)? mem[9192] : 
                        (N270)? mem[9265] : 
                        (N272)? mem[9338] : 1'b0;
  assign r_data_o[66] = (N145)? mem[66] : 
                        (N147)? mem[139] : 
                        (N149)? mem[212] : 
                        (N151)? mem[285] : 
                        (N153)? mem[358] : 
                        (N155)? mem[431] : 
                        (N157)? mem[504] : 
                        (N159)? mem[577] : 
                        (N161)? mem[650] : 
                        (N163)? mem[723] : 
                        (N165)? mem[796] : 
                        (N167)? mem[869] : 
                        (N169)? mem[942] : 
                        (N171)? mem[1015] : 
                        (N173)? mem[1088] : 
                        (N175)? mem[1161] : 
                        (N177)? mem[1234] : 
                        (N179)? mem[1307] : 
                        (N181)? mem[1380] : 
                        (N183)? mem[1453] : 
                        (N185)? mem[1526] : 
                        (N187)? mem[1599] : 
                        (N189)? mem[1672] : 
                        (N191)? mem[1745] : 
                        (N193)? mem[1818] : 
                        (N195)? mem[1891] : 
                        (N197)? mem[1964] : 
                        (N199)? mem[2037] : 
                        (N201)? mem[2110] : 
                        (N203)? mem[2183] : 
                        (N205)? mem[2256] : 
                        (N207)? mem[2329] : 
                        (N209)? mem[2402] : 
                        (N211)? mem[2475] : 
                        (N213)? mem[2548] : 
                        (N215)? mem[2621] : 
                        (N217)? mem[2694] : 
                        (N219)? mem[2767] : 
                        (N221)? mem[2840] : 
                        (N223)? mem[2913] : 
                        (N225)? mem[2986] : 
                        (N227)? mem[3059] : 
                        (N229)? mem[3132] : 
                        (N231)? mem[3205] : 
                        (N233)? mem[3278] : 
                        (N235)? mem[3351] : 
                        (N237)? mem[3424] : 
                        (N239)? mem[3497] : 
                        (N241)? mem[3570] : 
                        (N243)? mem[3643] : 
                        (N245)? mem[3716] : 
                        (N247)? mem[3789] : 
                        (N249)? mem[3862] : 
                        (N251)? mem[3935] : 
                        (N253)? mem[4008] : 
                        (N255)? mem[4081] : 
                        (N257)? mem[4154] : 
                        (N259)? mem[4227] : 
                        (N261)? mem[4300] : 
                        (N263)? mem[4373] : 
                        (N265)? mem[4446] : 
                        (N267)? mem[4519] : 
                        (N269)? mem[4592] : 
                        (N271)? mem[4665] : 
                        (N146)? mem[4738] : 
                        (N148)? mem[4811] : 
                        (N150)? mem[4884] : 
                        (N152)? mem[4957] : 
                        (N154)? mem[5030] : 
                        (N156)? mem[5103] : 
                        (N158)? mem[5176] : 
                        (N160)? mem[5249] : 
                        (N162)? mem[5322] : 
                        (N164)? mem[5395] : 
                        (N166)? mem[5468] : 
                        (N168)? mem[5541] : 
                        (N170)? mem[5614] : 
                        (N172)? mem[5687] : 
                        (N174)? mem[5760] : 
                        (N176)? mem[5833] : 
                        (N178)? mem[5906] : 
                        (N180)? mem[5979] : 
                        (N182)? mem[6052] : 
                        (N184)? mem[6125] : 
                        (N186)? mem[6198] : 
                        (N188)? mem[6271] : 
                        (N190)? mem[6344] : 
                        (N192)? mem[6417] : 
                        (N194)? mem[6490] : 
                        (N196)? mem[6563] : 
                        (N198)? mem[6636] : 
                        (N200)? mem[6709] : 
                        (N202)? mem[6782] : 
                        (N204)? mem[6855] : 
                        (N206)? mem[6928] : 
                        (N208)? mem[7001] : 
                        (N210)? mem[7074] : 
                        (N212)? mem[7147] : 
                        (N214)? mem[7220] : 
                        (N216)? mem[7293] : 
                        (N218)? mem[7366] : 
                        (N220)? mem[7439] : 
                        (N222)? mem[7512] : 
                        (N224)? mem[7585] : 
                        (N226)? mem[7658] : 
                        (N228)? mem[7731] : 
                        (N230)? mem[7804] : 
                        (N232)? mem[7877] : 
                        (N234)? mem[7950] : 
                        (N236)? mem[8023] : 
                        (N238)? mem[8096] : 
                        (N240)? mem[8169] : 
                        (N242)? mem[8242] : 
                        (N244)? mem[8315] : 
                        (N246)? mem[8388] : 
                        (N248)? mem[8461] : 
                        (N250)? mem[8534] : 
                        (N252)? mem[8607] : 
                        (N254)? mem[8680] : 
                        (N256)? mem[8753] : 
                        (N258)? mem[8826] : 
                        (N260)? mem[8899] : 
                        (N262)? mem[8972] : 
                        (N264)? mem[9045] : 
                        (N266)? mem[9118] : 
                        (N268)? mem[9191] : 
                        (N270)? mem[9264] : 
                        (N272)? mem[9337] : 1'b0;
  assign r_data_o[65] = (N145)? mem[65] : 
                        (N147)? mem[138] : 
                        (N149)? mem[211] : 
                        (N151)? mem[284] : 
                        (N153)? mem[357] : 
                        (N155)? mem[430] : 
                        (N157)? mem[503] : 
                        (N159)? mem[576] : 
                        (N161)? mem[649] : 
                        (N163)? mem[722] : 
                        (N165)? mem[795] : 
                        (N167)? mem[868] : 
                        (N169)? mem[941] : 
                        (N171)? mem[1014] : 
                        (N173)? mem[1087] : 
                        (N175)? mem[1160] : 
                        (N177)? mem[1233] : 
                        (N179)? mem[1306] : 
                        (N181)? mem[1379] : 
                        (N183)? mem[1452] : 
                        (N185)? mem[1525] : 
                        (N187)? mem[1598] : 
                        (N189)? mem[1671] : 
                        (N191)? mem[1744] : 
                        (N193)? mem[1817] : 
                        (N195)? mem[1890] : 
                        (N197)? mem[1963] : 
                        (N199)? mem[2036] : 
                        (N201)? mem[2109] : 
                        (N203)? mem[2182] : 
                        (N205)? mem[2255] : 
                        (N207)? mem[2328] : 
                        (N209)? mem[2401] : 
                        (N211)? mem[2474] : 
                        (N213)? mem[2547] : 
                        (N215)? mem[2620] : 
                        (N217)? mem[2693] : 
                        (N219)? mem[2766] : 
                        (N221)? mem[2839] : 
                        (N223)? mem[2912] : 
                        (N225)? mem[2985] : 
                        (N227)? mem[3058] : 
                        (N229)? mem[3131] : 
                        (N231)? mem[3204] : 
                        (N233)? mem[3277] : 
                        (N235)? mem[3350] : 
                        (N237)? mem[3423] : 
                        (N239)? mem[3496] : 
                        (N241)? mem[3569] : 
                        (N243)? mem[3642] : 
                        (N245)? mem[3715] : 
                        (N247)? mem[3788] : 
                        (N249)? mem[3861] : 
                        (N251)? mem[3934] : 
                        (N253)? mem[4007] : 
                        (N255)? mem[4080] : 
                        (N257)? mem[4153] : 
                        (N259)? mem[4226] : 
                        (N261)? mem[4299] : 
                        (N263)? mem[4372] : 
                        (N265)? mem[4445] : 
                        (N267)? mem[4518] : 
                        (N269)? mem[4591] : 
                        (N271)? mem[4664] : 
                        (N146)? mem[4737] : 
                        (N148)? mem[4810] : 
                        (N150)? mem[4883] : 
                        (N152)? mem[4956] : 
                        (N154)? mem[5029] : 
                        (N156)? mem[5102] : 
                        (N158)? mem[5175] : 
                        (N160)? mem[5248] : 
                        (N162)? mem[5321] : 
                        (N164)? mem[5394] : 
                        (N166)? mem[5467] : 
                        (N168)? mem[5540] : 
                        (N170)? mem[5613] : 
                        (N172)? mem[5686] : 
                        (N174)? mem[5759] : 
                        (N176)? mem[5832] : 
                        (N178)? mem[5905] : 
                        (N180)? mem[5978] : 
                        (N182)? mem[6051] : 
                        (N184)? mem[6124] : 
                        (N186)? mem[6197] : 
                        (N188)? mem[6270] : 
                        (N190)? mem[6343] : 
                        (N192)? mem[6416] : 
                        (N194)? mem[6489] : 
                        (N196)? mem[6562] : 
                        (N198)? mem[6635] : 
                        (N200)? mem[6708] : 
                        (N202)? mem[6781] : 
                        (N204)? mem[6854] : 
                        (N206)? mem[6927] : 
                        (N208)? mem[7000] : 
                        (N210)? mem[7073] : 
                        (N212)? mem[7146] : 
                        (N214)? mem[7219] : 
                        (N216)? mem[7292] : 
                        (N218)? mem[7365] : 
                        (N220)? mem[7438] : 
                        (N222)? mem[7511] : 
                        (N224)? mem[7584] : 
                        (N226)? mem[7657] : 
                        (N228)? mem[7730] : 
                        (N230)? mem[7803] : 
                        (N232)? mem[7876] : 
                        (N234)? mem[7949] : 
                        (N236)? mem[8022] : 
                        (N238)? mem[8095] : 
                        (N240)? mem[8168] : 
                        (N242)? mem[8241] : 
                        (N244)? mem[8314] : 
                        (N246)? mem[8387] : 
                        (N248)? mem[8460] : 
                        (N250)? mem[8533] : 
                        (N252)? mem[8606] : 
                        (N254)? mem[8679] : 
                        (N256)? mem[8752] : 
                        (N258)? mem[8825] : 
                        (N260)? mem[8898] : 
                        (N262)? mem[8971] : 
                        (N264)? mem[9044] : 
                        (N266)? mem[9117] : 
                        (N268)? mem[9190] : 
                        (N270)? mem[9263] : 
                        (N272)? mem[9336] : 1'b0;
  assign r_data_o[64] = (N145)? mem[64] : 
                        (N147)? mem[137] : 
                        (N149)? mem[210] : 
                        (N151)? mem[283] : 
                        (N153)? mem[356] : 
                        (N155)? mem[429] : 
                        (N157)? mem[502] : 
                        (N159)? mem[575] : 
                        (N161)? mem[648] : 
                        (N163)? mem[721] : 
                        (N165)? mem[794] : 
                        (N167)? mem[867] : 
                        (N169)? mem[940] : 
                        (N171)? mem[1013] : 
                        (N173)? mem[1086] : 
                        (N175)? mem[1159] : 
                        (N177)? mem[1232] : 
                        (N179)? mem[1305] : 
                        (N181)? mem[1378] : 
                        (N183)? mem[1451] : 
                        (N185)? mem[1524] : 
                        (N187)? mem[1597] : 
                        (N189)? mem[1670] : 
                        (N191)? mem[1743] : 
                        (N193)? mem[1816] : 
                        (N195)? mem[1889] : 
                        (N197)? mem[1962] : 
                        (N199)? mem[2035] : 
                        (N201)? mem[2108] : 
                        (N203)? mem[2181] : 
                        (N205)? mem[2254] : 
                        (N207)? mem[2327] : 
                        (N209)? mem[2400] : 
                        (N211)? mem[2473] : 
                        (N213)? mem[2546] : 
                        (N215)? mem[2619] : 
                        (N217)? mem[2692] : 
                        (N219)? mem[2765] : 
                        (N221)? mem[2838] : 
                        (N223)? mem[2911] : 
                        (N225)? mem[2984] : 
                        (N227)? mem[3057] : 
                        (N229)? mem[3130] : 
                        (N231)? mem[3203] : 
                        (N233)? mem[3276] : 
                        (N235)? mem[3349] : 
                        (N237)? mem[3422] : 
                        (N239)? mem[3495] : 
                        (N241)? mem[3568] : 
                        (N243)? mem[3641] : 
                        (N245)? mem[3714] : 
                        (N247)? mem[3787] : 
                        (N249)? mem[3860] : 
                        (N251)? mem[3933] : 
                        (N253)? mem[4006] : 
                        (N255)? mem[4079] : 
                        (N257)? mem[4152] : 
                        (N259)? mem[4225] : 
                        (N261)? mem[4298] : 
                        (N263)? mem[4371] : 
                        (N265)? mem[4444] : 
                        (N267)? mem[4517] : 
                        (N269)? mem[4590] : 
                        (N271)? mem[4663] : 
                        (N146)? mem[4736] : 
                        (N148)? mem[4809] : 
                        (N150)? mem[4882] : 
                        (N152)? mem[4955] : 
                        (N154)? mem[5028] : 
                        (N156)? mem[5101] : 
                        (N158)? mem[5174] : 
                        (N160)? mem[5247] : 
                        (N162)? mem[5320] : 
                        (N164)? mem[5393] : 
                        (N166)? mem[5466] : 
                        (N168)? mem[5539] : 
                        (N170)? mem[5612] : 
                        (N172)? mem[5685] : 
                        (N174)? mem[5758] : 
                        (N176)? mem[5831] : 
                        (N178)? mem[5904] : 
                        (N180)? mem[5977] : 
                        (N182)? mem[6050] : 
                        (N184)? mem[6123] : 
                        (N186)? mem[6196] : 
                        (N188)? mem[6269] : 
                        (N190)? mem[6342] : 
                        (N192)? mem[6415] : 
                        (N194)? mem[6488] : 
                        (N196)? mem[6561] : 
                        (N198)? mem[6634] : 
                        (N200)? mem[6707] : 
                        (N202)? mem[6780] : 
                        (N204)? mem[6853] : 
                        (N206)? mem[6926] : 
                        (N208)? mem[6999] : 
                        (N210)? mem[7072] : 
                        (N212)? mem[7145] : 
                        (N214)? mem[7218] : 
                        (N216)? mem[7291] : 
                        (N218)? mem[7364] : 
                        (N220)? mem[7437] : 
                        (N222)? mem[7510] : 
                        (N224)? mem[7583] : 
                        (N226)? mem[7656] : 
                        (N228)? mem[7729] : 
                        (N230)? mem[7802] : 
                        (N232)? mem[7875] : 
                        (N234)? mem[7948] : 
                        (N236)? mem[8021] : 
                        (N238)? mem[8094] : 
                        (N240)? mem[8167] : 
                        (N242)? mem[8240] : 
                        (N244)? mem[8313] : 
                        (N246)? mem[8386] : 
                        (N248)? mem[8459] : 
                        (N250)? mem[8532] : 
                        (N252)? mem[8605] : 
                        (N254)? mem[8678] : 
                        (N256)? mem[8751] : 
                        (N258)? mem[8824] : 
                        (N260)? mem[8897] : 
                        (N262)? mem[8970] : 
                        (N264)? mem[9043] : 
                        (N266)? mem[9116] : 
                        (N268)? mem[9189] : 
                        (N270)? mem[9262] : 
                        (N272)? mem[9335] : 1'b0;
  assign r_data_o[63] = (N145)? mem[63] : 
                        (N147)? mem[136] : 
                        (N149)? mem[209] : 
                        (N151)? mem[282] : 
                        (N153)? mem[355] : 
                        (N155)? mem[428] : 
                        (N157)? mem[501] : 
                        (N159)? mem[574] : 
                        (N161)? mem[647] : 
                        (N163)? mem[720] : 
                        (N165)? mem[793] : 
                        (N167)? mem[866] : 
                        (N169)? mem[939] : 
                        (N171)? mem[1012] : 
                        (N173)? mem[1085] : 
                        (N175)? mem[1158] : 
                        (N177)? mem[1231] : 
                        (N179)? mem[1304] : 
                        (N181)? mem[1377] : 
                        (N183)? mem[1450] : 
                        (N185)? mem[1523] : 
                        (N187)? mem[1596] : 
                        (N189)? mem[1669] : 
                        (N191)? mem[1742] : 
                        (N193)? mem[1815] : 
                        (N195)? mem[1888] : 
                        (N197)? mem[1961] : 
                        (N199)? mem[2034] : 
                        (N201)? mem[2107] : 
                        (N203)? mem[2180] : 
                        (N205)? mem[2253] : 
                        (N207)? mem[2326] : 
                        (N209)? mem[2399] : 
                        (N211)? mem[2472] : 
                        (N213)? mem[2545] : 
                        (N215)? mem[2618] : 
                        (N217)? mem[2691] : 
                        (N219)? mem[2764] : 
                        (N221)? mem[2837] : 
                        (N223)? mem[2910] : 
                        (N225)? mem[2983] : 
                        (N227)? mem[3056] : 
                        (N229)? mem[3129] : 
                        (N231)? mem[3202] : 
                        (N233)? mem[3275] : 
                        (N235)? mem[3348] : 
                        (N237)? mem[3421] : 
                        (N239)? mem[3494] : 
                        (N241)? mem[3567] : 
                        (N243)? mem[3640] : 
                        (N245)? mem[3713] : 
                        (N247)? mem[3786] : 
                        (N249)? mem[3859] : 
                        (N251)? mem[3932] : 
                        (N253)? mem[4005] : 
                        (N255)? mem[4078] : 
                        (N257)? mem[4151] : 
                        (N259)? mem[4224] : 
                        (N261)? mem[4297] : 
                        (N263)? mem[4370] : 
                        (N265)? mem[4443] : 
                        (N267)? mem[4516] : 
                        (N269)? mem[4589] : 
                        (N271)? mem[4662] : 
                        (N146)? mem[4735] : 
                        (N148)? mem[4808] : 
                        (N150)? mem[4881] : 
                        (N152)? mem[4954] : 
                        (N154)? mem[5027] : 
                        (N156)? mem[5100] : 
                        (N158)? mem[5173] : 
                        (N160)? mem[5246] : 
                        (N162)? mem[5319] : 
                        (N164)? mem[5392] : 
                        (N166)? mem[5465] : 
                        (N168)? mem[5538] : 
                        (N170)? mem[5611] : 
                        (N172)? mem[5684] : 
                        (N174)? mem[5757] : 
                        (N176)? mem[5830] : 
                        (N178)? mem[5903] : 
                        (N180)? mem[5976] : 
                        (N182)? mem[6049] : 
                        (N184)? mem[6122] : 
                        (N186)? mem[6195] : 
                        (N188)? mem[6268] : 
                        (N190)? mem[6341] : 
                        (N192)? mem[6414] : 
                        (N194)? mem[6487] : 
                        (N196)? mem[6560] : 
                        (N198)? mem[6633] : 
                        (N200)? mem[6706] : 
                        (N202)? mem[6779] : 
                        (N204)? mem[6852] : 
                        (N206)? mem[6925] : 
                        (N208)? mem[6998] : 
                        (N210)? mem[7071] : 
                        (N212)? mem[7144] : 
                        (N214)? mem[7217] : 
                        (N216)? mem[7290] : 
                        (N218)? mem[7363] : 
                        (N220)? mem[7436] : 
                        (N222)? mem[7509] : 
                        (N224)? mem[7582] : 
                        (N226)? mem[7655] : 
                        (N228)? mem[7728] : 
                        (N230)? mem[7801] : 
                        (N232)? mem[7874] : 
                        (N234)? mem[7947] : 
                        (N236)? mem[8020] : 
                        (N238)? mem[8093] : 
                        (N240)? mem[8166] : 
                        (N242)? mem[8239] : 
                        (N244)? mem[8312] : 
                        (N246)? mem[8385] : 
                        (N248)? mem[8458] : 
                        (N250)? mem[8531] : 
                        (N252)? mem[8604] : 
                        (N254)? mem[8677] : 
                        (N256)? mem[8750] : 
                        (N258)? mem[8823] : 
                        (N260)? mem[8896] : 
                        (N262)? mem[8969] : 
                        (N264)? mem[9042] : 
                        (N266)? mem[9115] : 
                        (N268)? mem[9188] : 
                        (N270)? mem[9261] : 
                        (N272)? mem[9334] : 1'b0;
  assign r_data_o[62] = (N145)? mem[62] : 
                        (N147)? mem[135] : 
                        (N149)? mem[208] : 
                        (N151)? mem[281] : 
                        (N153)? mem[354] : 
                        (N155)? mem[427] : 
                        (N157)? mem[500] : 
                        (N159)? mem[573] : 
                        (N161)? mem[646] : 
                        (N163)? mem[719] : 
                        (N165)? mem[792] : 
                        (N167)? mem[865] : 
                        (N169)? mem[938] : 
                        (N171)? mem[1011] : 
                        (N173)? mem[1084] : 
                        (N175)? mem[1157] : 
                        (N177)? mem[1230] : 
                        (N179)? mem[1303] : 
                        (N181)? mem[1376] : 
                        (N183)? mem[1449] : 
                        (N185)? mem[1522] : 
                        (N187)? mem[1595] : 
                        (N189)? mem[1668] : 
                        (N191)? mem[1741] : 
                        (N193)? mem[1814] : 
                        (N195)? mem[1887] : 
                        (N197)? mem[1960] : 
                        (N199)? mem[2033] : 
                        (N201)? mem[2106] : 
                        (N203)? mem[2179] : 
                        (N205)? mem[2252] : 
                        (N207)? mem[2325] : 
                        (N209)? mem[2398] : 
                        (N211)? mem[2471] : 
                        (N213)? mem[2544] : 
                        (N215)? mem[2617] : 
                        (N217)? mem[2690] : 
                        (N219)? mem[2763] : 
                        (N221)? mem[2836] : 
                        (N223)? mem[2909] : 
                        (N225)? mem[2982] : 
                        (N227)? mem[3055] : 
                        (N229)? mem[3128] : 
                        (N231)? mem[3201] : 
                        (N233)? mem[3274] : 
                        (N235)? mem[3347] : 
                        (N237)? mem[3420] : 
                        (N239)? mem[3493] : 
                        (N241)? mem[3566] : 
                        (N243)? mem[3639] : 
                        (N245)? mem[3712] : 
                        (N247)? mem[3785] : 
                        (N249)? mem[3858] : 
                        (N251)? mem[3931] : 
                        (N253)? mem[4004] : 
                        (N255)? mem[4077] : 
                        (N257)? mem[4150] : 
                        (N259)? mem[4223] : 
                        (N261)? mem[4296] : 
                        (N263)? mem[4369] : 
                        (N265)? mem[4442] : 
                        (N267)? mem[4515] : 
                        (N269)? mem[4588] : 
                        (N271)? mem[4661] : 
                        (N146)? mem[4734] : 
                        (N148)? mem[4807] : 
                        (N150)? mem[4880] : 
                        (N152)? mem[4953] : 
                        (N154)? mem[5026] : 
                        (N156)? mem[5099] : 
                        (N158)? mem[5172] : 
                        (N160)? mem[5245] : 
                        (N162)? mem[5318] : 
                        (N164)? mem[5391] : 
                        (N166)? mem[5464] : 
                        (N168)? mem[5537] : 
                        (N170)? mem[5610] : 
                        (N172)? mem[5683] : 
                        (N174)? mem[5756] : 
                        (N176)? mem[5829] : 
                        (N178)? mem[5902] : 
                        (N180)? mem[5975] : 
                        (N182)? mem[6048] : 
                        (N184)? mem[6121] : 
                        (N186)? mem[6194] : 
                        (N188)? mem[6267] : 
                        (N190)? mem[6340] : 
                        (N192)? mem[6413] : 
                        (N194)? mem[6486] : 
                        (N196)? mem[6559] : 
                        (N198)? mem[6632] : 
                        (N200)? mem[6705] : 
                        (N202)? mem[6778] : 
                        (N204)? mem[6851] : 
                        (N206)? mem[6924] : 
                        (N208)? mem[6997] : 
                        (N210)? mem[7070] : 
                        (N212)? mem[7143] : 
                        (N214)? mem[7216] : 
                        (N216)? mem[7289] : 
                        (N218)? mem[7362] : 
                        (N220)? mem[7435] : 
                        (N222)? mem[7508] : 
                        (N224)? mem[7581] : 
                        (N226)? mem[7654] : 
                        (N228)? mem[7727] : 
                        (N230)? mem[7800] : 
                        (N232)? mem[7873] : 
                        (N234)? mem[7946] : 
                        (N236)? mem[8019] : 
                        (N238)? mem[8092] : 
                        (N240)? mem[8165] : 
                        (N242)? mem[8238] : 
                        (N244)? mem[8311] : 
                        (N246)? mem[8384] : 
                        (N248)? mem[8457] : 
                        (N250)? mem[8530] : 
                        (N252)? mem[8603] : 
                        (N254)? mem[8676] : 
                        (N256)? mem[8749] : 
                        (N258)? mem[8822] : 
                        (N260)? mem[8895] : 
                        (N262)? mem[8968] : 
                        (N264)? mem[9041] : 
                        (N266)? mem[9114] : 
                        (N268)? mem[9187] : 
                        (N270)? mem[9260] : 
                        (N272)? mem[9333] : 1'b0;
  assign r_data_o[61] = (N145)? mem[61] : 
                        (N147)? mem[134] : 
                        (N149)? mem[207] : 
                        (N151)? mem[280] : 
                        (N153)? mem[353] : 
                        (N155)? mem[426] : 
                        (N157)? mem[499] : 
                        (N159)? mem[572] : 
                        (N161)? mem[645] : 
                        (N163)? mem[718] : 
                        (N165)? mem[791] : 
                        (N167)? mem[864] : 
                        (N169)? mem[937] : 
                        (N171)? mem[1010] : 
                        (N173)? mem[1083] : 
                        (N175)? mem[1156] : 
                        (N177)? mem[1229] : 
                        (N179)? mem[1302] : 
                        (N181)? mem[1375] : 
                        (N183)? mem[1448] : 
                        (N185)? mem[1521] : 
                        (N187)? mem[1594] : 
                        (N189)? mem[1667] : 
                        (N191)? mem[1740] : 
                        (N193)? mem[1813] : 
                        (N195)? mem[1886] : 
                        (N197)? mem[1959] : 
                        (N199)? mem[2032] : 
                        (N201)? mem[2105] : 
                        (N203)? mem[2178] : 
                        (N205)? mem[2251] : 
                        (N207)? mem[2324] : 
                        (N209)? mem[2397] : 
                        (N211)? mem[2470] : 
                        (N213)? mem[2543] : 
                        (N215)? mem[2616] : 
                        (N217)? mem[2689] : 
                        (N219)? mem[2762] : 
                        (N221)? mem[2835] : 
                        (N223)? mem[2908] : 
                        (N225)? mem[2981] : 
                        (N227)? mem[3054] : 
                        (N229)? mem[3127] : 
                        (N231)? mem[3200] : 
                        (N233)? mem[3273] : 
                        (N235)? mem[3346] : 
                        (N237)? mem[3419] : 
                        (N239)? mem[3492] : 
                        (N241)? mem[3565] : 
                        (N243)? mem[3638] : 
                        (N245)? mem[3711] : 
                        (N247)? mem[3784] : 
                        (N249)? mem[3857] : 
                        (N251)? mem[3930] : 
                        (N253)? mem[4003] : 
                        (N255)? mem[4076] : 
                        (N257)? mem[4149] : 
                        (N259)? mem[4222] : 
                        (N261)? mem[4295] : 
                        (N263)? mem[4368] : 
                        (N265)? mem[4441] : 
                        (N267)? mem[4514] : 
                        (N269)? mem[4587] : 
                        (N271)? mem[4660] : 
                        (N146)? mem[4733] : 
                        (N148)? mem[4806] : 
                        (N150)? mem[4879] : 
                        (N152)? mem[4952] : 
                        (N154)? mem[5025] : 
                        (N156)? mem[5098] : 
                        (N158)? mem[5171] : 
                        (N160)? mem[5244] : 
                        (N162)? mem[5317] : 
                        (N164)? mem[5390] : 
                        (N166)? mem[5463] : 
                        (N168)? mem[5536] : 
                        (N170)? mem[5609] : 
                        (N172)? mem[5682] : 
                        (N174)? mem[5755] : 
                        (N176)? mem[5828] : 
                        (N178)? mem[5901] : 
                        (N180)? mem[5974] : 
                        (N182)? mem[6047] : 
                        (N184)? mem[6120] : 
                        (N186)? mem[6193] : 
                        (N188)? mem[6266] : 
                        (N190)? mem[6339] : 
                        (N192)? mem[6412] : 
                        (N194)? mem[6485] : 
                        (N196)? mem[6558] : 
                        (N198)? mem[6631] : 
                        (N200)? mem[6704] : 
                        (N202)? mem[6777] : 
                        (N204)? mem[6850] : 
                        (N206)? mem[6923] : 
                        (N208)? mem[6996] : 
                        (N210)? mem[7069] : 
                        (N212)? mem[7142] : 
                        (N214)? mem[7215] : 
                        (N216)? mem[7288] : 
                        (N218)? mem[7361] : 
                        (N220)? mem[7434] : 
                        (N222)? mem[7507] : 
                        (N224)? mem[7580] : 
                        (N226)? mem[7653] : 
                        (N228)? mem[7726] : 
                        (N230)? mem[7799] : 
                        (N232)? mem[7872] : 
                        (N234)? mem[7945] : 
                        (N236)? mem[8018] : 
                        (N238)? mem[8091] : 
                        (N240)? mem[8164] : 
                        (N242)? mem[8237] : 
                        (N244)? mem[8310] : 
                        (N246)? mem[8383] : 
                        (N248)? mem[8456] : 
                        (N250)? mem[8529] : 
                        (N252)? mem[8602] : 
                        (N254)? mem[8675] : 
                        (N256)? mem[8748] : 
                        (N258)? mem[8821] : 
                        (N260)? mem[8894] : 
                        (N262)? mem[8967] : 
                        (N264)? mem[9040] : 
                        (N266)? mem[9113] : 
                        (N268)? mem[9186] : 
                        (N270)? mem[9259] : 
                        (N272)? mem[9332] : 1'b0;
  assign r_data_o[60] = (N145)? mem[60] : 
                        (N147)? mem[133] : 
                        (N149)? mem[206] : 
                        (N151)? mem[279] : 
                        (N153)? mem[352] : 
                        (N155)? mem[425] : 
                        (N157)? mem[498] : 
                        (N159)? mem[571] : 
                        (N161)? mem[644] : 
                        (N163)? mem[717] : 
                        (N165)? mem[790] : 
                        (N167)? mem[863] : 
                        (N169)? mem[936] : 
                        (N171)? mem[1009] : 
                        (N173)? mem[1082] : 
                        (N175)? mem[1155] : 
                        (N177)? mem[1228] : 
                        (N179)? mem[1301] : 
                        (N181)? mem[1374] : 
                        (N183)? mem[1447] : 
                        (N185)? mem[1520] : 
                        (N187)? mem[1593] : 
                        (N189)? mem[1666] : 
                        (N191)? mem[1739] : 
                        (N193)? mem[1812] : 
                        (N195)? mem[1885] : 
                        (N197)? mem[1958] : 
                        (N199)? mem[2031] : 
                        (N201)? mem[2104] : 
                        (N203)? mem[2177] : 
                        (N205)? mem[2250] : 
                        (N207)? mem[2323] : 
                        (N209)? mem[2396] : 
                        (N211)? mem[2469] : 
                        (N213)? mem[2542] : 
                        (N215)? mem[2615] : 
                        (N217)? mem[2688] : 
                        (N219)? mem[2761] : 
                        (N221)? mem[2834] : 
                        (N223)? mem[2907] : 
                        (N225)? mem[2980] : 
                        (N227)? mem[3053] : 
                        (N229)? mem[3126] : 
                        (N231)? mem[3199] : 
                        (N233)? mem[3272] : 
                        (N235)? mem[3345] : 
                        (N237)? mem[3418] : 
                        (N239)? mem[3491] : 
                        (N241)? mem[3564] : 
                        (N243)? mem[3637] : 
                        (N245)? mem[3710] : 
                        (N247)? mem[3783] : 
                        (N249)? mem[3856] : 
                        (N251)? mem[3929] : 
                        (N253)? mem[4002] : 
                        (N255)? mem[4075] : 
                        (N257)? mem[4148] : 
                        (N259)? mem[4221] : 
                        (N261)? mem[4294] : 
                        (N263)? mem[4367] : 
                        (N265)? mem[4440] : 
                        (N267)? mem[4513] : 
                        (N269)? mem[4586] : 
                        (N271)? mem[4659] : 
                        (N146)? mem[4732] : 
                        (N148)? mem[4805] : 
                        (N150)? mem[4878] : 
                        (N152)? mem[4951] : 
                        (N154)? mem[5024] : 
                        (N156)? mem[5097] : 
                        (N158)? mem[5170] : 
                        (N160)? mem[5243] : 
                        (N162)? mem[5316] : 
                        (N164)? mem[5389] : 
                        (N166)? mem[5462] : 
                        (N168)? mem[5535] : 
                        (N170)? mem[5608] : 
                        (N172)? mem[5681] : 
                        (N174)? mem[5754] : 
                        (N176)? mem[5827] : 
                        (N178)? mem[5900] : 
                        (N180)? mem[5973] : 
                        (N182)? mem[6046] : 
                        (N184)? mem[6119] : 
                        (N186)? mem[6192] : 
                        (N188)? mem[6265] : 
                        (N190)? mem[6338] : 
                        (N192)? mem[6411] : 
                        (N194)? mem[6484] : 
                        (N196)? mem[6557] : 
                        (N198)? mem[6630] : 
                        (N200)? mem[6703] : 
                        (N202)? mem[6776] : 
                        (N204)? mem[6849] : 
                        (N206)? mem[6922] : 
                        (N208)? mem[6995] : 
                        (N210)? mem[7068] : 
                        (N212)? mem[7141] : 
                        (N214)? mem[7214] : 
                        (N216)? mem[7287] : 
                        (N218)? mem[7360] : 
                        (N220)? mem[7433] : 
                        (N222)? mem[7506] : 
                        (N224)? mem[7579] : 
                        (N226)? mem[7652] : 
                        (N228)? mem[7725] : 
                        (N230)? mem[7798] : 
                        (N232)? mem[7871] : 
                        (N234)? mem[7944] : 
                        (N236)? mem[8017] : 
                        (N238)? mem[8090] : 
                        (N240)? mem[8163] : 
                        (N242)? mem[8236] : 
                        (N244)? mem[8309] : 
                        (N246)? mem[8382] : 
                        (N248)? mem[8455] : 
                        (N250)? mem[8528] : 
                        (N252)? mem[8601] : 
                        (N254)? mem[8674] : 
                        (N256)? mem[8747] : 
                        (N258)? mem[8820] : 
                        (N260)? mem[8893] : 
                        (N262)? mem[8966] : 
                        (N264)? mem[9039] : 
                        (N266)? mem[9112] : 
                        (N268)? mem[9185] : 
                        (N270)? mem[9258] : 
                        (N272)? mem[9331] : 1'b0;
  assign r_data_o[59] = (N145)? mem[59] : 
                        (N147)? mem[132] : 
                        (N149)? mem[205] : 
                        (N151)? mem[278] : 
                        (N153)? mem[351] : 
                        (N155)? mem[424] : 
                        (N157)? mem[497] : 
                        (N159)? mem[570] : 
                        (N161)? mem[643] : 
                        (N163)? mem[716] : 
                        (N165)? mem[789] : 
                        (N167)? mem[862] : 
                        (N169)? mem[935] : 
                        (N171)? mem[1008] : 
                        (N173)? mem[1081] : 
                        (N175)? mem[1154] : 
                        (N177)? mem[1227] : 
                        (N179)? mem[1300] : 
                        (N181)? mem[1373] : 
                        (N183)? mem[1446] : 
                        (N185)? mem[1519] : 
                        (N187)? mem[1592] : 
                        (N189)? mem[1665] : 
                        (N191)? mem[1738] : 
                        (N193)? mem[1811] : 
                        (N195)? mem[1884] : 
                        (N197)? mem[1957] : 
                        (N199)? mem[2030] : 
                        (N201)? mem[2103] : 
                        (N203)? mem[2176] : 
                        (N205)? mem[2249] : 
                        (N207)? mem[2322] : 
                        (N209)? mem[2395] : 
                        (N211)? mem[2468] : 
                        (N213)? mem[2541] : 
                        (N215)? mem[2614] : 
                        (N217)? mem[2687] : 
                        (N219)? mem[2760] : 
                        (N221)? mem[2833] : 
                        (N223)? mem[2906] : 
                        (N225)? mem[2979] : 
                        (N227)? mem[3052] : 
                        (N229)? mem[3125] : 
                        (N231)? mem[3198] : 
                        (N233)? mem[3271] : 
                        (N235)? mem[3344] : 
                        (N237)? mem[3417] : 
                        (N239)? mem[3490] : 
                        (N241)? mem[3563] : 
                        (N243)? mem[3636] : 
                        (N245)? mem[3709] : 
                        (N247)? mem[3782] : 
                        (N249)? mem[3855] : 
                        (N251)? mem[3928] : 
                        (N253)? mem[4001] : 
                        (N255)? mem[4074] : 
                        (N257)? mem[4147] : 
                        (N259)? mem[4220] : 
                        (N261)? mem[4293] : 
                        (N263)? mem[4366] : 
                        (N265)? mem[4439] : 
                        (N267)? mem[4512] : 
                        (N269)? mem[4585] : 
                        (N271)? mem[4658] : 
                        (N146)? mem[4731] : 
                        (N148)? mem[4804] : 
                        (N150)? mem[4877] : 
                        (N152)? mem[4950] : 
                        (N154)? mem[5023] : 
                        (N156)? mem[5096] : 
                        (N158)? mem[5169] : 
                        (N160)? mem[5242] : 
                        (N162)? mem[5315] : 
                        (N164)? mem[5388] : 
                        (N166)? mem[5461] : 
                        (N168)? mem[5534] : 
                        (N170)? mem[5607] : 
                        (N172)? mem[5680] : 
                        (N174)? mem[5753] : 
                        (N176)? mem[5826] : 
                        (N178)? mem[5899] : 
                        (N180)? mem[5972] : 
                        (N182)? mem[6045] : 
                        (N184)? mem[6118] : 
                        (N186)? mem[6191] : 
                        (N188)? mem[6264] : 
                        (N190)? mem[6337] : 
                        (N192)? mem[6410] : 
                        (N194)? mem[6483] : 
                        (N196)? mem[6556] : 
                        (N198)? mem[6629] : 
                        (N200)? mem[6702] : 
                        (N202)? mem[6775] : 
                        (N204)? mem[6848] : 
                        (N206)? mem[6921] : 
                        (N208)? mem[6994] : 
                        (N210)? mem[7067] : 
                        (N212)? mem[7140] : 
                        (N214)? mem[7213] : 
                        (N216)? mem[7286] : 
                        (N218)? mem[7359] : 
                        (N220)? mem[7432] : 
                        (N222)? mem[7505] : 
                        (N224)? mem[7578] : 
                        (N226)? mem[7651] : 
                        (N228)? mem[7724] : 
                        (N230)? mem[7797] : 
                        (N232)? mem[7870] : 
                        (N234)? mem[7943] : 
                        (N236)? mem[8016] : 
                        (N238)? mem[8089] : 
                        (N240)? mem[8162] : 
                        (N242)? mem[8235] : 
                        (N244)? mem[8308] : 
                        (N246)? mem[8381] : 
                        (N248)? mem[8454] : 
                        (N250)? mem[8527] : 
                        (N252)? mem[8600] : 
                        (N254)? mem[8673] : 
                        (N256)? mem[8746] : 
                        (N258)? mem[8819] : 
                        (N260)? mem[8892] : 
                        (N262)? mem[8965] : 
                        (N264)? mem[9038] : 
                        (N266)? mem[9111] : 
                        (N268)? mem[9184] : 
                        (N270)? mem[9257] : 
                        (N272)? mem[9330] : 1'b0;
  assign r_data_o[58] = (N145)? mem[58] : 
                        (N147)? mem[131] : 
                        (N149)? mem[204] : 
                        (N151)? mem[277] : 
                        (N153)? mem[350] : 
                        (N155)? mem[423] : 
                        (N157)? mem[496] : 
                        (N159)? mem[569] : 
                        (N161)? mem[642] : 
                        (N163)? mem[715] : 
                        (N165)? mem[788] : 
                        (N167)? mem[861] : 
                        (N169)? mem[934] : 
                        (N171)? mem[1007] : 
                        (N173)? mem[1080] : 
                        (N175)? mem[1153] : 
                        (N177)? mem[1226] : 
                        (N179)? mem[1299] : 
                        (N181)? mem[1372] : 
                        (N183)? mem[1445] : 
                        (N185)? mem[1518] : 
                        (N187)? mem[1591] : 
                        (N189)? mem[1664] : 
                        (N191)? mem[1737] : 
                        (N193)? mem[1810] : 
                        (N195)? mem[1883] : 
                        (N197)? mem[1956] : 
                        (N199)? mem[2029] : 
                        (N201)? mem[2102] : 
                        (N203)? mem[2175] : 
                        (N205)? mem[2248] : 
                        (N207)? mem[2321] : 
                        (N209)? mem[2394] : 
                        (N211)? mem[2467] : 
                        (N213)? mem[2540] : 
                        (N215)? mem[2613] : 
                        (N217)? mem[2686] : 
                        (N219)? mem[2759] : 
                        (N221)? mem[2832] : 
                        (N223)? mem[2905] : 
                        (N225)? mem[2978] : 
                        (N227)? mem[3051] : 
                        (N229)? mem[3124] : 
                        (N231)? mem[3197] : 
                        (N233)? mem[3270] : 
                        (N235)? mem[3343] : 
                        (N237)? mem[3416] : 
                        (N239)? mem[3489] : 
                        (N241)? mem[3562] : 
                        (N243)? mem[3635] : 
                        (N245)? mem[3708] : 
                        (N247)? mem[3781] : 
                        (N249)? mem[3854] : 
                        (N251)? mem[3927] : 
                        (N253)? mem[4000] : 
                        (N255)? mem[4073] : 
                        (N257)? mem[4146] : 
                        (N259)? mem[4219] : 
                        (N261)? mem[4292] : 
                        (N263)? mem[4365] : 
                        (N265)? mem[4438] : 
                        (N267)? mem[4511] : 
                        (N269)? mem[4584] : 
                        (N271)? mem[4657] : 
                        (N146)? mem[4730] : 
                        (N148)? mem[4803] : 
                        (N150)? mem[4876] : 
                        (N152)? mem[4949] : 
                        (N154)? mem[5022] : 
                        (N156)? mem[5095] : 
                        (N158)? mem[5168] : 
                        (N160)? mem[5241] : 
                        (N162)? mem[5314] : 
                        (N164)? mem[5387] : 
                        (N166)? mem[5460] : 
                        (N168)? mem[5533] : 
                        (N170)? mem[5606] : 
                        (N172)? mem[5679] : 
                        (N174)? mem[5752] : 
                        (N176)? mem[5825] : 
                        (N178)? mem[5898] : 
                        (N180)? mem[5971] : 
                        (N182)? mem[6044] : 
                        (N184)? mem[6117] : 
                        (N186)? mem[6190] : 
                        (N188)? mem[6263] : 
                        (N190)? mem[6336] : 
                        (N192)? mem[6409] : 
                        (N194)? mem[6482] : 
                        (N196)? mem[6555] : 
                        (N198)? mem[6628] : 
                        (N200)? mem[6701] : 
                        (N202)? mem[6774] : 
                        (N204)? mem[6847] : 
                        (N206)? mem[6920] : 
                        (N208)? mem[6993] : 
                        (N210)? mem[7066] : 
                        (N212)? mem[7139] : 
                        (N214)? mem[7212] : 
                        (N216)? mem[7285] : 
                        (N218)? mem[7358] : 
                        (N220)? mem[7431] : 
                        (N222)? mem[7504] : 
                        (N224)? mem[7577] : 
                        (N226)? mem[7650] : 
                        (N228)? mem[7723] : 
                        (N230)? mem[7796] : 
                        (N232)? mem[7869] : 
                        (N234)? mem[7942] : 
                        (N236)? mem[8015] : 
                        (N238)? mem[8088] : 
                        (N240)? mem[8161] : 
                        (N242)? mem[8234] : 
                        (N244)? mem[8307] : 
                        (N246)? mem[8380] : 
                        (N248)? mem[8453] : 
                        (N250)? mem[8526] : 
                        (N252)? mem[8599] : 
                        (N254)? mem[8672] : 
                        (N256)? mem[8745] : 
                        (N258)? mem[8818] : 
                        (N260)? mem[8891] : 
                        (N262)? mem[8964] : 
                        (N264)? mem[9037] : 
                        (N266)? mem[9110] : 
                        (N268)? mem[9183] : 
                        (N270)? mem[9256] : 
                        (N272)? mem[9329] : 1'b0;
  assign r_data_o[57] = (N145)? mem[57] : 
                        (N147)? mem[130] : 
                        (N149)? mem[203] : 
                        (N151)? mem[276] : 
                        (N153)? mem[349] : 
                        (N155)? mem[422] : 
                        (N157)? mem[495] : 
                        (N159)? mem[568] : 
                        (N161)? mem[641] : 
                        (N163)? mem[714] : 
                        (N165)? mem[787] : 
                        (N167)? mem[860] : 
                        (N169)? mem[933] : 
                        (N171)? mem[1006] : 
                        (N173)? mem[1079] : 
                        (N175)? mem[1152] : 
                        (N177)? mem[1225] : 
                        (N179)? mem[1298] : 
                        (N181)? mem[1371] : 
                        (N183)? mem[1444] : 
                        (N185)? mem[1517] : 
                        (N187)? mem[1590] : 
                        (N189)? mem[1663] : 
                        (N191)? mem[1736] : 
                        (N193)? mem[1809] : 
                        (N195)? mem[1882] : 
                        (N197)? mem[1955] : 
                        (N199)? mem[2028] : 
                        (N201)? mem[2101] : 
                        (N203)? mem[2174] : 
                        (N205)? mem[2247] : 
                        (N207)? mem[2320] : 
                        (N209)? mem[2393] : 
                        (N211)? mem[2466] : 
                        (N213)? mem[2539] : 
                        (N215)? mem[2612] : 
                        (N217)? mem[2685] : 
                        (N219)? mem[2758] : 
                        (N221)? mem[2831] : 
                        (N223)? mem[2904] : 
                        (N225)? mem[2977] : 
                        (N227)? mem[3050] : 
                        (N229)? mem[3123] : 
                        (N231)? mem[3196] : 
                        (N233)? mem[3269] : 
                        (N235)? mem[3342] : 
                        (N237)? mem[3415] : 
                        (N239)? mem[3488] : 
                        (N241)? mem[3561] : 
                        (N243)? mem[3634] : 
                        (N245)? mem[3707] : 
                        (N247)? mem[3780] : 
                        (N249)? mem[3853] : 
                        (N251)? mem[3926] : 
                        (N253)? mem[3999] : 
                        (N255)? mem[4072] : 
                        (N257)? mem[4145] : 
                        (N259)? mem[4218] : 
                        (N261)? mem[4291] : 
                        (N263)? mem[4364] : 
                        (N265)? mem[4437] : 
                        (N267)? mem[4510] : 
                        (N269)? mem[4583] : 
                        (N271)? mem[4656] : 
                        (N146)? mem[4729] : 
                        (N148)? mem[4802] : 
                        (N150)? mem[4875] : 
                        (N152)? mem[4948] : 
                        (N154)? mem[5021] : 
                        (N156)? mem[5094] : 
                        (N158)? mem[5167] : 
                        (N160)? mem[5240] : 
                        (N162)? mem[5313] : 
                        (N164)? mem[5386] : 
                        (N166)? mem[5459] : 
                        (N168)? mem[5532] : 
                        (N170)? mem[5605] : 
                        (N172)? mem[5678] : 
                        (N174)? mem[5751] : 
                        (N176)? mem[5824] : 
                        (N178)? mem[5897] : 
                        (N180)? mem[5970] : 
                        (N182)? mem[6043] : 
                        (N184)? mem[6116] : 
                        (N186)? mem[6189] : 
                        (N188)? mem[6262] : 
                        (N190)? mem[6335] : 
                        (N192)? mem[6408] : 
                        (N194)? mem[6481] : 
                        (N196)? mem[6554] : 
                        (N198)? mem[6627] : 
                        (N200)? mem[6700] : 
                        (N202)? mem[6773] : 
                        (N204)? mem[6846] : 
                        (N206)? mem[6919] : 
                        (N208)? mem[6992] : 
                        (N210)? mem[7065] : 
                        (N212)? mem[7138] : 
                        (N214)? mem[7211] : 
                        (N216)? mem[7284] : 
                        (N218)? mem[7357] : 
                        (N220)? mem[7430] : 
                        (N222)? mem[7503] : 
                        (N224)? mem[7576] : 
                        (N226)? mem[7649] : 
                        (N228)? mem[7722] : 
                        (N230)? mem[7795] : 
                        (N232)? mem[7868] : 
                        (N234)? mem[7941] : 
                        (N236)? mem[8014] : 
                        (N238)? mem[8087] : 
                        (N240)? mem[8160] : 
                        (N242)? mem[8233] : 
                        (N244)? mem[8306] : 
                        (N246)? mem[8379] : 
                        (N248)? mem[8452] : 
                        (N250)? mem[8525] : 
                        (N252)? mem[8598] : 
                        (N254)? mem[8671] : 
                        (N256)? mem[8744] : 
                        (N258)? mem[8817] : 
                        (N260)? mem[8890] : 
                        (N262)? mem[8963] : 
                        (N264)? mem[9036] : 
                        (N266)? mem[9109] : 
                        (N268)? mem[9182] : 
                        (N270)? mem[9255] : 
                        (N272)? mem[9328] : 1'b0;
  assign r_data_o[56] = (N145)? mem[56] : 
                        (N147)? mem[129] : 
                        (N149)? mem[202] : 
                        (N151)? mem[275] : 
                        (N153)? mem[348] : 
                        (N155)? mem[421] : 
                        (N157)? mem[494] : 
                        (N159)? mem[567] : 
                        (N161)? mem[640] : 
                        (N163)? mem[713] : 
                        (N165)? mem[786] : 
                        (N167)? mem[859] : 
                        (N169)? mem[932] : 
                        (N171)? mem[1005] : 
                        (N173)? mem[1078] : 
                        (N175)? mem[1151] : 
                        (N177)? mem[1224] : 
                        (N179)? mem[1297] : 
                        (N181)? mem[1370] : 
                        (N183)? mem[1443] : 
                        (N185)? mem[1516] : 
                        (N187)? mem[1589] : 
                        (N189)? mem[1662] : 
                        (N191)? mem[1735] : 
                        (N193)? mem[1808] : 
                        (N195)? mem[1881] : 
                        (N197)? mem[1954] : 
                        (N199)? mem[2027] : 
                        (N201)? mem[2100] : 
                        (N203)? mem[2173] : 
                        (N205)? mem[2246] : 
                        (N207)? mem[2319] : 
                        (N209)? mem[2392] : 
                        (N211)? mem[2465] : 
                        (N213)? mem[2538] : 
                        (N215)? mem[2611] : 
                        (N217)? mem[2684] : 
                        (N219)? mem[2757] : 
                        (N221)? mem[2830] : 
                        (N223)? mem[2903] : 
                        (N225)? mem[2976] : 
                        (N227)? mem[3049] : 
                        (N229)? mem[3122] : 
                        (N231)? mem[3195] : 
                        (N233)? mem[3268] : 
                        (N235)? mem[3341] : 
                        (N237)? mem[3414] : 
                        (N239)? mem[3487] : 
                        (N241)? mem[3560] : 
                        (N243)? mem[3633] : 
                        (N245)? mem[3706] : 
                        (N247)? mem[3779] : 
                        (N249)? mem[3852] : 
                        (N251)? mem[3925] : 
                        (N253)? mem[3998] : 
                        (N255)? mem[4071] : 
                        (N257)? mem[4144] : 
                        (N259)? mem[4217] : 
                        (N261)? mem[4290] : 
                        (N263)? mem[4363] : 
                        (N265)? mem[4436] : 
                        (N267)? mem[4509] : 
                        (N269)? mem[4582] : 
                        (N271)? mem[4655] : 
                        (N146)? mem[4728] : 
                        (N148)? mem[4801] : 
                        (N150)? mem[4874] : 
                        (N152)? mem[4947] : 
                        (N154)? mem[5020] : 
                        (N156)? mem[5093] : 
                        (N158)? mem[5166] : 
                        (N160)? mem[5239] : 
                        (N162)? mem[5312] : 
                        (N164)? mem[5385] : 
                        (N166)? mem[5458] : 
                        (N168)? mem[5531] : 
                        (N170)? mem[5604] : 
                        (N172)? mem[5677] : 
                        (N174)? mem[5750] : 
                        (N176)? mem[5823] : 
                        (N178)? mem[5896] : 
                        (N180)? mem[5969] : 
                        (N182)? mem[6042] : 
                        (N184)? mem[6115] : 
                        (N186)? mem[6188] : 
                        (N188)? mem[6261] : 
                        (N190)? mem[6334] : 
                        (N192)? mem[6407] : 
                        (N194)? mem[6480] : 
                        (N196)? mem[6553] : 
                        (N198)? mem[6626] : 
                        (N200)? mem[6699] : 
                        (N202)? mem[6772] : 
                        (N204)? mem[6845] : 
                        (N206)? mem[6918] : 
                        (N208)? mem[6991] : 
                        (N210)? mem[7064] : 
                        (N212)? mem[7137] : 
                        (N214)? mem[7210] : 
                        (N216)? mem[7283] : 
                        (N218)? mem[7356] : 
                        (N220)? mem[7429] : 
                        (N222)? mem[7502] : 
                        (N224)? mem[7575] : 
                        (N226)? mem[7648] : 
                        (N228)? mem[7721] : 
                        (N230)? mem[7794] : 
                        (N232)? mem[7867] : 
                        (N234)? mem[7940] : 
                        (N236)? mem[8013] : 
                        (N238)? mem[8086] : 
                        (N240)? mem[8159] : 
                        (N242)? mem[8232] : 
                        (N244)? mem[8305] : 
                        (N246)? mem[8378] : 
                        (N248)? mem[8451] : 
                        (N250)? mem[8524] : 
                        (N252)? mem[8597] : 
                        (N254)? mem[8670] : 
                        (N256)? mem[8743] : 
                        (N258)? mem[8816] : 
                        (N260)? mem[8889] : 
                        (N262)? mem[8962] : 
                        (N264)? mem[9035] : 
                        (N266)? mem[9108] : 
                        (N268)? mem[9181] : 
                        (N270)? mem[9254] : 
                        (N272)? mem[9327] : 1'b0;
  assign r_data_o[55] = (N145)? mem[55] : 
                        (N147)? mem[128] : 
                        (N149)? mem[201] : 
                        (N151)? mem[274] : 
                        (N153)? mem[347] : 
                        (N155)? mem[420] : 
                        (N157)? mem[493] : 
                        (N159)? mem[566] : 
                        (N161)? mem[639] : 
                        (N163)? mem[712] : 
                        (N165)? mem[785] : 
                        (N167)? mem[858] : 
                        (N169)? mem[931] : 
                        (N171)? mem[1004] : 
                        (N173)? mem[1077] : 
                        (N175)? mem[1150] : 
                        (N177)? mem[1223] : 
                        (N179)? mem[1296] : 
                        (N181)? mem[1369] : 
                        (N183)? mem[1442] : 
                        (N185)? mem[1515] : 
                        (N187)? mem[1588] : 
                        (N189)? mem[1661] : 
                        (N191)? mem[1734] : 
                        (N193)? mem[1807] : 
                        (N195)? mem[1880] : 
                        (N197)? mem[1953] : 
                        (N199)? mem[2026] : 
                        (N201)? mem[2099] : 
                        (N203)? mem[2172] : 
                        (N205)? mem[2245] : 
                        (N207)? mem[2318] : 
                        (N209)? mem[2391] : 
                        (N211)? mem[2464] : 
                        (N213)? mem[2537] : 
                        (N215)? mem[2610] : 
                        (N217)? mem[2683] : 
                        (N219)? mem[2756] : 
                        (N221)? mem[2829] : 
                        (N223)? mem[2902] : 
                        (N225)? mem[2975] : 
                        (N227)? mem[3048] : 
                        (N229)? mem[3121] : 
                        (N231)? mem[3194] : 
                        (N233)? mem[3267] : 
                        (N235)? mem[3340] : 
                        (N237)? mem[3413] : 
                        (N239)? mem[3486] : 
                        (N241)? mem[3559] : 
                        (N243)? mem[3632] : 
                        (N245)? mem[3705] : 
                        (N247)? mem[3778] : 
                        (N249)? mem[3851] : 
                        (N251)? mem[3924] : 
                        (N253)? mem[3997] : 
                        (N255)? mem[4070] : 
                        (N257)? mem[4143] : 
                        (N259)? mem[4216] : 
                        (N261)? mem[4289] : 
                        (N263)? mem[4362] : 
                        (N265)? mem[4435] : 
                        (N267)? mem[4508] : 
                        (N269)? mem[4581] : 
                        (N271)? mem[4654] : 
                        (N146)? mem[4727] : 
                        (N148)? mem[4800] : 
                        (N150)? mem[4873] : 
                        (N152)? mem[4946] : 
                        (N154)? mem[5019] : 
                        (N156)? mem[5092] : 
                        (N158)? mem[5165] : 
                        (N160)? mem[5238] : 
                        (N162)? mem[5311] : 
                        (N164)? mem[5384] : 
                        (N166)? mem[5457] : 
                        (N168)? mem[5530] : 
                        (N170)? mem[5603] : 
                        (N172)? mem[5676] : 
                        (N174)? mem[5749] : 
                        (N176)? mem[5822] : 
                        (N178)? mem[5895] : 
                        (N180)? mem[5968] : 
                        (N182)? mem[6041] : 
                        (N184)? mem[6114] : 
                        (N186)? mem[6187] : 
                        (N188)? mem[6260] : 
                        (N190)? mem[6333] : 
                        (N192)? mem[6406] : 
                        (N194)? mem[6479] : 
                        (N196)? mem[6552] : 
                        (N198)? mem[6625] : 
                        (N200)? mem[6698] : 
                        (N202)? mem[6771] : 
                        (N204)? mem[6844] : 
                        (N206)? mem[6917] : 
                        (N208)? mem[6990] : 
                        (N210)? mem[7063] : 
                        (N212)? mem[7136] : 
                        (N214)? mem[7209] : 
                        (N216)? mem[7282] : 
                        (N218)? mem[7355] : 
                        (N220)? mem[7428] : 
                        (N222)? mem[7501] : 
                        (N224)? mem[7574] : 
                        (N226)? mem[7647] : 
                        (N228)? mem[7720] : 
                        (N230)? mem[7793] : 
                        (N232)? mem[7866] : 
                        (N234)? mem[7939] : 
                        (N236)? mem[8012] : 
                        (N238)? mem[8085] : 
                        (N240)? mem[8158] : 
                        (N242)? mem[8231] : 
                        (N244)? mem[8304] : 
                        (N246)? mem[8377] : 
                        (N248)? mem[8450] : 
                        (N250)? mem[8523] : 
                        (N252)? mem[8596] : 
                        (N254)? mem[8669] : 
                        (N256)? mem[8742] : 
                        (N258)? mem[8815] : 
                        (N260)? mem[8888] : 
                        (N262)? mem[8961] : 
                        (N264)? mem[9034] : 
                        (N266)? mem[9107] : 
                        (N268)? mem[9180] : 
                        (N270)? mem[9253] : 
                        (N272)? mem[9326] : 1'b0;
  assign r_data_o[54] = (N145)? mem[54] : 
                        (N147)? mem[127] : 
                        (N149)? mem[200] : 
                        (N151)? mem[273] : 
                        (N153)? mem[346] : 
                        (N155)? mem[419] : 
                        (N157)? mem[492] : 
                        (N159)? mem[565] : 
                        (N161)? mem[638] : 
                        (N163)? mem[711] : 
                        (N165)? mem[784] : 
                        (N167)? mem[857] : 
                        (N169)? mem[930] : 
                        (N171)? mem[1003] : 
                        (N173)? mem[1076] : 
                        (N175)? mem[1149] : 
                        (N177)? mem[1222] : 
                        (N179)? mem[1295] : 
                        (N181)? mem[1368] : 
                        (N183)? mem[1441] : 
                        (N185)? mem[1514] : 
                        (N187)? mem[1587] : 
                        (N189)? mem[1660] : 
                        (N191)? mem[1733] : 
                        (N193)? mem[1806] : 
                        (N195)? mem[1879] : 
                        (N197)? mem[1952] : 
                        (N199)? mem[2025] : 
                        (N201)? mem[2098] : 
                        (N203)? mem[2171] : 
                        (N205)? mem[2244] : 
                        (N207)? mem[2317] : 
                        (N209)? mem[2390] : 
                        (N211)? mem[2463] : 
                        (N213)? mem[2536] : 
                        (N215)? mem[2609] : 
                        (N217)? mem[2682] : 
                        (N219)? mem[2755] : 
                        (N221)? mem[2828] : 
                        (N223)? mem[2901] : 
                        (N225)? mem[2974] : 
                        (N227)? mem[3047] : 
                        (N229)? mem[3120] : 
                        (N231)? mem[3193] : 
                        (N233)? mem[3266] : 
                        (N235)? mem[3339] : 
                        (N237)? mem[3412] : 
                        (N239)? mem[3485] : 
                        (N241)? mem[3558] : 
                        (N243)? mem[3631] : 
                        (N245)? mem[3704] : 
                        (N247)? mem[3777] : 
                        (N249)? mem[3850] : 
                        (N251)? mem[3923] : 
                        (N253)? mem[3996] : 
                        (N255)? mem[4069] : 
                        (N257)? mem[4142] : 
                        (N259)? mem[4215] : 
                        (N261)? mem[4288] : 
                        (N263)? mem[4361] : 
                        (N265)? mem[4434] : 
                        (N267)? mem[4507] : 
                        (N269)? mem[4580] : 
                        (N271)? mem[4653] : 
                        (N146)? mem[4726] : 
                        (N148)? mem[4799] : 
                        (N150)? mem[4872] : 
                        (N152)? mem[4945] : 
                        (N154)? mem[5018] : 
                        (N156)? mem[5091] : 
                        (N158)? mem[5164] : 
                        (N160)? mem[5237] : 
                        (N162)? mem[5310] : 
                        (N164)? mem[5383] : 
                        (N166)? mem[5456] : 
                        (N168)? mem[5529] : 
                        (N170)? mem[5602] : 
                        (N172)? mem[5675] : 
                        (N174)? mem[5748] : 
                        (N176)? mem[5821] : 
                        (N178)? mem[5894] : 
                        (N180)? mem[5967] : 
                        (N182)? mem[6040] : 
                        (N184)? mem[6113] : 
                        (N186)? mem[6186] : 
                        (N188)? mem[6259] : 
                        (N190)? mem[6332] : 
                        (N192)? mem[6405] : 
                        (N194)? mem[6478] : 
                        (N196)? mem[6551] : 
                        (N198)? mem[6624] : 
                        (N200)? mem[6697] : 
                        (N202)? mem[6770] : 
                        (N204)? mem[6843] : 
                        (N206)? mem[6916] : 
                        (N208)? mem[6989] : 
                        (N210)? mem[7062] : 
                        (N212)? mem[7135] : 
                        (N214)? mem[7208] : 
                        (N216)? mem[7281] : 
                        (N218)? mem[7354] : 
                        (N220)? mem[7427] : 
                        (N222)? mem[7500] : 
                        (N224)? mem[7573] : 
                        (N226)? mem[7646] : 
                        (N228)? mem[7719] : 
                        (N230)? mem[7792] : 
                        (N232)? mem[7865] : 
                        (N234)? mem[7938] : 
                        (N236)? mem[8011] : 
                        (N238)? mem[8084] : 
                        (N240)? mem[8157] : 
                        (N242)? mem[8230] : 
                        (N244)? mem[8303] : 
                        (N246)? mem[8376] : 
                        (N248)? mem[8449] : 
                        (N250)? mem[8522] : 
                        (N252)? mem[8595] : 
                        (N254)? mem[8668] : 
                        (N256)? mem[8741] : 
                        (N258)? mem[8814] : 
                        (N260)? mem[8887] : 
                        (N262)? mem[8960] : 
                        (N264)? mem[9033] : 
                        (N266)? mem[9106] : 
                        (N268)? mem[9179] : 
                        (N270)? mem[9252] : 
                        (N272)? mem[9325] : 1'b0;
  assign r_data_o[53] = (N145)? mem[53] : 
                        (N147)? mem[126] : 
                        (N149)? mem[199] : 
                        (N151)? mem[272] : 
                        (N153)? mem[345] : 
                        (N155)? mem[418] : 
                        (N157)? mem[491] : 
                        (N159)? mem[564] : 
                        (N161)? mem[637] : 
                        (N163)? mem[710] : 
                        (N165)? mem[783] : 
                        (N167)? mem[856] : 
                        (N169)? mem[929] : 
                        (N171)? mem[1002] : 
                        (N173)? mem[1075] : 
                        (N175)? mem[1148] : 
                        (N177)? mem[1221] : 
                        (N179)? mem[1294] : 
                        (N181)? mem[1367] : 
                        (N183)? mem[1440] : 
                        (N185)? mem[1513] : 
                        (N187)? mem[1586] : 
                        (N189)? mem[1659] : 
                        (N191)? mem[1732] : 
                        (N193)? mem[1805] : 
                        (N195)? mem[1878] : 
                        (N197)? mem[1951] : 
                        (N199)? mem[2024] : 
                        (N201)? mem[2097] : 
                        (N203)? mem[2170] : 
                        (N205)? mem[2243] : 
                        (N207)? mem[2316] : 
                        (N209)? mem[2389] : 
                        (N211)? mem[2462] : 
                        (N213)? mem[2535] : 
                        (N215)? mem[2608] : 
                        (N217)? mem[2681] : 
                        (N219)? mem[2754] : 
                        (N221)? mem[2827] : 
                        (N223)? mem[2900] : 
                        (N225)? mem[2973] : 
                        (N227)? mem[3046] : 
                        (N229)? mem[3119] : 
                        (N231)? mem[3192] : 
                        (N233)? mem[3265] : 
                        (N235)? mem[3338] : 
                        (N237)? mem[3411] : 
                        (N239)? mem[3484] : 
                        (N241)? mem[3557] : 
                        (N243)? mem[3630] : 
                        (N245)? mem[3703] : 
                        (N247)? mem[3776] : 
                        (N249)? mem[3849] : 
                        (N251)? mem[3922] : 
                        (N253)? mem[3995] : 
                        (N255)? mem[4068] : 
                        (N257)? mem[4141] : 
                        (N259)? mem[4214] : 
                        (N261)? mem[4287] : 
                        (N263)? mem[4360] : 
                        (N265)? mem[4433] : 
                        (N267)? mem[4506] : 
                        (N269)? mem[4579] : 
                        (N271)? mem[4652] : 
                        (N146)? mem[4725] : 
                        (N148)? mem[4798] : 
                        (N150)? mem[4871] : 
                        (N152)? mem[4944] : 
                        (N154)? mem[5017] : 
                        (N156)? mem[5090] : 
                        (N158)? mem[5163] : 
                        (N160)? mem[5236] : 
                        (N162)? mem[5309] : 
                        (N164)? mem[5382] : 
                        (N166)? mem[5455] : 
                        (N168)? mem[5528] : 
                        (N170)? mem[5601] : 
                        (N172)? mem[5674] : 
                        (N174)? mem[5747] : 
                        (N176)? mem[5820] : 
                        (N178)? mem[5893] : 
                        (N180)? mem[5966] : 
                        (N182)? mem[6039] : 
                        (N184)? mem[6112] : 
                        (N186)? mem[6185] : 
                        (N188)? mem[6258] : 
                        (N190)? mem[6331] : 
                        (N192)? mem[6404] : 
                        (N194)? mem[6477] : 
                        (N196)? mem[6550] : 
                        (N198)? mem[6623] : 
                        (N200)? mem[6696] : 
                        (N202)? mem[6769] : 
                        (N204)? mem[6842] : 
                        (N206)? mem[6915] : 
                        (N208)? mem[6988] : 
                        (N210)? mem[7061] : 
                        (N212)? mem[7134] : 
                        (N214)? mem[7207] : 
                        (N216)? mem[7280] : 
                        (N218)? mem[7353] : 
                        (N220)? mem[7426] : 
                        (N222)? mem[7499] : 
                        (N224)? mem[7572] : 
                        (N226)? mem[7645] : 
                        (N228)? mem[7718] : 
                        (N230)? mem[7791] : 
                        (N232)? mem[7864] : 
                        (N234)? mem[7937] : 
                        (N236)? mem[8010] : 
                        (N238)? mem[8083] : 
                        (N240)? mem[8156] : 
                        (N242)? mem[8229] : 
                        (N244)? mem[8302] : 
                        (N246)? mem[8375] : 
                        (N248)? mem[8448] : 
                        (N250)? mem[8521] : 
                        (N252)? mem[8594] : 
                        (N254)? mem[8667] : 
                        (N256)? mem[8740] : 
                        (N258)? mem[8813] : 
                        (N260)? mem[8886] : 
                        (N262)? mem[8959] : 
                        (N264)? mem[9032] : 
                        (N266)? mem[9105] : 
                        (N268)? mem[9178] : 
                        (N270)? mem[9251] : 
                        (N272)? mem[9324] : 1'b0;
  assign r_data_o[52] = (N145)? mem[52] : 
                        (N147)? mem[125] : 
                        (N149)? mem[198] : 
                        (N151)? mem[271] : 
                        (N153)? mem[344] : 
                        (N155)? mem[417] : 
                        (N157)? mem[490] : 
                        (N159)? mem[563] : 
                        (N161)? mem[636] : 
                        (N163)? mem[709] : 
                        (N165)? mem[782] : 
                        (N167)? mem[855] : 
                        (N169)? mem[928] : 
                        (N171)? mem[1001] : 
                        (N173)? mem[1074] : 
                        (N175)? mem[1147] : 
                        (N177)? mem[1220] : 
                        (N179)? mem[1293] : 
                        (N181)? mem[1366] : 
                        (N183)? mem[1439] : 
                        (N185)? mem[1512] : 
                        (N187)? mem[1585] : 
                        (N189)? mem[1658] : 
                        (N191)? mem[1731] : 
                        (N193)? mem[1804] : 
                        (N195)? mem[1877] : 
                        (N197)? mem[1950] : 
                        (N199)? mem[2023] : 
                        (N201)? mem[2096] : 
                        (N203)? mem[2169] : 
                        (N205)? mem[2242] : 
                        (N207)? mem[2315] : 
                        (N209)? mem[2388] : 
                        (N211)? mem[2461] : 
                        (N213)? mem[2534] : 
                        (N215)? mem[2607] : 
                        (N217)? mem[2680] : 
                        (N219)? mem[2753] : 
                        (N221)? mem[2826] : 
                        (N223)? mem[2899] : 
                        (N225)? mem[2972] : 
                        (N227)? mem[3045] : 
                        (N229)? mem[3118] : 
                        (N231)? mem[3191] : 
                        (N233)? mem[3264] : 
                        (N235)? mem[3337] : 
                        (N237)? mem[3410] : 
                        (N239)? mem[3483] : 
                        (N241)? mem[3556] : 
                        (N243)? mem[3629] : 
                        (N245)? mem[3702] : 
                        (N247)? mem[3775] : 
                        (N249)? mem[3848] : 
                        (N251)? mem[3921] : 
                        (N253)? mem[3994] : 
                        (N255)? mem[4067] : 
                        (N257)? mem[4140] : 
                        (N259)? mem[4213] : 
                        (N261)? mem[4286] : 
                        (N263)? mem[4359] : 
                        (N265)? mem[4432] : 
                        (N267)? mem[4505] : 
                        (N269)? mem[4578] : 
                        (N271)? mem[4651] : 
                        (N146)? mem[4724] : 
                        (N148)? mem[4797] : 
                        (N150)? mem[4870] : 
                        (N152)? mem[4943] : 
                        (N154)? mem[5016] : 
                        (N156)? mem[5089] : 
                        (N158)? mem[5162] : 
                        (N160)? mem[5235] : 
                        (N162)? mem[5308] : 
                        (N164)? mem[5381] : 
                        (N166)? mem[5454] : 
                        (N168)? mem[5527] : 
                        (N170)? mem[5600] : 
                        (N172)? mem[5673] : 
                        (N174)? mem[5746] : 
                        (N176)? mem[5819] : 
                        (N178)? mem[5892] : 
                        (N180)? mem[5965] : 
                        (N182)? mem[6038] : 
                        (N184)? mem[6111] : 
                        (N186)? mem[6184] : 
                        (N188)? mem[6257] : 
                        (N190)? mem[6330] : 
                        (N192)? mem[6403] : 
                        (N194)? mem[6476] : 
                        (N196)? mem[6549] : 
                        (N198)? mem[6622] : 
                        (N200)? mem[6695] : 
                        (N202)? mem[6768] : 
                        (N204)? mem[6841] : 
                        (N206)? mem[6914] : 
                        (N208)? mem[6987] : 
                        (N210)? mem[7060] : 
                        (N212)? mem[7133] : 
                        (N214)? mem[7206] : 
                        (N216)? mem[7279] : 
                        (N218)? mem[7352] : 
                        (N220)? mem[7425] : 
                        (N222)? mem[7498] : 
                        (N224)? mem[7571] : 
                        (N226)? mem[7644] : 
                        (N228)? mem[7717] : 
                        (N230)? mem[7790] : 
                        (N232)? mem[7863] : 
                        (N234)? mem[7936] : 
                        (N236)? mem[8009] : 
                        (N238)? mem[8082] : 
                        (N240)? mem[8155] : 
                        (N242)? mem[8228] : 
                        (N244)? mem[8301] : 
                        (N246)? mem[8374] : 
                        (N248)? mem[8447] : 
                        (N250)? mem[8520] : 
                        (N252)? mem[8593] : 
                        (N254)? mem[8666] : 
                        (N256)? mem[8739] : 
                        (N258)? mem[8812] : 
                        (N260)? mem[8885] : 
                        (N262)? mem[8958] : 
                        (N264)? mem[9031] : 
                        (N266)? mem[9104] : 
                        (N268)? mem[9177] : 
                        (N270)? mem[9250] : 
                        (N272)? mem[9323] : 1'b0;
  assign r_data_o[51] = (N145)? mem[51] : 
                        (N147)? mem[124] : 
                        (N149)? mem[197] : 
                        (N151)? mem[270] : 
                        (N153)? mem[343] : 
                        (N155)? mem[416] : 
                        (N157)? mem[489] : 
                        (N159)? mem[562] : 
                        (N161)? mem[635] : 
                        (N163)? mem[708] : 
                        (N165)? mem[781] : 
                        (N167)? mem[854] : 
                        (N169)? mem[927] : 
                        (N171)? mem[1000] : 
                        (N173)? mem[1073] : 
                        (N175)? mem[1146] : 
                        (N177)? mem[1219] : 
                        (N179)? mem[1292] : 
                        (N181)? mem[1365] : 
                        (N183)? mem[1438] : 
                        (N185)? mem[1511] : 
                        (N187)? mem[1584] : 
                        (N189)? mem[1657] : 
                        (N191)? mem[1730] : 
                        (N193)? mem[1803] : 
                        (N195)? mem[1876] : 
                        (N197)? mem[1949] : 
                        (N199)? mem[2022] : 
                        (N201)? mem[2095] : 
                        (N203)? mem[2168] : 
                        (N205)? mem[2241] : 
                        (N207)? mem[2314] : 
                        (N209)? mem[2387] : 
                        (N211)? mem[2460] : 
                        (N213)? mem[2533] : 
                        (N215)? mem[2606] : 
                        (N217)? mem[2679] : 
                        (N219)? mem[2752] : 
                        (N221)? mem[2825] : 
                        (N223)? mem[2898] : 
                        (N225)? mem[2971] : 
                        (N227)? mem[3044] : 
                        (N229)? mem[3117] : 
                        (N231)? mem[3190] : 
                        (N233)? mem[3263] : 
                        (N235)? mem[3336] : 
                        (N237)? mem[3409] : 
                        (N239)? mem[3482] : 
                        (N241)? mem[3555] : 
                        (N243)? mem[3628] : 
                        (N245)? mem[3701] : 
                        (N247)? mem[3774] : 
                        (N249)? mem[3847] : 
                        (N251)? mem[3920] : 
                        (N253)? mem[3993] : 
                        (N255)? mem[4066] : 
                        (N257)? mem[4139] : 
                        (N259)? mem[4212] : 
                        (N261)? mem[4285] : 
                        (N263)? mem[4358] : 
                        (N265)? mem[4431] : 
                        (N267)? mem[4504] : 
                        (N269)? mem[4577] : 
                        (N271)? mem[4650] : 
                        (N146)? mem[4723] : 
                        (N148)? mem[4796] : 
                        (N150)? mem[4869] : 
                        (N152)? mem[4942] : 
                        (N154)? mem[5015] : 
                        (N156)? mem[5088] : 
                        (N158)? mem[5161] : 
                        (N160)? mem[5234] : 
                        (N162)? mem[5307] : 
                        (N164)? mem[5380] : 
                        (N166)? mem[5453] : 
                        (N168)? mem[5526] : 
                        (N170)? mem[5599] : 
                        (N172)? mem[5672] : 
                        (N174)? mem[5745] : 
                        (N176)? mem[5818] : 
                        (N178)? mem[5891] : 
                        (N180)? mem[5964] : 
                        (N182)? mem[6037] : 
                        (N184)? mem[6110] : 
                        (N186)? mem[6183] : 
                        (N188)? mem[6256] : 
                        (N190)? mem[6329] : 
                        (N192)? mem[6402] : 
                        (N194)? mem[6475] : 
                        (N196)? mem[6548] : 
                        (N198)? mem[6621] : 
                        (N200)? mem[6694] : 
                        (N202)? mem[6767] : 
                        (N204)? mem[6840] : 
                        (N206)? mem[6913] : 
                        (N208)? mem[6986] : 
                        (N210)? mem[7059] : 
                        (N212)? mem[7132] : 
                        (N214)? mem[7205] : 
                        (N216)? mem[7278] : 
                        (N218)? mem[7351] : 
                        (N220)? mem[7424] : 
                        (N222)? mem[7497] : 
                        (N224)? mem[7570] : 
                        (N226)? mem[7643] : 
                        (N228)? mem[7716] : 
                        (N230)? mem[7789] : 
                        (N232)? mem[7862] : 
                        (N234)? mem[7935] : 
                        (N236)? mem[8008] : 
                        (N238)? mem[8081] : 
                        (N240)? mem[8154] : 
                        (N242)? mem[8227] : 
                        (N244)? mem[8300] : 
                        (N246)? mem[8373] : 
                        (N248)? mem[8446] : 
                        (N250)? mem[8519] : 
                        (N252)? mem[8592] : 
                        (N254)? mem[8665] : 
                        (N256)? mem[8738] : 
                        (N258)? mem[8811] : 
                        (N260)? mem[8884] : 
                        (N262)? mem[8957] : 
                        (N264)? mem[9030] : 
                        (N266)? mem[9103] : 
                        (N268)? mem[9176] : 
                        (N270)? mem[9249] : 
                        (N272)? mem[9322] : 1'b0;
  assign r_data_o[50] = (N145)? mem[50] : 
                        (N147)? mem[123] : 
                        (N149)? mem[196] : 
                        (N151)? mem[269] : 
                        (N153)? mem[342] : 
                        (N155)? mem[415] : 
                        (N157)? mem[488] : 
                        (N159)? mem[561] : 
                        (N161)? mem[634] : 
                        (N163)? mem[707] : 
                        (N165)? mem[780] : 
                        (N167)? mem[853] : 
                        (N169)? mem[926] : 
                        (N171)? mem[999] : 
                        (N173)? mem[1072] : 
                        (N175)? mem[1145] : 
                        (N177)? mem[1218] : 
                        (N179)? mem[1291] : 
                        (N181)? mem[1364] : 
                        (N183)? mem[1437] : 
                        (N185)? mem[1510] : 
                        (N187)? mem[1583] : 
                        (N189)? mem[1656] : 
                        (N191)? mem[1729] : 
                        (N193)? mem[1802] : 
                        (N195)? mem[1875] : 
                        (N197)? mem[1948] : 
                        (N199)? mem[2021] : 
                        (N201)? mem[2094] : 
                        (N203)? mem[2167] : 
                        (N205)? mem[2240] : 
                        (N207)? mem[2313] : 
                        (N209)? mem[2386] : 
                        (N211)? mem[2459] : 
                        (N213)? mem[2532] : 
                        (N215)? mem[2605] : 
                        (N217)? mem[2678] : 
                        (N219)? mem[2751] : 
                        (N221)? mem[2824] : 
                        (N223)? mem[2897] : 
                        (N225)? mem[2970] : 
                        (N227)? mem[3043] : 
                        (N229)? mem[3116] : 
                        (N231)? mem[3189] : 
                        (N233)? mem[3262] : 
                        (N235)? mem[3335] : 
                        (N237)? mem[3408] : 
                        (N239)? mem[3481] : 
                        (N241)? mem[3554] : 
                        (N243)? mem[3627] : 
                        (N245)? mem[3700] : 
                        (N247)? mem[3773] : 
                        (N249)? mem[3846] : 
                        (N251)? mem[3919] : 
                        (N253)? mem[3992] : 
                        (N255)? mem[4065] : 
                        (N257)? mem[4138] : 
                        (N259)? mem[4211] : 
                        (N261)? mem[4284] : 
                        (N263)? mem[4357] : 
                        (N265)? mem[4430] : 
                        (N267)? mem[4503] : 
                        (N269)? mem[4576] : 
                        (N271)? mem[4649] : 
                        (N146)? mem[4722] : 
                        (N148)? mem[4795] : 
                        (N150)? mem[4868] : 
                        (N152)? mem[4941] : 
                        (N154)? mem[5014] : 
                        (N156)? mem[5087] : 
                        (N158)? mem[5160] : 
                        (N160)? mem[5233] : 
                        (N162)? mem[5306] : 
                        (N164)? mem[5379] : 
                        (N166)? mem[5452] : 
                        (N168)? mem[5525] : 
                        (N170)? mem[5598] : 
                        (N172)? mem[5671] : 
                        (N174)? mem[5744] : 
                        (N176)? mem[5817] : 
                        (N178)? mem[5890] : 
                        (N180)? mem[5963] : 
                        (N182)? mem[6036] : 
                        (N184)? mem[6109] : 
                        (N186)? mem[6182] : 
                        (N188)? mem[6255] : 
                        (N190)? mem[6328] : 
                        (N192)? mem[6401] : 
                        (N194)? mem[6474] : 
                        (N196)? mem[6547] : 
                        (N198)? mem[6620] : 
                        (N200)? mem[6693] : 
                        (N202)? mem[6766] : 
                        (N204)? mem[6839] : 
                        (N206)? mem[6912] : 
                        (N208)? mem[6985] : 
                        (N210)? mem[7058] : 
                        (N212)? mem[7131] : 
                        (N214)? mem[7204] : 
                        (N216)? mem[7277] : 
                        (N218)? mem[7350] : 
                        (N220)? mem[7423] : 
                        (N222)? mem[7496] : 
                        (N224)? mem[7569] : 
                        (N226)? mem[7642] : 
                        (N228)? mem[7715] : 
                        (N230)? mem[7788] : 
                        (N232)? mem[7861] : 
                        (N234)? mem[7934] : 
                        (N236)? mem[8007] : 
                        (N238)? mem[8080] : 
                        (N240)? mem[8153] : 
                        (N242)? mem[8226] : 
                        (N244)? mem[8299] : 
                        (N246)? mem[8372] : 
                        (N248)? mem[8445] : 
                        (N250)? mem[8518] : 
                        (N252)? mem[8591] : 
                        (N254)? mem[8664] : 
                        (N256)? mem[8737] : 
                        (N258)? mem[8810] : 
                        (N260)? mem[8883] : 
                        (N262)? mem[8956] : 
                        (N264)? mem[9029] : 
                        (N266)? mem[9102] : 
                        (N268)? mem[9175] : 
                        (N270)? mem[9248] : 
                        (N272)? mem[9321] : 1'b0;
  assign r_data_o[49] = (N145)? mem[49] : 
                        (N147)? mem[122] : 
                        (N149)? mem[195] : 
                        (N151)? mem[268] : 
                        (N153)? mem[341] : 
                        (N155)? mem[414] : 
                        (N157)? mem[487] : 
                        (N159)? mem[560] : 
                        (N161)? mem[633] : 
                        (N163)? mem[706] : 
                        (N165)? mem[779] : 
                        (N167)? mem[852] : 
                        (N169)? mem[925] : 
                        (N171)? mem[998] : 
                        (N173)? mem[1071] : 
                        (N175)? mem[1144] : 
                        (N177)? mem[1217] : 
                        (N179)? mem[1290] : 
                        (N181)? mem[1363] : 
                        (N183)? mem[1436] : 
                        (N185)? mem[1509] : 
                        (N187)? mem[1582] : 
                        (N189)? mem[1655] : 
                        (N191)? mem[1728] : 
                        (N193)? mem[1801] : 
                        (N195)? mem[1874] : 
                        (N197)? mem[1947] : 
                        (N199)? mem[2020] : 
                        (N201)? mem[2093] : 
                        (N203)? mem[2166] : 
                        (N205)? mem[2239] : 
                        (N207)? mem[2312] : 
                        (N209)? mem[2385] : 
                        (N211)? mem[2458] : 
                        (N213)? mem[2531] : 
                        (N215)? mem[2604] : 
                        (N217)? mem[2677] : 
                        (N219)? mem[2750] : 
                        (N221)? mem[2823] : 
                        (N223)? mem[2896] : 
                        (N225)? mem[2969] : 
                        (N227)? mem[3042] : 
                        (N229)? mem[3115] : 
                        (N231)? mem[3188] : 
                        (N233)? mem[3261] : 
                        (N235)? mem[3334] : 
                        (N237)? mem[3407] : 
                        (N239)? mem[3480] : 
                        (N241)? mem[3553] : 
                        (N243)? mem[3626] : 
                        (N245)? mem[3699] : 
                        (N247)? mem[3772] : 
                        (N249)? mem[3845] : 
                        (N251)? mem[3918] : 
                        (N253)? mem[3991] : 
                        (N255)? mem[4064] : 
                        (N257)? mem[4137] : 
                        (N259)? mem[4210] : 
                        (N261)? mem[4283] : 
                        (N263)? mem[4356] : 
                        (N265)? mem[4429] : 
                        (N267)? mem[4502] : 
                        (N269)? mem[4575] : 
                        (N271)? mem[4648] : 
                        (N146)? mem[4721] : 
                        (N148)? mem[4794] : 
                        (N150)? mem[4867] : 
                        (N152)? mem[4940] : 
                        (N154)? mem[5013] : 
                        (N156)? mem[5086] : 
                        (N158)? mem[5159] : 
                        (N160)? mem[5232] : 
                        (N162)? mem[5305] : 
                        (N164)? mem[5378] : 
                        (N166)? mem[5451] : 
                        (N168)? mem[5524] : 
                        (N170)? mem[5597] : 
                        (N172)? mem[5670] : 
                        (N174)? mem[5743] : 
                        (N176)? mem[5816] : 
                        (N178)? mem[5889] : 
                        (N180)? mem[5962] : 
                        (N182)? mem[6035] : 
                        (N184)? mem[6108] : 
                        (N186)? mem[6181] : 
                        (N188)? mem[6254] : 
                        (N190)? mem[6327] : 
                        (N192)? mem[6400] : 
                        (N194)? mem[6473] : 
                        (N196)? mem[6546] : 
                        (N198)? mem[6619] : 
                        (N200)? mem[6692] : 
                        (N202)? mem[6765] : 
                        (N204)? mem[6838] : 
                        (N206)? mem[6911] : 
                        (N208)? mem[6984] : 
                        (N210)? mem[7057] : 
                        (N212)? mem[7130] : 
                        (N214)? mem[7203] : 
                        (N216)? mem[7276] : 
                        (N218)? mem[7349] : 
                        (N220)? mem[7422] : 
                        (N222)? mem[7495] : 
                        (N224)? mem[7568] : 
                        (N226)? mem[7641] : 
                        (N228)? mem[7714] : 
                        (N230)? mem[7787] : 
                        (N232)? mem[7860] : 
                        (N234)? mem[7933] : 
                        (N236)? mem[8006] : 
                        (N238)? mem[8079] : 
                        (N240)? mem[8152] : 
                        (N242)? mem[8225] : 
                        (N244)? mem[8298] : 
                        (N246)? mem[8371] : 
                        (N248)? mem[8444] : 
                        (N250)? mem[8517] : 
                        (N252)? mem[8590] : 
                        (N254)? mem[8663] : 
                        (N256)? mem[8736] : 
                        (N258)? mem[8809] : 
                        (N260)? mem[8882] : 
                        (N262)? mem[8955] : 
                        (N264)? mem[9028] : 
                        (N266)? mem[9101] : 
                        (N268)? mem[9174] : 
                        (N270)? mem[9247] : 
                        (N272)? mem[9320] : 1'b0;
  assign r_data_o[48] = (N145)? mem[48] : 
                        (N147)? mem[121] : 
                        (N149)? mem[194] : 
                        (N151)? mem[267] : 
                        (N153)? mem[340] : 
                        (N155)? mem[413] : 
                        (N157)? mem[486] : 
                        (N159)? mem[559] : 
                        (N161)? mem[632] : 
                        (N163)? mem[705] : 
                        (N165)? mem[778] : 
                        (N167)? mem[851] : 
                        (N169)? mem[924] : 
                        (N171)? mem[997] : 
                        (N173)? mem[1070] : 
                        (N175)? mem[1143] : 
                        (N177)? mem[1216] : 
                        (N179)? mem[1289] : 
                        (N181)? mem[1362] : 
                        (N183)? mem[1435] : 
                        (N185)? mem[1508] : 
                        (N187)? mem[1581] : 
                        (N189)? mem[1654] : 
                        (N191)? mem[1727] : 
                        (N193)? mem[1800] : 
                        (N195)? mem[1873] : 
                        (N197)? mem[1946] : 
                        (N199)? mem[2019] : 
                        (N201)? mem[2092] : 
                        (N203)? mem[2165] : 
                        (N205)? mem[2238] : 
                        (N207)? mem[2311] : 
                        (N209)? mem[2384] : 
                        (N211)? mem[2457] : 
                        (N213)? mem[2530] : 
                        (N215)? mem[2603] : 
                        (N217)? mem[2676] : 
                        (N219)? mem[2749] : 
                        (N221)? mem[2822] : 
                        (N223)? mem[2895] : 
                        (N225)? mem[2968] : 
                        (N227)? mem[3041] : 
                        (N229)? mem[3114] : 
                        (N231)? mem[3187] : 
                        (N233)? mem[3260] : 
                        (N235)? mem[3333] : 
                        (N237)? mem[3406] : 
                        (N239)? mem[3479] : 
                        (N241)? mem[3552] : 
                        (N243)? mem[3625] : 
                        (N245)? mem[3698] : 
                        (N247)? mem[3771] : 
                        (N249)? mem[3844] : 
                        (N251)? mem[3917] : 
                        (N253)? mem[3990] : 
                        (N255)? mem[4063] : 
                        (N257)? mem[4136] : 
                        (N259)? mem[4209] : 
                        (N261)? mem[4282] : 
                        (N263)? mem[4355] : 
                        (N265)? mem[4428] : 
                        (N267)? mem[4501] : 
                        (N269)? mem[4574] : 
                        (N271)? mem[4647] : 
                        (N146)? mem[4720] : 
                        (N148)? mem[4793] : 
                        (N150)? mem[4866] : 
                        (N152)? mem[4939] : 
                        (N154)? mem[5012] : 
                        (N156)? mem[5085] : 
                        (N158)? mem[5158] : 
                        (N160)? mem[5231] : 
                        (N162)? mem[5304] : 
                        (N164)? mem[5377] : 
                        (N166)? mem[5450] : 
                        (N168)? mem[5523] : 
                        (N170)? mem[5596] : 
                        (N172)? mem[5669] : 
                        (N174)? mem[5742] : 
                        (N176)? mem[5815] : 
                        (N178)? mem[5888] : 
                        (N180)? mem[5961] : 
                        (N182)? mem[6034] : 
                        (N184)? mem[6107] : 
                        (N186)? mem[6180] : 
                        (N188)? mem[6253] : 
                        (N190)? mem[6326] : 
                        (N192)? mem[6399] : 
                        (N194)? mem[6472] : 
                        (N196)? mem[6545] : 
                        (N198)? mem[6618] : 
                        (N200)? mem[6691] : 
                        (N202)? mem[6764] : 
                        (N204)? mem[6837] : 
                        (N206)? mem[6910] : 
                        (N208)? mem[6983] : 
                        (N210)? mem[7056] : 
                        (N212)? mem[7129] : 
                        (N214)? mem[7202] : 
                        (N216)? mem[7275] : 
                        (N218)? mem[7348] : 
                        (N220)? mem[7421] : 
                        (N222)? mem[7494] : 
                        (N224)? mem[7567] : 
                        (N226)? mem[7640] : 
                        (N228)? mem[7713] : 
                        (N230)? mem[7786] : 
                        (N232)? mem[7859] : 
                        (N234)? mem[7932] : 
                        (N236)? mem[8005] : 
                        (N238)? mem[8078] : 
                        (N240)? mem[8151] : 
                        (N242)? mem[8224] : 
                        (N244)? mem[8297] : 
                        (N246)? mem[8370] : 
                        (N248)? mem[8443] : 
                        (N250)? mem[8516] : 
                        (N252)? mem[8589] : 
                        (N254)? mem[8662] : 
                        (N256)? mem[8735] : 
                        (N258)? mem[8808] : 
                        (N260)? mem[8881] : 
                        (N262)? mem[8954] : 
                        (N264)? mem[9027] : 
                        (N266)? mem[9100] : 
                        (N268)? mem[9173] : 
                        (N270)? mem[9246] : 
                        (N272)? mem[9319] : 1'b0;
  assign r_data_o[47] = (N145)? mem[47] : 
                        (N147)? mem[120] : 
                        (N149)? mem[193] : 
                        (N151)? mem[266] : 
                        (N153)? mem[339] : 
                        (N155)? mem[412] : 
                        (N157)? mem[485] : 
                        (N159)? mem[558] : 
                        (N161)? mem[631] : 
                        (N163)? mem[704] : 
                        (N165)? mem[777] : 
                        (N167)? mem[850] : 
                        (N169)? mem[923] : 
                        (N171)? mem[996] : 
                        (N173)? mem[1069] : 
                        (N175)? mem[1142] : 
                        (N177)? mem[1215] : 
                        (N179)? mem[1288] : 
                        (N181)? mem[1361] : 
                        (N183)? mem[1434] : 
                        (N185)? mem[1507] : 
                        (N187)? mem[1580] : 
                        (N189)? mem[1653] : 
                        (N191)? mem[1726] : 
                        (N193)? mem[1799] : 
                        (N195)? mem[1872] : 
                        (N197)? mem[1945] : 
                        (N199)? mem[2018] : 
                        (N201)? mem[2091] : 
                        (N203)? mem[2164] : 
                        (N205)? mem[2237] : 
                        (N207)? mem[2310] : 
                        (N209)? mem[2383] : 
                        (N211)? mem[2456] : 
                        (N213)? mem[2529] : 
                        (N215)? mem[2602] : 
                        (N217)? mem[2675] : 
                        (N219)? mem[2748] : 
                        (N221)? mem[2821] : 
                        (N223)? mem[2894] : 
                        (N225)? mem[2967] : 
                        (N227)? mem[3040] : 
                        (N229)? mem[3113] : 
                        (N231)? mem[3186] : 
                        (N233)? mem[3259] : 
                        (N235)? mem[3332] : 
                        (N237)? mem[3405] : 
                        (N239)? mem[3478] : 
                        (N241)? mem[3551] : 
                        (N243)? mem[3624] : 
                        (N245)? mem[3697] : 
                        (N247)? mem[3770] : 
                        (N249)? mem[3843] : 
                        (N251)? mem[3916] : 
                        (N253)? mem[3989] : 
                        (N255)? mem[4062] : 
                        (N257)? mem[4135] : 
                        (N259)? mem[4208] : 
                        (N261)? mem[4281] : 
                        (N263)? mem[4354] : 
                        (N265)? mem[4427] : 
                        (N267)? mem[4500] : 
                        (N269)? mem[4573] : 
                        (N271)? mem[4646] : 
                        (N146)? mem[4719] : 
                        (N148)? mem[4792] : 
                        (N150)? mem[4865] : 
                        (N152)? mem[4938] : 
                        (N154)? mem[5011] : 
                        (N156)? mem[5084] : 
                        (N158)? mem[5157] : 
                        (N160)? mem[5230] : 
                        (N162)? mem[5303] : 
                        (N164)? mem[5376] : 
                        (N166)? mem[5449] : 
                        (N168)? mem[5522] : 
                        (N170)? mem[5595] : 
                        (N172)? mem[5668] : 
                        (N174)? mem[5741] : 
                        (N176)? mem[5814] : 
                        (N178)? mem[5887] : 
                        (N180)? mem[5960] : 
                        (N182)? mem[6033] : 
                        (N184)? mem[6106] : 
                        (N186)? mem[6179] : 
                        (N188)? mem[6252] : 
                        (N190)? mem[6325] : 
                        (N192)? mem[6398] : 
                        (N194)? mem[6471] : 
                        (N196)? mem[6544] : 
                        (N198)? mem[6617] : 
                        (N200)? mem[6690] : 
                        (N202)? mem[6763] : 
                        (N204)? mem[6836] : 
                        (N206)? mem[6909] : 
                        (N208)? mem[6982] : 
                        (N210)? mem[7055] : 
                        (N212)? mem[7128] : 
                        (N214)? mem[7201] : 
                        (N216)? mem[7274] : 
                        (N218)? mem[7347] : 
                        (N220)? mem[7420] : 
                        (N222)? mem[7493] : 
                        (N224)? mem[7566] : 
                        (N226)? mem[7639] : 
                        (N228)? mem[7712] : 
                        (N230)? mem[7785] : 
                        (N232)? mem[7858] : 
                        (N234)? mem[7931] : 
                        (N236)? mem[8004] : 
                        (N238)? mem[8077] : 
                        (N240)? mem[8150] : 
                        (N242)? mem[8223] : 
                        (N244)? mem[8296] : 
                        (N246)? mem[8369] : 
                        (N248)? mem[8442] : 
                        (N250)? mem[8515] : 
                        (N252)? mem[8588] : 
                        (N254)? mem[8661] : 
                        (N256)? mem[8734] : 
                        (N258)? mem[8807] : 
                        (N260)? mem[8880] : 
                        (N262)? mem[8953] : 
                        (N264)? mem[9026] : 
                        (N266)? mem[9099] : 
                        (N268)? mem[9172] : 
                        (N270)? mem[9245] : 
                        (N272)? mem[9318] : 1'b0;
  assign r_data_o[46] = (N145)? mem[46] : 
                        (N147)? mem[119] : 
                        (N149)? mem[192] : 
                        (N151)? mem[265] : 
                        (N153)? mem[338] : 
                        (N155)? mem[411] : 
                        (N157)? mem[484] : 
                        (N159)? mem[557] : 
                        (N161)? mem[630] : 
                        (N163)? mem[703] : 
                        (N165)? mem[776] : 
                        (N167)? mem[849] : 
                        (N169)? mem[922] : 
                        (N171)? mem[995] : 
                        (N173)? mem[1068] : 
                        (N175)? mem[1141] : 
                        (N177)? mem[1214] : 
                        (N179)? mem[1287] : 
                        (N181)? mem[1360] : 
                        (N183)? mem[1433] : 
                        (N185)? mem[1506] : 
                        (N187)? mem[1579] : 
                        (N189)? mem[1652] : 
                        (N191)? mem[1725] : 
                        (N193)? mem[1798] : 
                        (N195)? mem[1871] : 
                        (N197)? mem[1944] : 
                        (N199)? mem[2017] : 
                        (N201)? mem[2090] : 
                        (N203)? mem[2163] : 
                        (N205)? mem[2236] : 
                        (N207)? mem[2309] : 
                        (N209)? mem[2382] : 
                        (N211)? mem[2455] : 
                        (N213)? mem[2528] : 
                        (N215)? mem[2601] : 
                        (N217)? mem[2674] : 
                        (N219)? mem[2747] : 
                        (N221)? mem[2820] : 
                        (N223)? mem[2893] : 
                        (N225)? mem[2966] : 
                        (N227)? mem[3039] : 
                        (N229)? mem[3112] : 
                        (N231)? mem[3185] : 
                        (N233)? mem[3258] : 
                        (N235)? mem[3331] : 
                        (N237)? mem[3404] : 
                        (N239)? mem[3477] : 
                        (N241)? mem[3550] : 
                        (N243)? mem[3623] : 
                        (N245)? mem[3696] : 
                        (N247)? mem[3769] : 
                        (N249)? mem[3842] : 
                        (N251)? mem[3915] : 
                        (N253)? mem[3988] : 
                        (N255)? mem[4061] : 
                        (N257)? mem[4134] : 
                        (N259)? mem[4207] : 
                        (N261)? mem[4280] : 
                        (N263)? mem[4353] : 
                        (N265)? mem[4426] : 
                        (N267)? mem[4499] : 
                        (N269)? mem[4572] : 
                        (N271)? mem[4645] : 
                        (N146)? mem[4718] : 
                        (N148)? mem[4791] : 
                        (N150)? mem[4864] : 
                        (N152)? mem[4937] : 
                        (N154)? mem[5010] : 
                        (N156)? mem[5083] : 
                        (N158)? mem[5156] : 
                        (N160)? mem[5229] : 
                        (N162)? mem[5302] : 
                        (N164)? mem[5375] : 
                        (N166)? mem[5448] : 
                        (N168)? mem[5521] : 
                        (N170)? mem[5594] : 
                        (N172)? mem[5667] : 
                        (N174)? mem[5740] : 
                        (N176)? mem[5813] : 
                        (N178)? mem[5886] : 
                        (N180)? mem[5959] : 
                        (N182)? mem[6032] : 
                        (N184)? mem[6105] : 
                        (N186)? mem[6178] : 
                        (N188)? mem[6251] : 
                        (N190)? mem[6324] : 
                        (N192)? mem[6397] : 
                        (N194)? mem[6470] : 
                        (N196)? mem[6543] : 
                        (N198)? mem[6616] : 
                        (N200)? mem[6689] : 
                        (N202)? mem[6762] : 
                        (N204)? mem[6835] : 
                        (N206)? mem[6908] : 
                        (N208)? mem[6981] : 
                        (N210)? mem[7054] : 
                        (N212)? mem[7127] : 
                        (N214)? mem[7200] : 
                        (N216)? mem[7273] : 
                        (N218)? mem[7346] : 
                        (N220)? mem[7419] : 
                        (N222)? mem[7492] : 
                        (N224)? mem[7565] : 
                        (N226)? mem[7638] : 
                        (N228)? mem[7711] : 
                        (N230)? mem[7784] : 
                        (N232)? mem[7857] : 
                        (N234)? mem[7930] : 
                        (N236)? mem[8003] : 
                        (N238)? mem[8076] : 
                        (N240)? mem[8149] : 
                        (N242)? mem[8222] : 
                        (N244)? mem[8295] : 
                        (N246)? mem[8368] : 
                        (N248)? mem[8441] : 
                        (N250)? mem[8514] : 
                        (N252)? mem[8587] : 
                        (N254)? mem[8660] : 
                        (N256)? mem[8733] : 
                        (N258)? mem[8806] : 
                        (N260)? mem[8879] : 
                        (N262)? mem[8952] : 
                        (N264)? mem[9025] : 
                        (N266)? mem[9098] : 
                        (N268)? mem[9171] : 
                        (N270)? mem[9244] : 
                        (N272)? mem[9317] : 1'b0;
  assign r_data_o[45] = (N145)? mem[45] : 
                        (N147)? mem[118] : 
                        (N149)? mem[191] : 
                        (N151)? mem[264] : 
                        (N153)? mem[337] : 
                        (N155)? mem[410] : 
                        (N157)? mem[483] : 
                        (N159)? mem[556] : 
                        (N161)? mem[629] : 
                        (N163)? mem[702] : 
                        (N165)? mem[775] : 
                        (N167)? mem[848] : 
                        (N169)? mem[921] : 
                        (N171)? mem[994] : 
                        (N173)? mem[1067] : 
                        (N175)? mem[1140] : 
                        (N177)? mem[1213] : 
                        (N179)? mem[1286] : 
                        (N181)? mem[1359] : 
                        (N183)? mem[1432] : 
                        (N185)? mem[1505] : 
                        (N187)? mem[1578] : 
                        (N189)? mem[1651] : 
                        (N191)? mem[1724] : 
                        (N193)? mem[1797] : 
                        (N195)? mem[1870] : 
                        (N197)? mem[1943] : 
                        (N199)? mem[2016] : 
                        (N201)? mem[2089] : 
                        (N203)? mem[2162] : 
                        (N205)? mem[2235] : 
                        (N207)? mem[2308] : 
                        (N209)? mem[2381] : 
                        (N211)? mem[2454] : 
                        (N213)? mem[2527] : 
                        (N215)? mem[2600] : 
                        (N217)? mem[2673] : 
                        (N219)? mem[2746] : 
                        (N221)? mem[2819] : 
                        (N223)? mem[2892] : 
                        (N225)? mem[2965] : 
                        (N227)? mem[3038] : 
                        (N229)? mem[3111] : 
                        (N231)? mem[3184] : 
                        (N233)? mem[3257] : 
                        (N235)? mem[3330] : 
                        (N237)? mem[3403] : 
                        (N239)? mem[3476] : 
                        (N241)? mem[3549] : 
                        (N243)? mem[3622] : 
                        (N245)? mem[3695] : 
                        (N247)? mem[3768] : 
                        (N249)? mem[3841] : 
                        (N251)? mem[3914] : 
                        (N253)? mem[3987] : 
                        (N255)? mem[4060] : 
                        (N257)? mem[4133] : 
                        (N259)? mem[4206] : 
                        (N261)? mem[4279] : 
                        (N263)? mem[4352] : 
                        (N265)? mem[4425] : 
                        (N267)? mem[4498] : 
                        (N269)? mem[4571] : 
                        (N271)? mem[4644] : 
                        (N146)? mem[4717] : 
                        (N148)? mem[4790] : 
                        (N150)? mem[4863] : 
                        (N152)? mem[4936] : 
                        (N154)? mem[5009] : 
                        (N156)? mem[5082] : 
                        (N158)? mem[5155] : 
                        (N160)? mem[5228] : 
                        (N162)? mem[5301] : 
                        (N164)? mem[5374] : 
                        (N166)? mem[5447] : 
                        (N168)? mem[5520] : 
                        (N170)? mem[5593] : 
                        (N172)? mem[5666] : 
                        (N174)? mem[5739] : 
                        (N176)? mem[5812] : 
                        (N178)? mem[5885] : 
                        (N180)? mem[5958] : 
                        (N182)? mem[6031] : 
                        (N184)? mem[6104] : 
                        (N186)? mem[6177] : 
                        (N188)? mem[6250] : 
                        (N190)? mem[6323] : 
                        (N192)? mem[6396] : 
                        (N194)? mem[6469] : 
                        (N196)? mem[6542] : 
                        (N198)? mem[6615] : 
                        (N200)? mem[6688] : 
                        (N202)? mem[6761] : 
                        (N204)? mem[6834] : 
                        (N206)? mem[6907] : 
                        (N208)? mem[6980] : 
                        (N210)? mem[7053] : 
                        (N212)? mem[7126] : 
                        (N214)? mem[7199] : 
                        (N216)? mem[7272] : 
                        (N218)? mem[7345] : 
                        (N220)? mem[7418] : 
                        (N222)? mem[7491] : 
                        (N224)? mem[7564] : 
                        (N226)? mem[7637] : 
                        (N228)? mem[7710] : 
                        (N230)? mem[7783] : 
                        (N232)? mem[7856] : 
                        (N234)? mem[7929] : 
                        (N236)? mem[8002] : 
                        (N238)? mem[8075] : 
                        (N240)? mem[8148] : 
                        (N242)? mem[8221] : 
                        (N244)? mem[8294] : 
                        (N246)? mem[8367] : 
                        (N248)? mem[8440] : 
                        (N250)? mem[8513] : 
                        (N252)? mem[8586] : 
                        (N254)? mem[8659] : 
                        (N256)? mem[8732] : 
                        (N258)? mem[8805] : 
                        (N260)? mem[8878] : 
                        (N262)? mem[8951] : 
                        (N264)? mem[9024] : 
                        (N266)? mem[9097] : 
                        (N268)? mem[9170] : 
                        (N270)? mem[9243] : 
                        (N272)? mem[9316] : 1'b0;
  assign r_data_o[44] = (N145)? mem[44] : 
                        (N147)? mem[117] : 
                        (N149)? mem[190] : 
                        (N151)? mem[263] : 
                        (N153)? mem[336] : 
                        (N155)? mem[409] : 
                        (N157)? mem[482] : 
                        (N159)? mem[555] : 
                        (N161)? mem[628] : 
                        (N163)? mem[701] : 
                        (N165)? mem[774] : 
                        (N167)? mem[847] : 
                        (N169)? mem[920] : 
                        (N171)? mem[993] : 
                        (N173)? mem[1066] : 
                        (N175)? mem[1139] : 
                        (N177)? mem[1212] : 
                        (N179)? mem[1285] : 
                        (N181)? mem[1358] : 
                        (N183)? mem[1431] : 
                        (N185)? mem[1504] : 
                        (N187)? mem[1577] : 
                        (N189)? mem[1650] : 
                        (N191)? mem[1723] : 
                        (N193)? mem[1796] : 
                        (N195)? mem[1869] : 
                        (N197)? mem[1942] : 
                        (N199)? mem[2015] : 
                        (N201)? mem[2088] : 
                        (N203)? mem[2161] : 
                        (N205)? mem[2234] : 
                        (N207)? mem[2307] : 
                        (N209)? mem[2380] : 
                        (N211)? mem[2453] : 
                        (N213)? mem[2526] : 
                        (N215)? mem[2599] : 
                        (N217)? mem[2672] : 
                        (N219)? mem[2745] : 
                        (N221)? mem[2818] : 
                        (N223)? mem[2891] : 
                        (N225)? mem[2964] : 
                        (N227)? mem[3037] : 
                        (N229)? mem[3110] : 
                        (N231)? mem[3183] : 
                        (N233)? mem[3256] : 
                        (N235)? mem[3329] : 
                        (N237)? mem[3402] : 
                        (N239)? mem[3475] : 
                        (N241)? mem[3548] : 
                        (N243)? mem[3621] : 
                        (N245)? mem[3694] : 
                        (N247)? mem[3767] : 
                        (N249)? mem[3840] : 
                        (N251)? mem[3913] : 
                        (N253)? mem[3986] : 
                        (N255)? mem[4059] : 
                        (N257)? mem[4132] : 
                        (N259)? mem[4205] : 
                        (N261)? mem[4278] : 
                        (N263)? mem[4351] : 
                        (N265)? mem[4424] : 
                        (N267)? mem[4497] : 
                        (N269)? mem[4570] : 
                        (N271)? mem[4643] : 
                        (N146)? mem[4716] : 
                        (N148)? mem[4789] : 
                        (N150)? mem[4862] : 
                        (N152)? mem[4935] : 
                        (N154)? mem[5008] : 
                        (N156)? mem[5081] : 
                        (N158)? mem[5154] : 
                        (N160)? mem[5227] : 
                        (N162)? mem[5300] : 
                        (N164)? mem[5373] : 
                        (N166)? mem[5446] : 
                        (N168)? mem[5519] : 
                        (N170)? mem[5592] : 
                        (N172)? mem[5665] : 
                        (N174)? mem[5738] : 
                        (N176)? mem[5811] : 
                        (N178)? mem[5884] : 
                        (N180)? mem[5957] : 
                        (N182)? mem[6030] : 
                        (N184)? mem[6103] : 
                        (N186)? mem[6176] : 
                        (N188)? mem[6249] : 
                        (N190)? mem[6322] : 
                        (N192)? mem[6395] : 
                        (N194)? mem[6468] : 
                        (N196)? mem[6541] : 
                        (N198)? mem[6614] : 
                        (N200)? mem[6687] : 
                        (N202)? mem[6760] : 
                        (N204)? mem[6833] : 
                        (N206)? mem[6906] : 
                        (N208)? mem[6979] : 
                        (N210)? mem[7052] : 
                        (N212)? mem[7125] : 
                        (N214)? mem[7198] : 
                        (N216)? mem[7271] : 
                        (N218)? mem[7344] : 
                        (N220)? mem[7417] : 
                        (N222)? mem[7490] : 
                        (N224)? mem[7563] : 
                        (N226)? mem[7636] : 
                        (N228)? mem[7709] : 
                        (N230)? mem[7782] : 
                        (N232)? mem[7855] : 
                        (N234)? mem[7928] : 
                        (N236)? mem[8001] : 
                        (N238)? mem[8074] : 
                        (N240)? mem[8147] : 
                        (N242)? mem[8220] : 
                        (N244)? mem[8293] : 
                        (N246)? mem[8366] : 
                        (N248)? mem[8439] : 
                        (N250)? mem[8512] : 
                        (N252)? mem[8585] : 
                        (N254)? mem[8658] : 
                        (N256)? mem[8731] : 
                        (N258)? mem[8804] : 
                        (N260)? mem[8877] : 
                        (N262)? mem[8950] : 
                        (N264)? mem[9023] : 
                        (N266)? mem[9096] : 
                        (N268)? mem[9169] : 
                        (N270)? mem[9242] : 
                        (N272)? mem[9315] : 1'b0;
  assign r_data_o[43] = (N145)? mem[43] : 
                        (N147)? mem[116] : 
                        (N149)? mem[189] : 
                        (N151)? mem[262] : 
                        (N153)? mem[335] : 
                        (N155)? mem[408] : 
                        (N157)? mem[481] : 
                        (N159)? mem[554] : 
                        (N161)? mem[627] : 
                        (N163)? mem[700] : 
                        (N165)? mem[773] : 
                        (N167)? mem[846] : 
                        (N169)? mem[919] : 
                        (N171)? mem[992] : 
                        (N173)? mem[1065] : 
                        (N175)? mem[1138] : 
                        (N177)? mem[1211] : 
                        (N179)? mem[1284] : 
                        (N181)? mem[1357] : 
                        (N183)? mem[1430] : 
                        (N185)? mem[1503] : 
                        (N187)? mem[1576] : 
                        (N189)? mem[1649] : 
                        (N191)? mem[1722] : 
                        (N193)? mem[1795] : 
                        (N195)? mem[1868] : 
                        (N197)? mem[1941] : 
                        (N199)? mem[2014] : 
                        (N201)? mem[2087] : 
                        (N203)? mem[2160] : 
                        (N205)? mem[2233] : 
                        (N207)? mem[2306] : 
                        (N209)? mem[2379] : 
                        (N211)? mem[2452] : 
                        (N213)? mem[2525] : 
                        (N215)? mem[2598] : 
                        (N217)? mem[2671] : 
                        (N219)? mem[2744] : 
                        (N221)? mem[2817] : 
                        (N223)? mem[2890] : 
                        (N225)? mem[2963] : 
                        (N227)? mem[3036] : 
                        (N229)? mem[3109] : 
                        (N231)? mem[3182] : 
                        (N233)? mem[3255] : 
                        (N235)? mem[3328] : 
                        (N237)? mem[3401] : 
                        (N239)? mem[3474] : 
                        (N241)? mem[3547] : 
                        (N243)? mem[3620] : 
                        (N245)? mem[3693] : 
                        (N247)? mem[3766] : 
                        (N249)? mem[3839] : 
                        (N251)? mem[3912] : 
                        (N253)? mem[3985] : 
                        (N255)? mem[4058] : 
                        (N257)? mem[4131] : 
                        (N259)? mem[4204] : 
                        (N261)? mem[4277] : 
                        (N263)? mem[4350] : 
                        (N265)? mem[4423] : 
                        (N267)? mem[4496] : 
                        (N269)? mem[4569] : 
                        (N271)? mem[4642] : 
                        (N146)? mem[4715] : 
                        (N148)? mem[4788] : 
                        (N150)? mem[4861] : 
                        (N152)? mem[4934] : 
                        (N154)? mem[5007] : 
                        (N156)? mem[5080] : 
                        (N158)? mem[5153] : 
                        (N160)? mem[5226] : 
                        (N162)? mem[5299] : 
                        (N164)? mem[5372] : 
                        (N166)? mem[5445] : 
                        (N168)? mem[5518] : 
                        (N170)? mem[5591] : 
                        (N172)? mem[5664] : 
                        (N174)? mem[5737] : 
                        (N176)? mem[5810] : 
                        (N178)? mem[5883] : 
                        (N180)? mem[5956] : 
                        (N182)? mem[6029] : 
                        (N184)? mem[6102] : 
                        (N186)? mem[6175] : 
                        (N188)? mem[6248] : 
                        (N190)? mem[6321] : 
                        (N192)? mem[6394] : 
                        (N194)? mem[6467] : 
                        (N196)? mem[6540] : 
                        (N198)? mem[6613] : 
                        (N200)? mem[6686] : 
                        (N202)? mem[6759] : 
                        (N204)? mem[6832] : 
                        (N206)? mem[6905] : 
                        (N208)? mem[6978] : 
                        (N210)? mem[7051] : 
                        (N212)? mem[7124] : 
                        (N214)? mem[7197] : 
                        (N216)? mem[7270] : 
                        (N218)? mem[7343] : 
                        (N220)? mem[7416] : 
                        (N222)? mem[7489] : 
                        (N224)? mem[7562] : 
                        (N226)? mem[7635] : 
                        (N228)? mem[7708] : 
                        (N230)? mem[7781] : 
                        (N232)? mem[7854] : 
                        (N234)? mem[7927] : 
                        (N236)? mem[8000] : 
                        (N238)? mem[8073] : 
                        (N240)? mem[8146] : 
                        (N242)? mem[8219] : 
                        (N244)? mem[8292] : 
                        (N246)? mem[8365] : 
                        (N248)? mem[8438] : 
                        (N250)? mem[8511] : 
                        (N252)? mem[8584] : 
                        (N254)? mem[8657] : 
                        (N256)? mem[8730] : 
                        (N258)? mem[8803] : 
                        (N260)? mem[8876] : 
                        (N262)? mem[8949] : 
                        (N264)? mem[9022] : 
                        (N266)? mem[9095] : 
                        (N268)? mem[9168] : 
                        (N270)? mem[9241] : 
                        (N272)? mem[9314] : 1'b0;
  assign r_data_o[42] = (N145)? mem[42] : 
                        (N147)? mem[115] : 
                        (N149)? mem[188] : 
                        (N151)? mem[261] : 
                        (N153)? mem[334] : 
                        (N155)? mem[407] : 
                        (N157)? mem[480] : 
                        (N159)? mem[553] : 
                        (N161)? mem[626] : 
                        (N163)? mem[699] : 
                        (N165)? mem[772] : 
                        (N167)? mem[845] : 
                        (N169)? mem[918] : 
                        (N171)? mem[991] : 
                        (N173)? mem[1064] : 
                        (N175)? mem[1137] : 
                        (N177)? mem[1210] : 
                        (N179)? mem[1283] : 
                        (N181)? mem[1356] : 
                        (N183)? mem[1429] : 
                        (N185)? mem[1502] : 
                        (N187)? mem[1575] : 
                        (N189)? mem[1648] : 
                        (N191)? mem[1721] : 
                        (N193)? mem[1794] : 
                        (N195)? mem[1867] : 
                        (N197)? mem[1940] : 
                        (N199)? mem[2013] : 
                        (N201)? mem[2086] : 
                        (N203)? mem[2159] : 
                        (N205)? mem[2232] : 
                        (N207)? mem[2305] : 
                        (N209)? mem[2378] : 
                        (N211)? mem[2451] : 
                        (N213)? mem[2524] : 
                        (N215)? mem[2597] : 
                        (N217)? mem[2670] : 
                        (N219)? mem[2743] : 
                        (N221)? mem[2816] : 
                        (N223)? mem[2889] : 
                        (N225)? mem[2962] : 
                        (N227)? mem[3035] : 
                        (N229)? mem[3108] : 
                        (N231)? mem[3181] : 
                        (N233)? mem[3254] : 
                        (N235)? mem[3327] : 
                        (N237)? mem[3400] : 
                        (N239)? mem[3473] : 
                        (N241)? mem[3546] : 
                        (N243)? mem[3619] : 
                        (N245)? mem[3692] : 
                        (N247)? mem[3765] : 
                        (N249)? mem[3838] : 
                        (N251)? mem[3911] : 
                        (N253)? mem[3984] : 
                        (N255)? mem[4057] : 
                        (N257)? mem[4130] : 
                        (N259)? mem[4203] : 
                        (N261)? mem[4276] : 
                        (N263)? mem[4349] : 
                        (N265)? mem[4422] : 
                        (N267)? mem[4495] : 
                        (N269)? mem[4568] : 
                        (N271)? mem[4641] : 
                        (N146)? mem[4714] : 
                        (N148)? mem[4787] : 
                        (N150)? mem[4860] : 
                        (N152)? mem[4933] : 
                        (N154)? mem[5006] : 
                        (N156)? mem[5079] : 
                        (N158)? mem[5152] : 
                        (N160)? mem[5225] : 
                        (N162)? mem[5298] : 
                        (N164)? mem[5371] : 
                        (N166)? mem[5444] : 
                        (N168)? mem[5517] : 
                        (N170)? mem[5590] : 
                        (N172)? mem[5663] : 
                        (N174)? mem[5736] : 
                        (N176)? mem[5809] : 
                        (N178)? mem[5882] : 
                        (N180)? mem[5955] : 
                        (N182)? mem[6028] : 
                        (N184)? mem[6101] : 
                        (N186)? mem[6174] : 
                        (N188)? mem[6247] : 
                        (N190)? mem[6320] : 
                        (N192)? mem[6393] : 
                        (N194)? mem[6466] : 
                        (N196)? mem[6539] : 
                        (N198)? mem[6612] : 
                        (N200)? mem[6685] : 
                        (N202)? mem[6758] : 
                        (N204)? mem[6831] : 
                        (N206)? mem[6904] : 
                        (N208)? mem[6977] : 
                        (N210)? mem[7050] : 
                        (N212)? mem[7123] : 
                        (N214)? mem[7196] : 
                        (N216)? mem[7269] : 
                        (N218)? mem[7342] : 
                        (N220)? mem[7415] : 
                        (N222)? mem[7488] : 
                        (N224)? mem[7561] : 
                        (N226)? mem[7634] : 
                        (N228)? mem[7707] : 
                        (N230)? mem[7780] : 
                        (N232)? mem[7853] : 
                        (N234)? mem[7926] : 
                        (N236)? mem[7999] : 
                        (N238)? mem[8072] : 
                        (N240)? mem[8145] : 
                        (N242)? mem[8218] : 
                        (N244)? mem[8291] : 
                        (N246)? mem[8364] : 
                        (N248)? mem[8437] : 
                        (N250)? mem[8510] : 
                        (N252)? mem[8583] : 
                        (N254)? mem[8656] : 
                        (N256)? mem[8729] : 
                        (N258)? mem[8802] : 
                        (N260)? mem[8875] : 
                        (N262)? mem[8948] : 
                        (N264)? mem[9021] : 
                        (N266)? mem[9094] : 
                        (N268)? mem[9167] : 
                        (N270)? mem[9240] : 
                        (N272)? mem[9313] : 1'b0;
  assign r_data_o[41] = (N145)? mem[41] : 
                        (N147)? mem[114] : 
                        (N149)? mem[187] : 
                        (N151)? mem[260] : 
                        (N153)? mem[333] : 
                        (N155)? mem[406] : 
                        (N157)? mem[479] : 
                        (N159)? mem[552] : 
                        (N161)? mem[625] : 
                        (N163)? mem[698] : 
                        (N165)? mem[771] : 
                        (N167)? mem[844] : 
                        (N169)? mem[917] : 
                        (N171)? mem[990] : 
                        (N173)? mem[1063] : 
                        (N175)? mem[1136] : 
                        (N177)? mem[1209] : 
                        (N179)? mem[1282] : 
                        (N181)? mem[1355] : 
                        (N183)? mem[1428] : 
                        (N185)? mem[1501] : 
                        (N187)? mem[1574] : 
                        (N189)? mem[1647] : 
                        (N191)? mem[1720] : 
                        (N193)? mem[1793] : 
                        (N195)? mem[1866] : 
                        (N197)? mem[1939] : 
                        (N199)? mem[2012] : 
                        (N201)? mem[2085] : 
                        (N203)? mem[2158] : 
                        (N205)? mem[2231] : 
                        (N207)? mem[2304] : 
                        (N209)? mem[2377] : 
                        (N211)? mem[2450] : 
                        (N213)? mem[2523] : 
                        (N215)? mem[2596] : 
                        (N217)? mem[2669] : 
                        (N219)? mem[2742] : 
                        (N221)? mem[2815] : 
                        (N223)? mem[2888] : 
                        (N225)? mem[2961] : 
                        (N227)? mem[3034] : 
                        (N229)? mem[3107] : 
                        (N231)? mem[3180] : 
                        (N233)? mem[3253] : 
                        (N235)? mem[3326] : 
                        (N237)? mem[3399] : 
                        (N239)? mem[3472] : 
                        (N241)? mem[3545] : 
                        (N243)? mem[3618] : 
                        (N245)? mem[3691] : 
                        (N247)? mem[3764] : 
                        (N249)? mem[3837] : 
                        (N251)? mem[3910] : 
                        (N253)? mem[3983] : 
                        (N255)? mem[4056] : 
                        (N257)? mem[4129] : 
                        (N259)? mem[4202] : 
                        (N261)? mem[4275] : 
                        (N263)? mem[4348] : 
                        (N265)? mem[4421] : 
                        (N267)? mem[4494] : 
                        (N269)? mem[4567] : 
                        (N271)? mem[4640] : 
                        (N146)? mem[4713] : 
                        (N148)? mem[4786] : 
                        (N150)? mem[4859] : 
                        (N152)? mem[4932] : 
                        (N154)? mem[5005] : 
                        (N156)? mem[5078] : 
                        (N158)? mem[5151] : 
                        (N160)? mem[5224] : 
                        (N162)? mem[5297] : 
                        (N164)? mem[5370] : 
                        (N166)? mem[5443] : 
                        (N168)? mem[5516] : 
                        (N170)? mem[5589] : 
                        (N172)? mem[5662] : 
                        (N174)? mem[5735] : 
                        (N176)? mem[5808] : 
                        (N178)? mem[5881] : 
                        (N180)? mem[5954] : 
                        (N182)? mem[6027] : 
                        (N184)? mem[6100] : 
                        (N186)? mem[6173] : 
                        (N188)? mem[6246] : 
                        (N190)? mem[6319] : 
                        (N192)? mem[6392] : 
                        (N194)? mem[6465] : 
                        (N196)? mem[6538] : 
                        (N198)? mem[6611] : 
                        (N200)? mem[6684] : 
                        (N202)? mem[6757] : 
                        (N204)? mem[6830] : 
                        (N206)? mem[6903] : 
                        (N208)? mem[6976] : 
                        (N210)? mem[7049] : 
                        (N212)? mem[7122] : 
                        (N214)? mem[7195] : 
                        (N216)? mem[7268] : 
                        (N218)? mem[7341] : 
                        (N220)? mem[7414] : 
                        (N222)? mem[7487] : 
                        (N224)? mem[7560] : 
                        (N226)? mem[7633] : 
                        (N228)? mem[7706] : 
                        (N230)? mem[7779] : 
                        (N232)? mem[7852] : 
                        (N234)? mem[7925] : 
                        (N236)? mem[7998] : 
                        (N238)? mem[8071] : 
                        (N240)? mem[8144] : 
                        (N242)? mem[8217] : 
                        (N244)? mem[8290] : 
                        (N246)? mem[8363] : 
                        (N248)? mem[8436] : 
                        (N250)? mem[8509] : 
                        (N252)? mem[8582] : 
                        (N254)? mem[8655] : 
                        (N256)? mem[8728] : 
                        (N258)? mem[8801] : 
                        (N260)? mem[8874] : 
                        (N262)? mem[8947] : 
                        (N264)? mem[9020] : 
                        (N266)? mem[9093] : 
                        (N268)? mem[9166] : 
                        (N270)? mem[9239] : 
                        (N272)? mem[9312] : 1'b0;
  assign r_data_o[40] = (N145)? mem[40] : 
                        (N147)? mem[113] : 
                        (N149)? mem[186] : 
                        (N151)? mem[259] : 
                        (N153)? mem[332] : 
                        (N155)? mem[405] : 
                        (N157)? mem[478] : 
                        (N159)? mem[551] : 
                        (N161)? mem[624] : 
                        (N163)? mem[697] : 
                        (N165)? mem[770] : 
                        (N167)? mem[843] : 
                        (N169)? mem[916] : 
                        (N171)? mem[989] : 
                        (N173)? mem[1062] : 
                        (N175)? mem[1135] : 
                        (N177)? mem[1208] : 
                        (N179)? mem[1281] : 
                        (N181)? mem[1354] : 
                        (N183)? mem[1427] : 
                        (N185)? mem[1500] : 
                        (N187)? mem[1573] : 
                        (N189)? mem[1646] : 
                        (N191)? mem[1719] : 
                        (N193)? mem[1792] : 
                        (N195)? mem[1865] : 
                        (N197)? mem[1938] : 
                        (N199)? mem[2011] : 
                        (N201)? mem[2084] : 
                        (N203)? mem[2157] : 
                        (N205)? mem[2230] : 
                        (N207)? mem[2303] : 
                        (N209)? mem[2376] : 
                        (N211)? mem[2449] : 
                        (N213)? mem[2522] : 
                        (N215)? mem[2595] : 
                        (N217)? mem[2668] : 
                        (N219)? mem[2741] : 
                        (N221)? mem[2814] : 
                        (N223)? mem[2887] : 
                        (N225)? mem[2960] : 
                        (N227)? mem[3033] : 
                        (N229)? mem[3106] : 
                        (N231)? mem[3179] : 
                        (N233)? mem[3252] : 
                        (N235)? mem[3325] : 
                        (N237)? mem[3398] : 
                        (N239)? mem[3471] : 
                        (N241)? mem[3544] : 
                        (N243)? mem[3617] : 
                        (N245)? mem[3690] : 
                        (N247)? mem[3763] : 
                        (N249)? mem[3836] : 
                        (N251)? mem[3909] : 
                        (N253)? mem[3982] : 
                        (N255)? mem[4055] : 
                        (N257)? mem[4128] : 
                        (N259)? mem[4201] : 
                        (N261)? mem[4274] : 
                        (N263)? mem[4347] : 
                        (N265)? mem[4420] : 
                        (N267)? mem[4493] : 
                        (N269)? mem[4566] : 
                        (N271)? mem[4639] : 
                        (N146)? mem[4712] : 
                        (N148)? mem[4785] : 
                        (N150)? mem[4858] : 
                        (N152)? mem[4931] : 
                        (N154)? mem[5004] : 
                        (N156)? mem[5077] : 
                        (N158)? mem[5150] : 
                        (N160)? mem[5223] : 
                        (N162)? mem[5296] : 
                        (N164)? mem[5369] : 
                        (N166)? mem[5442] : 
                        (N168)? mem[5515] : 
                        (N170)? mem[5588] : 
                        (N172)? mem[5661] : 
                        (N174)? mem[5734] : 
                        (N176)? mem[5807] : 
                        (N178)? mem[5880] : 
                        (N180)? mem[5953] : 
                        (N182)? mem[6026] : 
                        (N184)? mem[6099] : 
                        (N186)? mem[6172] : 
                        (N188)? mem[6245] : 
                        (N190)? mem[6318] : 
                        (N192)? mem[6391] : 
                        (N194)? mem[6464] : 
                        (N196)? mem[6537] : 
                        (N198)? mem[6610] : 
                        (N200)? mem[6683] : 
                        (N202)? mem[6756] : 
                        (N204)? mem[6829] : 
                        (N206)? mem[6902] : 
                        (N208)? mem[6975] : 
                        (N210)? mem[7048] : 
                        (N212)? mem[7121] : 
                        (N214)? mem[7194] : 
                        (N216)? mem[7267] : 
                        (N218)? mem[7340] : 
                        (N220)? mem[7413] : 
                        (N222)? mem[7486] : 
                        (N224)? mem[7559] : 
                        (N226)? mem[7632] : 
                        (N228)? mem[7705] : 
                        (N230)? mem[7778] : 
                        (N232)? mem[7851] : 
                        (N234)? mem[7924] : 
                        (N236)? mem[7997] : 
                        (N238)? mem[8070] : 
                        (N240)? mem[8143] : 
                        (N242)? mem[8216] : 
                        (N244)? mem[8289] : 
                        (N246)? mem[8362] : 
                        (N248)? mem[8435] : 
                        (N250)? mem[8508] : 
                        (N252)? mem[8581] : 
                        (N254)? mem[8654] : 
                        (N256)? mem[8727] : 
                        (N258)? mem[8800] : 
                        (N260)? mem[8873] : 
                        (N262)? mem[8946] : 
                        (N264)? mem[9019] : 
                        (N266)? mem[9092] : 
                        (N268)? mem[9165] : 
                        (N270)? mem[9238] : 
                        (N272)? mem[9311] : 1'b0;
  assign r_data_o[39] = (N145)? mem[39] : 
                        (N147)? mem[112] : 
                        (N149)? mem[185] : 
                        (N151)? mem[258] : 
                        (N153)? mem[331] : 
                        (N155)? mem[404] : 
                        (N157)? mem[477] : 
                        (N159)? mem[550] : 
                        (N161)? mem[623] : 
                        (N163)? mem[696] : 
                        (N165)? mem[769] : 
                        (N167)? mem[842] : 
                        (N169)? mem[915] : 
                        (N171)? mem[988] : 
                        (N173)? mem[1061] : 
                        (N175)? mem[1134] : 
                        (N177)? mem[1207] : 
                        (N179)? mem[1280] : 
                        (N181)? mem[1353] : 
                        (N183)? mem[1426] : 
                        (N185)? mem[1499] : 
                        (N187)? mem[1572] : 
                        (N189)? mem[1645] : 
                        (N191)? mem[1718] : 
                        (N193)? mem[1791] : 
                        (N195)? mem[1864] : 
                        (N197)? mem[1937] : 
                        (N199)? mem[2010] : 
                        (N201)? mem[2083] : 
                        (N203)? mem[2156] : 
                        (N205)? mem[2229] : 
                        (N207)? mem[2302] : 
                        (N209)? mem[2375] : 
                        (N211)? mem[2448] : 
                        (N213)? mem[2521] : 
                        (N215)? mem[2594] : 
                        (N217)? mem[2667] : 
                        (N219)? mem[2740] : 
                        (N221)? mem[2813] : 
                        (N223)? mem[2886] : 
                        (N225)? mem[2959] : 
                        (N227)? mem[3032] : 
                        (N229)? mem[3105] : 
                        (N231)? mem[3178] : 
                        (N233)? mem[3251] : 
                        (N235)? mem[3324] : 
                        (N237)? mem[3397] : 
                        (N239)? mem[3470] : 
                        (N241)? mem[3543] : 
                        (N243)? mem[3616] : 
                        (N245)? mem[3689] : 
                        (N247)? mem[3762] : 
                        (N249)? mem[3835] : 
                        (N251)? mem[3908] : 
                        (N253)? mem[3981] : 
                        (N255)? mem[4054] : 
                        (N257)? mem[4127] : 
                        (N259)? mem[4200] : 
                        (N261)? mem[4273] : 
                        (N263)? mem[4346] : 
                        (N265)? mem[4419] : 
                        (N267)? mem[4492] : 
                        (N269)? mem[4565] : 
                        (N271)? mem[4638] : 
                        (N146)? mem[4711] : 
                        (N148)? mem[4784] : 
                        (N150)? mem[4857] : 
                        (N152)? mem[4930] : 
                        (N154)? mem[5003] : 
                        (N156)? mem[5076] : 
                        (N158)? mem[5149] : 
                        (N160)? mem[5222] : 
                        (N162)? mem[5295] : 
                        (N164)? mem[5368] : 
                        (N166)? mem[5441] : 
                        (N168)? mem[5514] : 
                        (N170)? mem[5587] : 
                        (N172)? mem[5660] : 
                        (N174)? mem[5733] : 
                        (N176)? mem[5806] : 
                        (N178)? mem[5879] : 
                        (N180)? mem[5952] : 
                        (N182)? mem[6025] : 
                        (N184)? mem[6098] : 
                        (N186)? mem[6171] : 
                        (N188)? mem[6244] : 
                        (N190)? mem[6317] : 
                        (N192)? mem[6390] : 
                        (N194)? mem[6463] : 
                        (N196)? mem[6536] : 
                        (N198)? mem[6609] : 
                        (N200)? mem[6682] : 
                        (N202)? mem[6755] : 
                        (N204)? mem[6828] : 
                        (N206)? mem[6901] : 
                        (N208)? mem[6974] : 
                        (N210)? mem[7047] : 
                        (N212)? mem[7120] : 
                        (N214)? mem[7193] : 
                        (N216)? mem[7266] : 
                        (N218)? mem[7339] : 
                        (N220)? mem[7412] : 
                        (N222)? mem[7485] : 
                        (N224)? mem[7558] : 
                        (N226)? mem[7631] : 
                        (N228)? mem[7704] : 
                        (N230)? mem[7777] : 
                        (N232)? mem[7850] : 
                        (N234)? mem[7923] : 
                        (N236)? mem[7996] : 
                        (N238)? mem[8069] : 
                        (N240)? mem[8142] : 
                        (N242)? mem[8215] : 
                        (N244)? mem[8288] : 
                        (N246)? mem[8361] : 
                        (N248)? mem[8434] : 
                        (N250)? mem[8507] : 
                        (N252)? mem[8580] : 
                        (N254)? mem[8653] : 
                        (N256)? mem[8726] : 
                        (N258)? mem[8799] : 
                        (N260)? mem[8872] : 
                        (N262)? mem[8945] : 
                        (N264)? mem[9018] : 
                        (N266)? mem[9091] : 
                        (N268)? mem[9164] : 
                        (N270)? mem[9237] : 
                        (N272)? mem[9310] : 1'b0;
  assign r_data_o[38] = (N145)? mem[38] : 
                        (N147)? mem[111] : 
                        (N149)? mem[184] : 
                        (N151)? mem[257] : 
                        (N153)? mem[330] : 
                        (N155)? mem[403] : 
                        (N157)? mem[476] : 
                        (N159)? mem[549] : 
                        (N161)? mem[622] : 
                        (N163)? mem[695] : 
                        (N165)? mem[768] : 
                        (N167)? mem[841] : 
                        (N169)? mem[914] : 
                        (N171)? mem[987] : 
                        (N173)? mem[1060] : 
                        (N175)? mem[1133] : 
                        (N177)? mem[1206] : 
                        (N179)? mem[1279] : 
                        (N181)? mem[1352] : 
                        (N183)? mem[1425] : 
                        (N185)? mem[1498] : 
                        (N187)? mem[1571] : 
                        (N189)? mem[1644] : 
                        (N191)? mem[1717] : 
                        (N193)? mem[1790] : 
                        (N195)? mem[1863] : 
                        (N197)? mem[1936] : 
                        (N199)? mem[2009] : 
                        (N201)? mem[2082] : 
                        (N203)? mem[2155] : 
                        (N205)? mem[2228] : 
                        (N207)? mem[2301] : 
                        (N209)? mem[2374] : 
                        (N211)? mem[2447] : 
                        (N213)? mem[2520] : 
                        (N215)? mem[2593] : 
                        (N217)? mem[2666] : 
                        (N219)? mem[2739] : 
                        (N221)? mem[2812] : 
                        (N223)? mem[2885] : 
                        (N225)? mem[2958] : 
                        (N227)? mem[3031] : 
                        (N229)? mem[3104] : 
                        (N231)? mem[3177] : 
                        (N233)? mem[3250] : 
                        (N235)? mem[3323] : 
                        (N237)? mem[3396] : 
                        (N239)? mem[3469] : 
                        (N241)? mem[3542] : 
                        (N243)? mem[3615] : 
                        (N245)? mem[3688] : 
                        (N247)? mem[3761] : 
                        (N249)? mem[3834] : 
                        (N251)? mem[3907] : 
                        (N253)? mem[3980] : 
                        (N255)? mem[4053] : 
                        (N257)? mem[4126] : 
                        (N259)? mem[4199] : 
                        (N261)? mem[4272] : 
                        (N263)? mem[4345] : 
                        (N265)? mem[4418] : 
                        (N267)? mem[4491] : 
                        (N269)? mem[4564] : 
                        (N271)? mem[4637] : 
                        (N146)? mem[4710] : 
                        (N148)? mem[4783] : 
                        (N150)? mem[4856] : 
                        (N152)? mem[4929] : 
                        (N154)? mem[5002] : 
                        (N156)? mem[5075] : 
                        (N158)? mem[5148] : 
                        (N160)? mem[5221] : 
                        (N162)? mem[5294] : 
                        (N164)? mem[5367] : 
                        (N166)? mem[5440] : 
                        (N168)? mem[5513] : 
                        (N170)? mem[5586] : 
                        (N172)? mem[5659] : 
                        (N174)? mem[5732] : 
                        (N176)? mem[5805] : 
                        (N178)? mem[5878] : 
                        (N180)? mem[5951] : 
                        (N182)? mem[6024] : 
                        (N184)? mem[6097] : 
                        (N186)? mem[6170] : 
                        (N188)? mem[6243] : 
                        (N190)? mem[6316] : 
                        (N192)? mem[6389] : 
                        (N194)? mem[6462] : 
                        (N196)? mem[6535] : 
                        (N198)? mem[6608] : 
                        (N200)? mem[6681] : 
                        (N202)? mem[6754] : 
                        (N204)? mem[6827] : 
                        (N206)? mem[6900] : 
                        (N208)? mem[6973] : 
                        (N210)? mem[7046] : 
                        (N212)? mem[7119] : 
                        (N214)? mem[7192] : 
                        (N216)? mem[7265] : 
                        (N218)? mem[7338] : 
                        (N220)? mem[7411] : 
                        (N222)? mem[7484] : 
                        (N224)? mem[7557] : 
                        (N226)? mem[7630] : 
                        (N228)? mem[7703] : 
                        (N230)? mem[7776] : 
                        (N232)? mem[7849] : 
                        (N234)? mem[7922] : 
                        (N236)? mem[7995] : 
                        (N238)? mem[8068] : 
                        (N240)? mem[8141] : 
                        (N242)? mem[8214] : 
                        (N244)? mem[8287] : 
                        (N246)? mem[8360] : 
                        (N248)? mem[8433] : 
                        (N250)? mem[8506] : 
                        (N252)? mem[8579] : 
                        (N254)? mem[8652] : 
                        (N256)? mem[8725] : 
                        (N258)? mem[8798] : 
                        (N260)? mem[8871] : 
                        (N262)? mem[8944] : 
                        (N264)? mem[9017] : 
                        (N266)? mem[9090] : 
                        (N268)? mem[9163] : 
                        (N270)? mem[9236] : 
                        (N272)? mem[9309] : 1'b0;
  assign r_data_o[37] = (N145)? mem[37] : 
                        (N147)? mem[110] : 
                        (N149)? mem[183] : 
                        (N151)? mem[256] : 
                        (N153)? mem[329] : 
                        (N155)? mem[402] : 
                        (N157)? mem[475] : 
                        (N159)? mem[548] : 
                        (N161)? mem[621] : 
                        (N163)? mem[694] : 
                        (N165)? mem[767] : 
                        (N167)? mem[840] : 
                        (N169)? mem[913] : 
                        (N171)? mem[986] : 
                        (N173)? mem[1059] : 
                        (N175)? mem[1132] : 
                        (N177)? mem[1205] : 
                        (N179)? mem[1278] : 
                        (N181)? mem[1351] : 
                        (N183)? mem[1424] : 
                        (N185)? mem[1497] : 
                        (N187)? mem[1570] : 
                        (N189)? mem[1643] : 
                        (N191)? mem[1716] : 
                        (N193)? mem[1789] : 
                        (N195)? mem[1862] : 
                        (N197)? mem[1935] : 
                        (N199)? mem[2008] : 
                        (N201)? mem[2081] : 
                        (N203)? mem[2154] : 
                        (N205)? mem[2227] : 
                        (N207)? mem[2300] : 
                        (N209)? mem[2373] : 
                        (N211)? mem[2446] : 
                        (N213)? mem[2519] : 
                        (N215)? mem[2592] : 
                        (N217)? mem[2665] : 
                        (N219)? mem[2738] : 
                        (N221)? mem[2811] : 
                        (N223)? mem[2884] : 
                        (N225)? mem[2957] : 
                        (N227)? mem[3030] : 
                        (N229)? mem[3103] : 
                        (N231)? mem[3176] : 
                        (N233)? mem[3249] : 
                        (N235)? mem[3322] : 
                        (N237)? mem[3395] : 
                        (N239)? mem[3468] : 
                        (N241)? mem[3541] : 
                        (N243)? mem[3614] : 
                        (N245)? mem[3687] : 
                        (N247)? mem[3760] : 
                        (N249)? mem[3833] : 
                        (N251)? mem[3906] : 
                        (N253)? mem[3979] : 
                        (N255)? mem[4052] : 
                        (N257)? mem[4125] : 
                        (N259)? mem[4198] : 
                        (N261)? mem[4271] : 
                        (N263)? mem[4344] : 
                        (N265)? mem[4417] : 
                        (N267)? mem[4490] : 
                        (N269)? mem[4563] : 
                        (N271)? mem[4636] : 
                        (N146)? mem[4709] : 
                        (N148)? mem[4782] : 
                        (N150)? mem[4855] : 
                        (N152)? mem[4928] : 
                        (N154)? mem[5001] : 
                        (N156)? mem[5074] : 
                        (N158)? mem[5147] : 
                        (N160)? mem[5220] : 
                        (N162)? mem[5293] : 
                        (N164)? mem[5366] : 
                        (N166)? mem[5439] : 
                        (N168)? mem[5512] : 
                        (N170)? mem[5585] : 
                        (N172)? mem[5658] : 
                        (N174)? mem[5731] : 
                        (N176)? mem[5804] : 
                        (N178)? mem[5877] : 
                        (N180)? mem[5950] : 
                        (N182)? mem[6023] : 
                        (N184)? mem[6096] : 
                        (N186)? mem[6169] : 
                        (N188)? mem[6242] : 
                        (N190)? mem[6315] : 
                        (N192)? mem[6388] : 
                        (N194)? mem[6461] : 
                        (N196)? mem[6534] : 
                        (N198)? mem[6607] : 
                        (N200)? mem[6680] : 
                        (N202)? mem[6753] : 
                        (N204)? mem[6826] : 
                        (N206)? mem[6899] : 
                        (N208)? mem[6972] : 
                        (N210)? mem[7045] : 
                        (N212)? mem[7118] : 
                        (N214)? mem[7191] : 
                        (N216)? mem[7264] : 
                        (N218)? mem[7337] : 
                        (N220)? mem[7410] : 
                        (N222)? mem[7483] : 
                        (N224)? mem[7556] : 
                        (N226)? mem[7629] : 
                        (N228)? mem[7702] : 
                        (N230)? mem[7775] : 
                        (N232)? mem[7848] : 
                        (N234)? mem[7921] : 
                        (N236)? mem[7994] : 
                        (N238)? mem[8067] : 
                        (N240)? mem[8140] : 
                        (N242)? mem[8213] : 
                        (N244)? mem[8286] : 
                        (N246)? mem[8359] : 
                        (N248)? mem[8432] : 
                        (N250)? mem[8505] : 
                        (N252)? mem[8578] : 
                        (N254)? mem[8651] : 
                        (N256)? mem[8724] : 
                        (N258)? mem[8797] : 
                        (N260)? mem[8870] : 
                        (N262)? mem[8943] : 
                        (N264)? mem[9016] : 
                        (N266)? mem[9089] : 
                        (N268)? mem[9162] : 
                        (N270)? mem[9235] : 
                        (N272)? mem[9308] : 1'b0;
  assign r_data_o[36] = (N145)? mem[36] : 
                        (N147)? mem[109] : 
                        (N149)? mem[182] : 
                        (N151)? mem[255] : 
                        (N153)? mem[328] : 
                        (N155)? mem[401] : 
                        (N157)? mem[474] : 
                        (N159)? mem[547] : 
                        (N161)? mem[620] : 
                        (N163)? mem[693] : 
                        (N165)? mem[766] : 
                        (N167)? mem[839] : 
                        (N169)? mem[912] : 
                        (N171)? mem[985] : 
                        (N173)? mem[1058] : 
                        (N175)? mem[1131] : 
                        (N177)? mem[1204] : 
                        (N179)? mem[1277] : 
                        (N181)? mem[1350] : 
                        (N183)? mem[1423] : 
                        (N185)? mem[1496] : 
                        (N187)? mem[1569] : 
                        (N189)? mem[1642] : 
                        (N191)? mem[1715] : 
                        (N193)? mem[1788] : 
                        (N195)? mem[1861] : 
                        (N197)? mem[1934] : 
                        (N199)? mem[2007] : 
                        (N201)? mem[2080] : 
                        (N203)? mem[2153] : 
                        (N205)? mem[2226] : 
                        (N207)? mem[2299] : 
                        (N209)? mem[2372] : 
                        (N211)? mem[2445] : 
                        (N213)? mem[2518] : 
                        (N215)? mem[2591] : 
                        (N217)? mem[2664] : 
                        (N219)? mem[2737] : 
                        (N221)? mem[2810] : 
                        (N223)? mem[2883] : 
                        (N225)? mem[2956] : 
                        (N227)? mem[3029] : 
                        (N229)? mem[3102] : 
                        (N231)? mem[3175] : 
                        (N233)? mem[3248] : 
                        (N235)? mem[3321] : 
                        (N237)? mem[3394] : 
                        (N239)? mem[3467] : 
                        (N241)? mem[3540] : 
                        (N243)? mem[3613] : 
                        (N245)? mem[3686] : 
                        (N247)? mem[3759] : 
                        (N249)? mem[3832] : 
                        (N251)? mem[3905] : 
                        (N253)? mem[3978] : 
                        (N255)? mem[4051] : 
                        (N257)? mem[4124] : 
                        (N259)? mem[4197] : 
                        (N261)? mem[4270] : 
                        (N263)? mem[4343] : 
                        (N265)? mem[4416] : 
                        (N267)? mem[4489] : 
                        (N269)? mem[4562] : 
                        (N271)? mem[4635] : 
                        (N146)? mem[4708] : 
                        (N148)? mem[4781] : 
                        (N150)? mem[4854] : 
                        (N152)? mem[4927] : 
                        (N154)? mem[5000] : 
                        (N156)? mem[5073] : 
                        (N158)? mem[5146] : 
                        (N160)? mem[5219] : 
                        (N162)? mem[5292] : 
                        (N164)? mem[5365] : 
                        (N166)? mem[5438] : 
                        (N168)? mem[5511] : 
                        (N170)? mem[5584] : 
                        (N172)? mem[5657] : 
                        (N174)? mem[5730] : 
                        (N176)? mem[5803] : 
                        (N178)? mem[5876] : 
                        (N180)? mem[5949] : 
                        (N182)? mem[6022] : 
                        (N184)? mem[6095] : 
                        (N186)? mem[6168] : 
                        (N188)? mem[6241] : 
                        (N190)? mem[6314] : 
                        (N192)? mem[6387] : 
                        (N194)? mem[6460] : 
                        (N196)? mem[6533] : 
                        (N198)? mem[6606] : 
                        (N200)? mem[6679] : 
                        (N202)? mem[6752] : 
                        (N204)? mem[6825] : 
                        (N206)? mem[6898] : 
                        (N208)? mem[6971] : 
                        (N210)? mem[7044] : 
                        (N212)? mem[7117] : 
                        (N214)? mem[7190] : 
                        (N216)? mem[7263] : 
                        (N218)? mem[7336] : 
                        (N220)? mem[7409] : 
                        (N222)? mem[7482] : 
                        (N224)? mem[7555] : 
                        (N226)? mem[7628] : 
                        (N228)? mem[7701] : 
                        (N230)? mem[7774] : 
                        (N232)? mem[7847] : 
                        (N234)? mem[7920] : 
                        (N236)? mem[7993] : 
                        (N238)? mem[8066] : 
                        (N240)? mem[8139] : 
                        (N242)? mem[8212] : 
                        (N244)? mem[8285] : 
                        (N246)? mem[8358] : 
                        (N248)? mem[8431] : 
                        (N250)? mem[8504] : 
                        (N252)? mem[8577] : 
                        (N254)? mem[8650] : 
                        (N256)? mem[8723] : 
                        (N258)? mem[8796] : 
                        (N260)? mem[8869] : 
                        (N262)? mem[8942] : 
                        (N264)? mem[9015] : 
                        (N266)? mem[9088] : 
                        (N268)? mem[9161] : 
                        (N270)? mem[9234] : 
                        (N272)? mem[9307] : 1'b0;
  assign r_data_o[35] = (N145)? mem[35] : 
                        (N147)? mem[108] : 
                        (N149)? mem[181] : 
                        (N151)? mem[254] : 
                        (N153)? mem[327] : 
                        (N155)? mem[400] : 
                        (N157)? mem[473] : 
                        (N159)? mem[546] : 
                        (N161)? mem[619] : 
                        (N163)? mem[692] : 
                        (N165)? mem[765] : 
                        (N167)? mem[838] : 
                        (N169)? mem[911] : 
                        (N171)? mem[984] : 
                        (N173)? mem[1057] : 
                        (N175)? mem[1130] : 
                        (N177)? mem[1203] : 
                        (N179)? mem[1276] : 
                        (N181)? mem[1349] : 
                        (N183)? mem[1422] : 
                        (N185)? mem[1495] : 
                        (N187)? mem[1568] : 
                        (N189)? mem[1641] : 
                        (N191)? mem[1714] : 
                        (N193)? mem[1787] : 
                        (N195)? mem[1860] : 
                        (N197)? mem[1933] : 
                        (N199)? mem[2006] : 
                        (N201)? mem[2079] : 
                        (N203)? mem[2152] : 
                        (N205)? mem[2225] : 
                        (N207)? mem[2298] : 
                        (N209)? mem[2371] : 
                        (N211)? mem[2444] : 
                        (N213)? mem[2517] : 
                        (N215)? mem[2590] : 
                        (N217)? mem[2663] : 
                        (N219)? mem[2736] : 
                        (N221)? mem[2809] : 
                        (N223)? mem[2882] : 
                        (N225)? mem[2955] : 
                        (N227)? mem[3028] : 
                        (N229)? mem[3101] : 
                        (N231)? mem[3174] : 
                        (N233)? mem[3247] : 
                        (N235)? mem[3320] : 
                        (N237)? mem[3393] : 
                        (N239)? mem[3466] : 
                        (N241)? mem[3539] : 
                        (N243)? mem[3612] : 
                        (N245)? mem[3685] : 
                        (N247)? mem[3758] : 
                        (N249)? mem[3831] : 
                        (N251)? mem[3904] : 
                        (N253)? mem[3977] : 
                        (N255)? mem[4050] : 
                        (N257)? mem[4123] : 
                        (N259)? mem[4196] : 
                        (N261)? mem[4269] : 
                        (N263)? mem[4342] : 
                        (N265)? mem[4415] : 
                        (N267)? mem[4488] : 
                        (N269)? mem[4561] : 
                        (N271)? mem[4634] : 
                        (N146)? mem[4707] : 
                        (N148)? mem[4780] : 
                        (N150)? mem[4853] : 
                        (N152)? mem[4926] : 
                        (N154)? mem[4999] : 
                        (N156)? mem[5072] : 
                        (N158)? mem[5145] : 
                        (N160)? mem[5218] : 
                        (N162)? mem[5291] : 
                        (N164)? mem[5364] : 
                        (N166)? mem[5437] : 
                        (N168)? mem[5510] : 
                        (N170)? mem[5583] : 
                        (N172)? mem[5656] : 
                        (N174)? mem[5729] : 
                        (N176)? mem[5802] : 
                        (N178)? mem[5875] : 
                        (N180)? mem[5948] : 
                        (N182)? mem[6021] : 
                        (N184)? mem[6094] : 
                        (N186)? mem[6167] : 
                        (N188)? mem[6240] : 
                        (N190)? mem[6313] : 
                        (N192)? mem[6386] : 
                        (N194)? mem[6459] : 
                        (N196)? mem[6532] : 
                        (N198)? mem[6605] : 
                        (N200)? mem[6678] : 
                        (N202)? mem[6751] : 
                        (N204)? mem[6824] : 
                        (N206)? mem[6897] : 
                        (N208)? mem[6970] : 
                        (N210)? mem[7043] : 
                        (N212)? mem[7116] : 
                        (N214)? mem[7189] : 
                        (N216)? mem[7262] : 
                        (N218)? mem[7335] : 
                        (N220)? mem[7408] : 
                        (N222)? mem[7481] : 
                        (N224)? mem[7554] : 
                        (N226)? mem[7627] : 
                        (N228)? mem[7700] : 
                        (N230)? mem[7773] : 
                        (N232)? mem[7846] : 
                        (N234)? mem[7919] : 
                        (N236)? mem[7992] : 
                        (N238)? mem[8065] : 
                        (N240)? mem[8138] : 
                        (N242)? mem[8211] : 
                        (N244)? mem[8284] : 
                        (N246)? mem[8357] : 
                        (N248)? mem[8430] : 
                        (N250)? mem[8503] : 
                        (N252)? mem[8576] : 
                        (N254)? mem[8649] : 
                        (N256)? mem[8722] : 
                        (N258)? mem[8795] : 
                        (N260)? mem[8868] : 
                        (N262)? mem[8941] : 
                        (N264)? mem[9014] : 
                        (N266)? mem[9087] : 
                        (N268)? mem[9160] : 
                        (N270)? mem[9233] : 
                        (N272)? mem[9306] : 1'b0;
  assign r_data_o[34] = (N145)? mem[34] : 
                        (N147)? mem[107] : 
                        (N149)? mem[180] : 
                        (N151)? mem[253] : 
                        (N153)? mem[326] : 
                        (N155)? mem[399] : 
                        (N157)? mem[472] : 
                        (N159)? mem[545] : 
                        (N161)? mem[618] : 
                        (N163)? mem[691] : 
                        (N165)? mem[764] : 
                        (N167)? mem[837] : 
                        (N169)? mem[910] : 
                        (N171)? mem[983] : 
                        (N173)? mem[1056] : 
                        (N175)? mem[1129] : 
                        (N177)? mem[1202] : 
                        (N179)? mem[1275] : 
                        (N181)? mem[1348] : 
                        (N183)? mem[1421] : 
                        (N185)? mem[1494] : 
                        (N187)? mem[1567] : 
                        (N189)? mem[1640] : 
                        (N191)? mem[1713] : 
                        (N193)? mem[1786] : 
                        (N195)? mem[1859] : 
                        (N197)? mem[1932] : 
                        (N199)? mem[2005] : 
                        (N201)? mem[2078] : 
                        (N203)? mem[2151] : 
                        (N205)? mem[2224] : 
                        (N207)? mem[2297] : 
                        (N209)? mem[2370] : 
                        (N211)? mem[2443] : 
                        (N213)? mem[2516] : 
                        (N215)? mem[2589] : 
                        (N217)? mem[2662] : 
                        (N219)? mem[2735] : 
                        (N221)? mem[2808] : 
                        (N223)? mem[2881] : 
                        (N225)? mem[2954] : 
                        (N227)? mem[3027] : 
                        (N229)? mem[3100] : 
                        (N231)? mem[3173] : 
                        (N233)? mem[3246] : 
                        (N235)? mem[3319] : 
                        (N237)? mem[3392] : 
                        (N239)? mem[3465] : 
                        (N241)? mem[3538] : 
                        (N243)? mem[3611] : 
                        (N245)? mem[3684] : 
                        (N247)? mem[3757] : 
                        (N249)? mem[3830] : 
                        (N251)? mem[3903] : 
                        (N253)? mem[3976] : 
                        (N255)? mem[4049] : 
                        (N257)? mem[4122] : 
                        (N259)? mem[4195] : 
                        (N261)? mem[4268] : 
                        (N263)? mem[4341] : 
                        (N265)? mem[4414] : 
                        (N267)? mem[4487] : 
                        (N269)? mem[4560] : 
                        (N271)? mem[4633] : 
                        (N146)? mem[4706] : 
                        (N148)? mem[4779] : 
                        (N150)? mem[4852] : 
                        (N152)? mem[4925] : 
                        (N154)? mem[4998] : 
                        (N156)? mem[5071] : 
                        (N158)? mem[5144] : 
                        (N160)? mem[5217] : 
                        (N162)? mem[5290] : 
                        (N164)? mem[5363] : 
                        (N166)? mem[5436] : 
                        (N168)? mem[5509] : 
                        (N170)? mem[5582] : 
                        (N172)? mem[5655] : 
                        (N174)? mem[5728] : 
                        (N176)? mem[5801] : 
                        (N178)? mem[5874] : 
                        (N180)? mem[5947] : 
                        (N182)? mem[6020] : 
                        (N184)? mem[6093] : 
                        (N186)? mem[6166] : 
                        (N188)? mem[6239] : 
                        (N190)? mem[6312] : 
                        (N192)? mem[6385] : 
                        (N194)? mem[6458] : 
                        (N196)? mem[6531] : 
                        (N198)? mem[6604] : 
                        (N200)? mem[6677] : 
                        (N202)? mem[6750] : 
                        (N204)? mem[6823] : 
                        (N206)? mem[6896] : 
                        (N208)? mem[6969] : 
                        (N210)? mem[7042] : 
                        (N212)? mem[7115] : 
                        (N214)? mem[7188] : 
                        (N216)? mem[7261] : 
                        (N218)? mem[7334] : 
                        (N220)? mem[7407] : 
                        (N222)? mem[7480] : 
                        (N224)? mem[7553] : 
                        (N226)? mem[7626] : 
                        (N228)? mem[7699] : 
                        (N230)? mem[7772] : 
                        (N232)? mem[7845] : 
                        (N234)? mem[7918] : 
                        (N236)? mem[7991] : 
                        (N238)? mem[8064] : 
                        (N240)? mem[8137] : 
                        (N242)? mem[8210] : 
                        (N244)? mem[8283] : 
                        (N246)? mem[8356] : 
                        (N248)? mem[8429] : 
                        (N250)? mem[8502] : 
                        (N252)? mem[8575] : 
                        (N254)? mem[8648] : 
                        (N256)? mem[8721] : 
                        (N258)? mem[8794] : 
                        (N260)? mem[8867] : 
                        (N262)? mem[8940] : 
                        (N264)? mem[9013] : 
                        (N266)? mem[9086] : 
                        (N268)? mem[9159] : 
                        (N270)? mem[9232] : 
                        (N272)? mem[9305] : 1'b0;
  assign r_data_o[33] = (N145)? mem[33] : 
                        (N147)? mem[106] : 
                        (N149)? mem[179] : 
                        (N151)? mem[252] : 
                        (N153)? mem[325] : 
                        (N155)? mem[398] : 
                        (N157)? mem[471] : 
                        (N159)? mem[544] : 
                        (N161)? mem[617] : 
                        (N163)? mem[690] : 
                        (N165)? mem[763] : 
                        (N167)? mem[836] : 
                        (N169)? mem[909] : 
                        (N171)? mem[982] : 
                        (N173)? mem[1055] : 
                        (N175)? mem[1128] : 
                        (N177)? mem[1201] : 
                        (N179)? mem[1274] : 
                        (N181)? mem[1347] : 
                        (N183)? mem[1420] : 
                        (N185)? mem[1493] : 
                        (N187)? mem[1566] : 
                        (N189)? mem[1639] : 
                        (N191)? mem[1712] : 
                        (N193)? mem[1785] : 
                        (N195)? mem[1858] : 
                        (N197)? mem[1931] : 
                        (N199)? mem[2004] : 
                        (N201)? mem[2077] : 
                        (N203)? mem[2150] : 
                        (N205)? mem[2223] : 
                        (N207)? mem[2296] : 
                        (N209)? mem[2369] : 
                        (N211)? mem[2442] : 
                        (N213)? mem[2515] : 
                        (N215)? mem[2588] : 
                        (N217)? mem[2661] : 
                        (N219)? mem[2734] : 
                        (N221)? mem[2807] : 
                        (N223)? mem[2880] : 
                        (N225)? mem[2953] : 
                        (N227)? mem[3026] : 
                        (N229)? mem[3099] : 
                        (N231)? mem[3172] : 
                        (N233)? mem[3245] : 
                        (N235)? mem[3318] : 
                        (N237)? mem[3391] : 
                        (N239)? mem[3464] : 
                        (N241)? mem[3537] : 
                        (N243)? mem[3610] : 
                        (N245)? mem[3683] : 
                        (N247)? mem[3756] : 
                        (N249)? mem[3829] : 
                        (N251)? mem[3902] : 
                        (N253)? mem[3975] : 
                        (N255)? mem[4048] : 
                        (N257)? mem[4121] : 
                        (N259)? mem[4194] : 
                        (N261)? mem[4267] : 
                        (N263)? mem[4340] : 
                        (N265)? mem[4413] : 
                        (N267)? mem[4486] : 
                        (N269)? mem[4559] : 
                        (N271)? mem[4632] : 
                        (N146)? mem[4705] : 
                        (N148)? mem[4778] : 
                        (N150)? mem[4851] : 
                        (N152)? mem[4924] : 
                        (N154)? mem[4997] : 
                        (N156)? mem[5070] : 
                        (N158)? mem[5143] : 
                        (N160)? mem[5216] : 
                        (N162)? mem[5289] : 
                        (N164)? mem[5362] : 
                        (N166)? mem[5435] : 
                        (N168)? mem[5508] : 
                        (N170)? mem[5581] : 
                        (N172)? mem[5654] : 
                        (N174)? mem[5727] : 
                        (N176)? mem[5800] : 
                        (N178)? mem[5873] : 
                        (N180)? mem[5946] : 
                        (N182)? mem[6019] : 
                        (N184)? mem[6092] : 
                        (N186)? mem[6165] : 
                        (N188)? mem[6238] : 
                        (N190)? mem[6311] : 
                        (N192)? mem[6384] : 
                        (N194)? mem[6457] : 
                        (N196)? mem[6530] : 
                        (N198)? mem[6603] : 
                        (N200)? mem[6676] : 
                        (N202)? mem[6749] : 
                        (N204)? mem[6822] : 
                        (N206)? mem[6895] : 
                        (N208)? mem[6968] : 
                        (N210)? mem[7041] : 
                        (N212)? mem[7114] : 
                        (N214)? mem[7187] : 
                        (N216)? mem[7260] : 
                        (N218)? mem[7333] : 
                        (N220)? mem[7406] : 
                        (N222)? mem[7479] : 
                        (N224)? mem[7552] : 
                        (N226)? mem[7625] : 
                        (N228)? mem[7698] : 
                        (N230)? mem[7771] : 
                        (N232)? mem[7844] : 
                        (N234)? mem[7917] : 
                        (N236)? mem[7990] : 
                        (N238)? mem[8063] : 
                        (N240)? mem[8136] : 
                        (N242)? mem[8209] : 
                        (N244)? mem[8282] : 
                        (N246)? mem[8355] : 
                        (N248)? mem[8428] : 
                        (N250)? mem[8501] : 
                        (N252)? mem[8574] : 
                        (N254)? mem[8647] : 
                        (N256)? mem[8720] : 
                        (N258)? mem[8793] : 
                        (N260)? mem[8866] : 
                        (N262)? mem[8939] : 
                        (N264)? mem[9012] : 
                        (N266)? mem[9085] : 
                        (N268)? mem[9158] : 
                        (N270)? mem[9231] : 
                        (N272)? mem[9304] : 1'b0;
  assign r_data_o[32] = (N145)? mem[32] : 
                        (N147)? mem[105] : 
                        (N149)? mem[178] : 
                        (N151)? mem[251] : 
                        (N153)? mem[324] : 
                        (N155)? mem[397] : 
                        (N157)? mem[470] : 
                        (N159)? mem[543] : 
                        (N161)? mem[616] : 
                        (N163)? mem[689] : 
                        (N165)? mem[762] : 
                        (N167)? mem[835] : 
                        (N169)? mem[908] : 
                        (N171)? mem[981] : 
                        (N173)? mem[1054] : 
                        (N175)? mem[1127] : 
                        (N177)? mem[1200] : 
                        (N179)? mem[1273] : 
                        (N181)? mem[1346] : 
                        (N183)? mem[1419] : 
                        (N185)? mem[1492] : 
                        (N187)? mem[1565] : 
                        (N189)? mem[1638] : 
                        (N191)? mem[1711] : 
                        (N193)? mem[1784] : 
                        (N195)? mem[1857] : 
                        (N197)? mem[1930] : 
                        (N199)? mem[2003] : 
                        (N201)? mem[2076] : 
                        (N203)? mem[2149] : 
                        (N205)? mem[2222] : 
                        (N207)? mem[2295] : 
                        (N209)? mem[2368] : 
                        (N211)? mem[2441] : 
                        (N213)? mem[2514] : 
                        (N215)? mem[2587] : 
                        (N217)? mem[2660] : 
                        (N219)? mem[2733] : 
                        (N221)? mem[2806] : 
                        (N223)? mem[2879] : 
                        (N225)? mem[2952] : 
                        (N227)? mem[3025] : 
                        (N229)? mem[3098] : 
                        (N231)? mem[3171] : 
                        (N233)? mem[3244] : 
                        (N235)? mem[3317] : 
                        (N237)? mem[3390] : 
                        (N239)? mem[3463] : 
                        (N241)? mem[3536] : 
                        (N243)? mem[3609] : 
                        (N245)? mem[3682] : 
                        (N247)? mem[3755] : 
                        (N249)? mem[3828] : 
                        (N251)? mem[3901] : 
                        (N253)? mem[3974] : 
                        (N255)? mem[4047] : 
                        (N257)? mem[4120] : 
                        (N259)? mem[4193] : 
                        (N261)? mem[4266] : 
                        (N263)? mem[4339] : 
                        (N265)? mem[4412] : 
                        (N267)? mem[4485] : 
                        (N269)? mem[4558] : 
                        (N271)? mem[4631] : 
                        (N146)? mem[4704] : 
                        (N148)? mem[4777] : 
                        (N150)? mem[4850] : 
                        (N152)? mem[4923] : 
                        (N154)? mem[4996] : 
                        (N156)? mem[5069] : 
                        (N158)? mem[5142] : 
                        (N160)? mem[5215] : 
                        (N162)? mem[5288] : 
                        (N164)? mem[5361] : 
                        (N166)? mem[5434] : 
                        (N168)? mem[5507] : 
                        (N170)? mem[5580] : 
                        (N172)? mem[5653] : 
                        (N174)? mem[5726] : 
                        (N176)? mem[5799] : 
                        (N178)? mem[5872] : 
                        (N180)? mem[5945] : 
                        (N182)? mem[6018] : 
                        (N184)? mem[6091] : 
                        (N186)? mem[6164] : 
                        (N188)? mem[6237] : 
                        (N190)? mem[6310] : 
                        (N192)? mem[6383] : 
                        (N194)? mem[6456] : 
                        (N196)? mem[6529] : 
                        (N198)? mem[6602] : 
                        (N200)? mem[6675] : 
                        (N202)? mem[6748] : 
                        (N204)? mem[6821] : 
                        (N206)? mem[6894] : 
                        (N208)? mem[6967] : 
                        (N210)? mem[7040] : 
                        (N212)? mem[7113] : 
                        (N214)? mem[7186] : 
                        (N216)? mem[7259] : 
                        (N218)? mem[7332] : 
                        (N220)? mem[7405] : 
                        (N222)? mem[7478] : 
                        (N224)? mem[7551] : 
                        (N226)? mem[7624] : 
                        (N228)? mem[7697] : 
                        (N230)? mem[7770] : 
                        (N232)? mem[7843] : 
                        (N234)? mem[7916] : 
                        (N236)? mem[7989] : 
                        (N238)? mem[8062] : 
                        (N240)? mem[8135] : 
                        (N242)? mem[8208] : 
                        (N244)? mem[8281] : 
                        (N246)? mem[8354] : 
                        (N248)? mem[8427] : 
                        (N250)? mem[8500] : 
                        (N252)? mem[8573] : 
                        (N254)? mem[8646] : 
                        (N256)? mem[8719] : 
                        (N258)? mem[8792] : 
                        (N260)? mem[8865] : 
                        (N262)? mem[8938] : 
                        (N264)? mem[9011] : 
                        (N266)? mem[9084] : 
                        (N268)? mem[9157] : 
                        (N270)? mem[9230] : 
                        (N272)? mem[9303] : 1'b0;
  assign r_data_o[31] = (N145)? mem[31] : 
                        (N147)? mem[104] : 
                        (N149)? mem[177] : 
                        (N151)? mem[250] : 
                        (N153)? mem[323] : 
                        (N155)? mem[396] : 
                        (N157)? mem[469] : 
                        (N159)? mem[542] : 
                        (N161)? mem[615] : 
                        (N163)? mem[688] : 
                        (N165)? mem[761] : 
                        (N167)? mem[834] : 
                        (N169)? mem[907] : 
                        (N171)? mem[980] : 
                        (N173)? mem[1053] : 
                        (N175)? mem[1126] : 
                        (N177)? mem[1199] : 
                        (N179)? mem[1272] : 
                        (N181)? mem[1345] : 
                        (N183)? mem[1418] : 
                        (N185)? mem[1491] : 
                        (N187)? mem[1564] : 
                        (N189)? mem[1637] : 
                        (N191)? mem[1710] : 
                        (N193)? mem[1783] : 
                        (N195)? mem[1856] : 
                        (N197)? mem[1929] : 
                        (N199)? mem[2002] : 
                        (N201)? mem[2075] : 
                        (N203)? mem[2148] : 
                        (N205)? mem[2221] : 
                        (N207)? mem[2294] : 
                        (N209)? mem[2367] : 
                        (N211)? mem[2440] : 
                        (N213)? mem[2513] : 
                        (N215)? mem[2586] : 
                        (N217)? mem[2659] : 
                        (N219)? mem[2732] : 
                        (N221)? mem[2805] : 
                        (N223)? mem[2878] : 
                        (N225)? mem[2951] : 
                        (N227)? mem[3024] : 
                        (N229)? mem[3097] : 
                        (N231)? mem[3170] : 
                        (N233)? mem[3243] : 
                        (N235)? mem[3316] : 
                        (N237)? mem[3389] : 
                        (N239)? mem[3462] : 
                        (N241)? mem[3535] : 
                        (N243)? mem[3608] : 
                        (N245)? mem[3681] : 
                        (N247)? mem[3754] : 
                        (N249)? mem[3827] : 
                        (N251)? mem[3900] : 
                        (N253)? mem[3973] : 
                        (N255)? mem[4046] : 
                        (N257)? mem[4119] : 
                        (N259)? mem[4192] : 
                        (N261)? mem[4265] : 
                        (N263)? mem[4338] : 
                        (N265)? mem[4411] : 
                        (N267)? mem[4484] : 
                        (N269)? mem[4557] : 
                        (N271)? mem[4630] : 
                        (N146)? mem[4703] : 
                        (N148)? mem[4776] : 
                        (N150)? mem[4849] : 
                        (N152)? mem[4922] : 
                        (N154)? mem[4995] : 
                        (N156)? mem[5068] : 
                        (N158)? mem[5141] : 
                        (N160)? mem[5214] : 
                        (N162)? mem[5287] : 
                        (N164)? mem[5360] : 
                        (N166)? mem[5433] : 
                        (N168)? mem[5506] : 
                        (N170)? mem[5579] : 
                        (N172)? mem[5652] : 
                        (N174)? mem[5725] : 
                        (N176)? mem[5798] : 
                        (N178)? mem[5871] : 
                        (N180)? mem[5944] : 
                        (N182)? mem[6017] : 
                        (N184)? mem[6090] : 
                        (N186)? mem[6163] : 
                        (N188)? mem[6236] : 
                        (N190)? mem[6309] : 
                        (N192)? mem[6382] : 
                        (N194)? mem[6455] : 
                        (N196)? mem[6528] : 
                        (N198)? mem[6601] : 
                        (N200)? mem[6674] : 
                        (N202)? mem[6747] : 
                        (N204)? mem[6820] : 
                        (N206)? mem[6893] : 
                        (N208)? mem[6966] : 
                        (N210)? mem[7039] : 
                        (N212)? mem[7112] : 
                        (N214)? mem[7185] : 
                        (N216)? mem[7258] : 
                        (N218)? mem[7331] : 
                        (N220)? mem[7404] : 
                        (N222)? mem[7477] : 
                        (N224)? mem[7550] : 
                        (N226)? mem[7623] : 
                        (N228)? mem[7696] : 
                        (N230)? mem[7769] : 
                        (N232)? mem[7842] : 
                        (N234)? mem[7915] : 
                        (N236)? mem[7988] : 
                        (N238)? mem[8061] : 
                        (N240)? mem[8134] : 
                        (N242)? mem[8207] : 
                        (N244)? mem[8280] : 
                        (N246)? mem[8353] : 
                        (N248)? mem[8426] : 
                        (N250)? mem[8499] : 
                        (N252)? mem[8572] : 
                        (N254)? mem[8645] : 
                        (N256)? mem[8718] : 
                        (N258)? mem[8791] : 
                        (N260)? mem[8864] : 
                        (N262)? mem[8937] : 
                        (N264)? mem[9010] : 
                        (N266)? mem[9083] : 
                        (N268)? mem[9156] : 
                        (N270)? mem[9229] : 
                        (N272)? mem[9302] : 1'b0;
  assign r_data_o[30] = (N145)? mem[30] : 
                        (N147)? mem[103] : 
                        (N149)? mem[176] : 
                        (N151)? mem[249] : 
                        (N153)? mem[322] : 
                        (N155)? mem[395] : 
                        (N157)? mem[468] : 
                        (N159)? mem[541] : 
                        (N161)? mem[614] : 
                        (N163)? mem[687] : 
                        (N165)? mem[760] : 
                        (N167)? mem[833] : 
                        (N169)? mem[906] : 
                        (N171)? mem[979] : 
                        (N173)? mem[1052] : 
                        (N175)? mem[1125] : 
                        (N177)? mem[1198] : 
                        (N179)? mem[1271] : 
                        (N181)? mem[1344] : 
                        (N183)? mem[1417] : 
                        (N185)? mem[1490] : 
                        (N187)? mem[1563] : 
                        (N189)? mem[1636] : 
                        (N191)? mem[1709] : 
                        (N193)? mem[1782] : 
                        (N195)? mem[1855] : 
                        (N197)? mem[1928] : 
                        (N199)? mem[2001] : 
                        (N201)? mem[2074] : 
                        (N203)? mem[2147] : 
                        (N205)? mem[2220] : 
                        (N207)? mem[2293] : 
                        (N209)? mem[2366] : 
                        (N211)? mem[2439] : 
                        (N213)? mem[2512] : 
                        (N215)? mem[2585] : 
                        (N217)? mem[2658] : 
                        (N219)? mem[2731] : 
                        (N221)? mem[2804] : 
                        (N223)? mem[2877] : 
                        (N225)? mem[2950] : 
                        (N227)? mem[3023] : 
                        (N229)? mem[3096] : 
                        (N231)? mem[3169] : 
                        (N233)? mem[3242] : 
                        (N235)? mem[3315] : 
                        (N237)? mem[3388] : 
                        (N239)? mem[3461] : 
                        (N241)? mem[3534] : 
                        (N243)? mem[3607] : 
                        (N245)? mem[3680] : 
                        (N247)? mem[3753] : 
                        (N249)? mem[3826] : 
                        (N251)? mem[3899] : 
                        (N253)? mem[3972] : 
                        (N255)? mem[4045] : 
                        (N257)? mem[4118] : 
                        (N259)? mem[4191] : 
                        (N261)? mem[4264] : 
                        (N263)? mem[4337] : 
                        (N265)? mem[4410] : 
                        (N267)? mem[4483] : 
                        (N269)? mem[4556] : 
                        (N271)? mem[4629] : 
                        (N146)? mem[4702] : 
                        (N148)? mem[4775] : 
                        (N150)? mem[4848] : 
                        (N152)? mem[4921] : 
                        (N154)? mem[4994] : 
                        (N156)? mem[5067] : 
                        (N158)? mem[5140] : 
                        (N160)? mem[5213] : 
                        (N162)? mem[5286] : 
                        (N164)? mem[5359] : 
                        (N166)? mem[5432] : 
                        (N168)? mem[5505] : 
                        (N170)? mem[5578] : 
                        (N172)? mem[5651] : 
                        (N174)? mem[5724] : 
                        (N176)? mem[5797] : 
                        (N178)? mem[5870] : 
                        (N180)? mem[5943] : 
                        (N182)? mem[6016] : 
                        (N184)? mem[6089] : 
                        (N186)? mem[6162] : 
                        (N188)? mem[6235] : 
                        (N190)? mem[6308] : 
                        (N192)? mem[6381] : 
                        (N194)? mem[6454] : 
                        (N196)? mem[6527] : 
                        (N198)? mem[6600] : 
                        (N200)? mem[6673] : 
                        (N202)? mem[6746] : 
                        (N204)? mem[6819] : 
                        (N206)? mem[6892] : 
                        (N208)? mem[6965] : 
                        (N210)? mem[7038] : 
                        (N212)? mem[7111] : 
                        (N214)? mem[7184] : 
                        (N216)? mem[7257] : 
                        (N218)? mem[7330] : 
                        (N220)? mem[7403] : 
                        (N222)? mem[7476] : 
                        (N224)? mem[7549] : 
                        (N226)? mem[7622] : 
                        (N228)? mem[7695] : 
                        (N230)? mem[7768] : 
                        (N232)? mem[7841] : 
                        (N234)? mem[7914] : 
                        (N236)? mem[7987] : 
                        (N238)? mem[8060] : 
                        (N240)? mem[8133] : 
                        (N242)? mem[8206] : 
                        (N244)? mem[8279] : 
                        (N246)? mem[8352] : 
                        (N248)? mem[8425] : 
                        (N250)? mem[8498] : 
                        (N252)? mem[8571] : 
                        (N254)? mem[8644] : 
                        (N256)? mem[8717] : 
                        (N258)? mem[8790] : 
                        (N260)? mem[8863] : 
                        (N262)? mem[8936] : 
                        (N264)? mem[9009] : 
                        (N266)? mem[9082] : 
                        (N268)? mem[9155] : 
                        (N270)? mem[9228] : 
                        (N272)? mem[9301] : 1'b0;
  assign r_data_o[29] = (N145)? mem[29] : 
                        (N147)? mem[102] : 
                        (N149)? mem[175] : 
                        (N151)? mem[248] : 
                        (N153)? mem[321] : 
                        (N155)? mem[394] : 
                        (N157)? mem[467] : 
                        (N159)? mem[540] : 
                        (N161)? mem[613] : 
                        (N163)? mem[686] : 
                        (N165)? mem[759] : 
                        (N167)? mem[832] : 
                        (N169)? mem[905] : 
                        (N171)? mem[978] : 
                        (N173)? mem[1051] : 
                        (N175)? mem[1124] : 
                        (N177)? mem[1197] : 
                        (N179)? mem[1270] : 
                        (N181)? mem[1343] : 
                        (N183)? mem[1416] : 
                        (N185)? mem[1489] : 
                        (N187)? mem[1562] : 
                        (N189)? mem[1635] : 
                        (N191)? mem[1708] : 
                        (N193)? mem[1781] : 
                        (N195)? mem[1854] : 
                        (N197)? mem[1927] : 
                        (N199)? mem[2000] : 
                        (N201)? mem[2073] : 
                        (N203)? mem[2146] : 
                        (N205)? mem[2219] : 
                        (N207)? mem[2292] : 
                        (N209)? mem[2365] : 
                        (N211)? mem[2438] : 
                        (N213)? mem[2511] : 
                        (N215)? mem[2584] : 
                        (N217)? mem[2657] : 
                        (N219)? mem[2730] : 
                        (N221)? mem[2803] : 
                        (N223)? mem[2876] : 
                        (N225)? mem[2949] : 
                        (N227)? mem[3022] : 
                        (N229)? mem[3095] : 
                        (N231)? mem[3168] : 
                        (N233)? mem[3241] : 
                        (N235)? mem[3314] : 
                        (N237)? mem[3387] : 
                        (N239)? mem[3460] : 
                        (N241)? mem[3533] : 
                        (N243)? mem[3606] : 
                        (N245)? mem[3679] : 
                        (N247)? mem[3752] : 
                        (N249)? mem[3825] : 
                        (N251)? mem[3898] : 
                        (N253)? mem[3971] : 
                        (N255)? mem[4044] : 
                        (N257)? mem[4117] : 
                        (N259)? mem[4190] : 
                        (N261)? mem[4263] : 
                        (N263)? mem[4336] : 
                        (N265)? mem[4409] : 
                        (N267)? mem[4482] : 
                        (N269)? mem[4555] : 
                        (N271)? mem[4628] : 
                        (N146)? mem[4701] : 
                        (N148)? mem[4774] : 
                        (N150)? mem[4847] : 
                        (N152)? mem[4920] : 
                        (N154)? mem[4993] : 
                        (N156)? mem[5066] : 
                        (N158)? mem[5139] : 
                        (N160)? mem[5212] : 
                        (N162)? mem[5285] : 
                        (N164)? mem[5358] : 
                        (N166)? mem[5431] : 
                        (N168)? mem[5504] : 
                        (N170)? mem[5577] : 
                        (N172)? mem[5650] : 
                        (N174)? mem[5723] : 
                        (N176)? mem[5796] : 
                        (N178)? mem[5869] : 
                        (N180)? mem[5942] : 
                        (N182)? mem[6015] : 
                        (N184)? mem[6088] : 
                        (N186)? mem[6161] : 
                        (N188)? mem[6234] : 
                        (N190)? mem[6307] : 
                        (N192)? mem[6380] : 
                        (N194)? mem[6453] : 
                        (N196)? mem[6526] : 
                        (N198)? mem[6599] : 
                        (N200)? mem[6672] : 
                        (N202)? mem[6745] : 
                        (N204)? mem[6818] : 
                        (N206)? mem[6891] : 
                        (N208)? mem[6964] : 
                        (N210)? mem[7037] : 
                        (N212)? mem[7110] : 
                        (N214)? mem[7183] : 
                        (N216)? mem[7256] : 
                        (N218)? mem[7329] : 
                        (N220)? mem[7402] : 
                        (N222)? mem[7475] : 
                        (N224)? mem[7548] : 
                        (N226)? mem[7621] : 
                        (N228)? mem[7694] : 
                        (N230)? mem[7767] : 
                        (N232)? mem[7840] : 
                        (N234)? mem[7913] : 
                        (N236)? mem[7986] : 
                        (N238)? mem[8059] : 
                        (N240)? mem[8132] : 
                        (N242)? mem[8205] : 
                        (N244)? mem[8278] : 
                        (N246)? mem[8351] : 
                        (N248)? mem[8424] : 
                        (N250)? mem[8497] : 
                        (N252)? mem[8570] : 
                        (N254)? mem[8643] : 
                        (N256)? mem[8716] : 
                        (N258)? mem[8789] : 
                        (N260)? mem[8862] : 
                        (N262)? mem[8935] : 
                        (N264)? mem[9008] : 
                        (N266)? mem[9081] : 
                        (N268)? mem[9154] : 
                        (N270)? mem[9227] : 
                        (N272)? mem[9300] : 1'b0;
  assign r_data_o[28] = (N145)? mem[28] : 
                        (N147)? mem[101] : 
                        (N149)? mem[174] : 
                        (N151)? mem[247] : 
                        (N153)? mem[320] : 
                        (N155)? mem[393] : 
                        (N157)? mem[466] : 
                        (N159)? mem[539] : 
                        (N161)? mem[612] : 
                        (N163)? mem[685] : 
                        (N165)? mem[758] : 
                        (N167)? mem[831] : 
                        (N169)? mem[904] : 
                        (N171)? mem[977] : 
                        (N173)? mem[1050] : 
                        (N175)? mem[1123] : 
                        (N177)? mem[1196] : 
                        (N179)? mem[1269] : 
                        (N181)? mem[1342] : 
                        (N183)? mem[1415] : 
                        (N185)? mem[1488] : 
                        (N187)? mem[1561] : 
                        (N189)? mem[1634] : 
                        (N191)? mem[1707] : 
                        (N193)? mem[1780] : 
                        (N195)? mem[1853] : 
                        (N197)? mem[1926] : 
                        (N199)? mem[1999] : 
                        (N201)? mem[2072] : 
                        (N203)? mem[2145] : 
                        (N205)? mem[2218] : 
                        (N207)? mem[2291] : 
                        (N209)? mem[2364] : 
                        (N211)? mem[2437] : 
                        (N213)? mem[2510] : 
                        (N215)? mem[2583] : 
                        (N217)? mem[2656] : 
                        (N219)? mem[2729] : 
                        (N221)? mem[2802] : 
                        (N223)? mem[2875] : 
                        (N225)? mem[2948] : 
                        (N227)? mem[3021] : 
                        (N229)? mem[3094] : 
                        (N231)? mem[3167] : 
                        (N233)? mem[3240] : 
                        (N235)? mem[3313] : 
                        (N237)? mem[3386] : 
                        (N239)? mem[3459] : 
                        (N241)? mem[3532] : 
                        (N243)? mem[3605] : 
                        (N245)? mem[3678] : 
                        (N247)? mem[3751] : 
                        (N249)? mem[3824] : 
                        (N251)? mem[3897] : 
                        (N253)? mem[3970] : 
                        (N255)? mem[4043] : 
                        (N257)? mem[4116] : 
                        (N259)? mem[4189] : 
                        (N261)? mem[4262] : 
                        (N263)? mem[4335] : 
                        (N265)? mem[4408] : 
                        (N267)? mem[4481] : 
                        (N269)? mem[4554] : 
                        (N271)? mem[4627] : 
                        (N146)? mem[4700] : 
                        (N148)? mem[4773] : 
                        (N150)? mem[4846] : 
                        (N152)? mem[4919] : 
                        (N154)? mem[4992] : 
                        (N156)? mem[5065] : 
                        (N158)? mem[5138] : 
                        (N160)? mem[5211] : 
                        (N162)? mem[5284] : 
                        (N164)? mem[5357] : 
                        (N166)? mem[5430] : 
                        (N168)? mem[5503] : 
                        (N170)? mem[5576] : 
                        (N172)? mem[5649] : 
                        (N174)? mem[5722] : 
                        (N176)? mem[5795] : 
                        (N178)? mem[5868] : 
                        (N180)? mem[5941] : 
                        (N182)? mem[6014] : 
                        (N184)? mem[6087] : 
                        (N186)? mem[6160] : 
                        (N188)? mem[6233] : 
                        (N190)? mem[6306] : 
                        (N192)? mem[6379] : 
                        (N194)? mem[6452] : 
                        (N196)? mem[6525] : 
                        (N198)? mem[6598] : 
                        (N200)? mem[6671] : 
                        (N202)? mem[6744] : 
                        (N204)? mem[6817] : 
                        (N206)? mem[6890] : 
                        (N208)? mem[6963] : 
                        (N210)? mem[7036] : 
                        (N212)? mem[7109] : 
                        (N214)? mem[7182] : 
                        (N216)? mem[7255] : 
                        (N218)? mem[7328] : 
                        (N220)? mem[7401] : 
                        (N222)? mem[7474] : 
                        (N224)? mem[7547] : 
                        (N226)? mem[7620] : 
                        (N228)? mem[7693] : 
                        (N230)? mem[7766] : 
                        (N232)? mem[7839] : 
                        (N234)? mem[7912] : 
                        (N236)? mem[7985] : 
                        (N238)? mem[8058] : 
                        (N240)? mem[8131] : 
                        (N242)? mem[8204] : 
                        (N244)? mem[8277] : 
                        (N246)? mem[8350] : 
                        (N248)? mem[8423] : 
                        (N250)? mem[8496] : 
                        (N252)? mem[8569] : 
                        (N254)? mem[8642] : 
                        (N256)? mem[8715] : 
                        (N258)? mem[8788] : 
                        (N260)? mem[8861] : 
                        (N262)? mem[8934] : 
                        (N264)? mem[9007] : 
                        (N266)? mem[9080] : 
                        (N268)? mem[9153] : 
                        (N270)? mem[9226] : 
                        (N272)? mem[9299] : 1'b0;
  assign r_data_o[27] = (N145)? mem[27] : 
                        (N147)? mem[100] : 
                        (N149)? mem[173] : 
                        (N151)? mem[246] : 
                        (N153)? mem[319] : 
                        (N155)? mem[392] : 
                        (N157)? mem[465] : 
                        (N159)? mem[538] : 
                        (N161)? mem[611] : 
                        (N163)? mem[684] : 
                        (N165)? mem[757] : 
                        (N167)? mem[830] : 
                        (N169)? mem[903] : 
                        (N171)? mem[976] : 
                        (N173)? mem[1049] : 
                        (N175)? mem[1122] : 
                        (N177)? mem[1195] : 
                        (N179)? mem[1268] : 
                        (N181)? mem[1341] : 
                        (N183)? mem[1414] : 
                        (N185)? mem[1487] : 
                        (N187)? mem[1560] : 
                        (N189)? mem[1633] : 
                        (N191)? mem[1706] : 
                        (N193)? mem[1779] : 
                        (N195)? mem[1852] : 
                        (N197)? mem[1925] : 
                        (N199)? mem[1998] : 
                        (N201)? mem[2071] : 
                        (N203)? mem[2144] : 
                        (N205)? mem[2217] : 
                        (N207)? mem[2290] : 
                        (N209)? mem[2363] : 
                        (N211)? mem[2436] : 
                        (N213)? mem[2509] : 
                        (N215)? mem[2582] : 
                        (N217)? mem[2655] : 
                        (N219)? mem[2728] : 
                        (N221)? mem[2801] : 
                        (N223)? mem[2874] : 
                        (N225)? mem[2947] : 
                        (N227)? mem[3020] : 
                        (N229)? mem[3093] : 
                        (N231)? mem[3166] : 
                        (N233)? mem[3239] : 
                        (N235)? mem[3312] : 
                        (N237)? mem[3385] : 
                        (N239)? mem[3458] : 
                        (N241)? mem[3531] : 
                        (N243)? mem[3604] : 
                        (N245)? mem[3677] : 
                        (N247)? mem[3750] : 
                        (N249)? mem[3823] : 
                        (N251)? mem[3896] : 
                        (N253)? mem[3969] : 
                        (N255)? mem[4042] : 
                        (N257)? mem[4115] : 
                        (N259)? mem[4188] : 
                        (N261)? mem[4261] : 
                        (N263)? mem[4334] : 
                        (N265)? mem[4407] : 
                        (N267)? mem[4480] : 
                        (N269)? mem[4553] : 
                        (N271)? mem[4626] : 
                        (N146)? mem[4699] : 
                        (N148)? mem[4772] : 
                        (N150)? mem[4845] : 
                        (N152)? mem[4918] : 
                        (N154)? mem[4991] : 
                        (N156)? mem[5064] : 
                        (N158)? mem[5137] : 
                        (N160)? mem[5210] : 
                        (N162)? mem[5283] : 
                        (N164)? mem[5356] : 
                        (N166)? mem[5429] : 
                        (N168)? mem[5502] : 
                        (N170)? mem[5575] : 
                        (N172)? mem[5648] : 
                        (N174)? mem[5721] : 
                        (N176)? mem[5794] : 
                        (N178)? mem[5867] : 
                        (N180)? mem[5940] : 
                        (N182)? mem[6013] : 
                        (N184)? mem[6086] : 
                        (N186)? mem[6159] : 
                        (N188)? mem[6232] : 
                        (N190)? mem[6305] : 
                        (N192)? mem[6378] : 
                        (N194)? mem[6451] : 
                        (N196)? mem[6524] : 
                        (N198)? mem[6597] : 
                        (N200)? mem[6670] : 
                        (N202)? mem[6743] : 
                        (N204)? mem[6816] : 
                        (N206)? mem[6889] : 
                        (N208)? mem[6962] : 
                        (N210)? mem[7035] : 
                        (N212)? mem[7108] : 
                        (N214)? mem[7181] : 
                        (N216)? mem[7254] : 
                        (N218)? mem[7327] : 
                        (N220)? mem[7400] : 
                        (N222)? mem[7473] : 
                        (N224)? mem[7546] : 
                        (N226)? mem[7619] : 
                        (N228)? mem[7692] : 
                        (N230)? mem[7765] : 
                        (N232)? mem[7838] : 
                        (N234)? mem[7911] : 
                        (N236)? mem[7984] : 
                        (N238)? mem[8057] : 
                        (N240)? mem[8130] : 
                        (N242)? mem[8203] : 
                        (N244)? mem[8276] : 
                        (N246)? mem[8349] : 
                        (N248)? mem[8422] : 
                        (N250)? mem[8495] : 
                        (N252)? mem[8568] : 
                        (N254)? mem[8641] : 
                        (N256)? mem[8714] : 
                        (N258)? mem[8787] : 
                        (N260)? mem[8860] : 
                        (N262)? mem[8933] : 
                        (N264)? mem[9006] : 
                        (N266)? mem[9079] : 
                        (N268)? mem[9152] : 
                        (N270)? mem[9225] : 
                        (N272)? mem[9298] : 1'b0;
  assign r_data_o[26] = (N145)? mem[26] : 
                        (N147)? mem[99] : 
                        (N149)? mem[172] : 
                        (N151)? mem[245] : 
                        (N153)? mem[318] : 
                        (N155)? mem[391] : 
                        (N157)? mem[464] : 
                        (N159)? mem[537] : 
                        (N161)? mem[610] : 
                        (N163)? mem[683] : 
                        (N165)? mem[756] : 
                        (N167)? mem[829] : 
                        (N169)? mem[902] : 
                        (N171)? mem[975] : 
                        (N173)? mem[1048] : 
                        (N175)? mem[1121] : 
                        (N177)? mem[1194] : 
                        (N179)? mem[1267] : 
                        (N181)? mem[1340] : 
                        (N183)? mem[1413] : 
                        (N185)? mem[1486] : 
                        (N187)? mem[1559] : 
                        (N189)? mem[1632] : 
                        (N191)? mem[1705] : 
                        (N193)? mem[1778] : 
                        (N195)? mem[1851] : 
                        (N197)? mem[1924] : 
                        (N199)? mem[1997] : 
                        (N201)? mem[2070] : 
                        (N203)? mem[2143] : 
                        (N205)? mem[2216] : 
                        (N207)? mem[2289] : 
                        (N209)? mem[2362] : 
                        (N211)? mem[2435] : 
                        (N213)? mem[2508] : 
                        (N215)? mem[2581] : 
                        (N217)? mem[2654] : 
                        (N219)? mem[2727] : 
                        (N221)? mem[2800] : 
                        (N223)? mem[2873] : 
                        (N225)? mem[2946] : 
                        (N227)? mem[3019] : 
                        (N229)? mem[3092] : 
                        (N231)? mem[3165] : 
                        (N233)? mem[3238] : 
                        (N235)? mem[3311] : 
                        (N237)? mem[3384] : 
                        (N239)? mem[3457] : 
                        (N241)? mem[3530] : 
                        (N243)? mem[3603] : 
                        (N245)? mem[3676] : 
                        (N247)? mem[3749] : 
                        (N249)? mem[3822] : 
                        (N251)? mem[3895] : 
                        (N253)? mem[3968] : 
                        (N255)? mem[4041] : 
                        (N257)? mem[4114] : 
                        (N259)? mem[4187] : 
                        (N261)? mem[4260] : 
                        (N263)? mem[4333] : 
                        (N265)? mem[4406] : 
                        (N267)? mem[4479] : 
                        (N269)? mem[4552] : 
                        (N271)? mem[4625] : 
                        (N146)? mem[4698] : 
                        (N148)? mem[4771] : 
                        (N150)? mem[4844] : 
                        (N152)? mem[4917] : 
                        (N154)? mem[4990] : 
                        (N156)? mem[5063] : 
                        (N158)? mem[5136] : 
                        (N160)? mem[5209] : 
                        (N162)? mem[5282] : 
                        (N164)? mem[5355] : 
                        (N166)? mem[5428] : 
                        (N168)? mem[5501] : 
                        (N170)? mem[5574] : 
                        (N172)? mem[5647] : 
                        (N174)? mem[5720] : 
                        (N176)? mem[5793] : 
                        (N178)? mem[5866] : 
                        (N180)? mem[5939] : 
                        (N182)? mem[6012] : 
                        (N184)? mem[6085] : 
                        (N186)? mem[6158] : 
                        (N188)? mem[6231] : 
                        (N190)? mem[6304] : 
                        (N192)? mem[6377] : 
                        (N194)? mem[6450] : 
                        (N196)? mem[6523] : 
                        (N198)? mem[6596] : 
                        (N200)? mem[6669] : 
                        (N202)? mem[6742] : 
                        (N204)? mem[6815] : 
                        (N206)? mem[6888] : 
                        (N208)? mem[6961] : 
                        (N210)? mem[7034] : 
                        (N212)? mem[7107] : 
                        (N214)? mem[7180] : 
                        (N216)? mem[7253] : 
                        (N218)? mem[7326] : 
                        (N220)? mem[7399] : 
                        (N222)? mem[7472] : 
                        (N224)? mem[7545] : 
                        (N226)? mem[7618] : 
                        (N228)? mem[7691] : 
                        (N230)? mem[7764] : 
                        (N232)? mem[7837] : 
                        (N234)? mem[7910] : 
                        (N236)? mem[7983] : 
                        (N238)? mem[8056] : 
                        (N240)? mem[8129] : 
                        (N242)? mem[8202] : 
                        (N244)? mem[8275] : 
                        (N246)? mem[8348] : 
                        (N248)? mem[8421] : 
                        (N250)? mem[8494] : 
                        (N252)? mem[8567] : 
                        (N254)? mem[8640] : 
                        (N256)? mem[8713] : 
                        (N258)? mem[8786] : 
                        (N260)? mem[8859] : 
                        (N262)? mem[8932] : 
                        (N264)? mem[9005] : 
                        (N266)? mem[9078] : 
                        (N268)? mem[9151] : 
                        (N270)? mem[9224] : 
                        (N272)? mem[9297] : 1'b0;
  assign r_data_o[25] = (N145)? mem[25] : 
                        (N147)? mem[98] : 
                        (N149)? mem[171] : 
                        (N151)? mem[244] : 
                        (N153)? mem[317] : 
                        (N155)? mem[390] : 
                        (N157)? mem[463] : 
                        (N159)? mem[536] : 
                        (N161)? mem[609] : 
                        (N163)? mem[682] : 
                        (N165)? mem[755] : 
                        (N167)? mem[828] : 
                        (N169)? mem[901] : 
                        (N171)? mem[974] : 
                        (N173)? mem[1047] : 
                        (N175)? mem[1120] : 
                        (N177)? mem[1193] : 
                        (N179)? mem[1266] : 
                        (N181)? mem[1339] : 
                        (N183)? mem[1412] : 
                        (N185)? mem[1485] : 
                        (N187)? mem[1558] : 
                        (N189)? mem[1631] : 
                        (N191)? mem[1704] : 
                        (N193)? mem[1777] : 
                        (N195)? mem[1850] : 
                        (N197)? mem[1923] : 
                        (N199)? mem[1996] : 
                        (N201)? mem[2069] : 
                        (N203)? mem[2142] : 
                        (N205)? mem[2215] : 
                        (N207)? mem[2288] : 
                        (N209)? mem[2361] : 
                        (N211)? mem[2434] : 
                        (N213)? mem[2507] : 
                        (N215)? mem[2580] : 
                        (N217)? mem[2653] : 
                        (N219)? mem[2726] : 
                        (N221)? mem[2799] : 
                        (N223)? mem[2872] : 
                        (N225)? mem[2945] : 
                        (N227)? mem[3018] : 
                        (N229)? mem[3091] : 
                        (N231)? mem[3164] : 
                        (N233)? mem[3237] : 
                        (N235)? mem[3310] : 
                        (N237)? mem[3383] : 
                        (N239)? mem[3456] : 
                        (N241)? mem[3529] : 
                        (N243)? mem[3602] : 
                        (N245)? mem[3675] : 
                        (N247)? mem[3748] : 
                        (N249)? mem[3821] : 
                        (N251)? mem[3894] : 
                        (N253)? mem[3967] : 
                        (N255)? mem[4040] : 
                        (N257)? mem[4113] : 
                        (N259)? mem[4186] : 
                        (N261)? mem[4259] : 
                        (N263)? mem[4332] : 
                        (N265)? mem[4405] : 
                        (N267)? mem[4478] : 
                        (N269)? mem[4551] : 
                        (N271)? mem[4624] : 
                        (N146)? mem[4697] : 
                        (N148)? mem[4770] : 
                        (N150)? mem[4843] : 
                        (N152)? mem[4916] : 
                        (N154)? mem[4989] : 
                        (N156)? mem[5062] : 
                        (N158)? mem[5135] : 
                        (N160)? mem[5208] : 
                        (N162)? mem[5281] : 
                        (N164)? mem[5354] : 
                        (N166)? mem[5427] : 
                        (N168)? mem[5500] : 
                        (N170)? mem[5573] : 
                        (N172)? mem[5646] : 
                        (N174)? mem[5719] : 
                        (N176)? mem[5792] : 
                        (N178)? mem[5865] : 
                        (N180)? mem[5938] : 
                        (N182)? mem[6011] : 
                        (N184)? mem[6084] : 
                        (N186)? mem[6157] : 
                        (N188)? mem[6230] : 
                        (N190)? mem[6303] : 
                        (N192)? mem[6376] : 
                        (N194)? mem[6449] : 
                        (N196)? mem[6522] : 
                        (N198)? mem[6595] : 
                        (N200)? mem[6668] : 
                        (N202)? mem[6741] : 
                        (N204)? mem[6814] : 
                        (N206)? mem[6887] : 
                        (N208)? mem[6960] : 
                        (N210)? mem[7033] : 
                        (N212)? mem[7106] : 
                        (N214)? mem[7179] : 
                        (N216)? mem[7252] : 
                        (N218)? mem[7325] : 
                        (N220)? mem[7398] : 
                        (N222)? mem[7471] : 
                        (N224)? mem[7544] : 
                        (N226)? mem[7617] : 
                        (N228)? mem[7690] : 
                        (N230)? mem[7763] : 
                        (N232)? mem[7836] : 
                        (N234)? mem[7909] : 
                        (N236)? mem[7982] : 
                        (N238)? mem[8055] : 
                        (N240)? mem[8128] : 
                        (N242)? mem[8201] : 
                        (N244)? mem[8274] : 
                        (N246)? mem[8347] : 
                        (N248)? mem[8420] : 
                        (N250)? mem[8493] : 
                        (N252)? mem[8566] : 
                        (N254)? mem[8639] : 
                        (N256)? mem[8712] : 
                        (N258)? mem[8785] : 
                        (N260)? mem[8858] : 
                        (N262)? mem[8931] : 
                        (N264)? mem[9004] : 
                        (N266)? mem[9077] : 
                        (N268)? mem[9150] : 
                        (N270)? mem[9223] : 
                        (N272)? mem[9296] : 1'b0;
  assign r_data_o[24] = (N145)? mem[24] : 
                        (N147)? mem[97] : 
                        (N149)? mem[170] : 
                        (N151)? mem[243] : 
                        (N153)? mem[316] : 
                        (N155)? mem[389] : 
                        (N157)? mem[462] : 
                        (N159)? mem[535] : 
                        (N161)? mem[608] : 
                        (N163)? mem[681] : 
                        (N165)? mem[754] : 
                        (N167)? mem[827] : 
                        (N169)? mem[900] : 
                        (N171)? mem[973] : 
                        (N173)? mem[1046] : 
                        (N175)? mem[1119] : 
                        (N177)? mem[1192] : 
                        (N179)? mem[1265] : 
                        (N181)? mem[1338] : 
                        (N183)? mem[1411] : 
                        (N185)? mem[1484] : 
                        (N187)? mem[1557] : 
                        (N189)? mem[1630] : 
                        (N191)? mem[1703] : 
                        (N193)? mem[1776] : 
                        (N195)? mem[1849] : 
                        (N197)? mem[1922] : 
                        (N199)? mem[1995] : 
                        (N201)? mem[2068] : 
                        (N203)? mem[2141] : 
                        (N205)? mem[2214] : 
                        (N207)? mem[2287] : 
                        (N209)? mem[2360] : 
                        (N211)? mem[2433] : 
                        (N213)? mem[2506] : 
                        (N215)? mem[2579] : 
                        (N217)? mem[2652] : 
                        (N219)? mem[2725] : 
                        (N221)? mem[2798] : 
                        (N223)? mem[2871] : 
                        (N225)? mem[2944] : 
                        (N227)? mem[3017] : 
                        (N229)? mem[3090] : 
                        (N231)? mem[3163] : 
                        (N233)? mem[3236] : 
                        (N235)? mem[3309] : 
                        (N237)? mem[3382] : 
                        (N239)? mem[3455] : 
                        (N241)? mem[3528] : 
                        (N243)? mem[3601] : 
                        (N245)? mem[3674] : 
                        (N247)? mem[3747] : 
                        (N249)? mem[3820] : 
                        (N251)? mem[3893] : 
                        (N253)? mem[3966] : 
                        (N255)? mem[4039] : 
                        (N257)? mem[4112] : 
                        (N259)? mem[4185] : 
                        (N261)? mem[4258] : 
                        (N263)? mem[4331] : 
                        (N265)? mem[4404] : 
                        (N267)? mem[4477] : 
                        (N269)? mem[4550] : 
                        (N271)? mem[4623] : 
                        (N146)? mem[4696] : 
                        (N148)? mem[4769] : 
                        (N150)? mem[4842] : 
                        (N152)? mem[4915] : 
                        (N154)? mem[4988] : 
                        (N156)? mem[5061] : 
                        (N158)? mem[5134] : 
                        (N160)? mem[5207] : 
                        (N162)? mem[5280] : 
                        (N164)? mem[5353] : 
                        (N166)? mem[5426] : 
                        (N168)? mem[5499] : 
                        (N170)? mem[5572] : 
                        (N172)? mem[5645] : 
                        (N174)? mem[5718] : 
                        (N176)? mem[5791] : 
                        (N178)? mem[5864] : 
                        (N180)? mem[5937] : 
                        (N182)? mem[6010] : 
                        (N184)? mem[6083] : 
                        (N186)? mem[6156] : 
                        (N188)? mem[6229] : 
                        (N190)? mem[6302] : 
                        (N192)? mem[6375] : 
                        (N194)? mem[6448] : 
                        (N196)? mem[6521] : 
                        (N198)? mem[6594] : 
                        (N200)? mem[6667] : 
                        (N202)? mem[6740] : 
                        (N204)? mem[6813] : 
                        (N206)? mem[6886] : 
                        (N208)? mem[6959] : 
                        (N210)? mem[7032] : 
                        (N212)? mem[7105] : 
                        (N214)? mem[7178] : 
                        (N216)? mem[7251] : 
                        (N218)? mem[7324] : 
                        (N220)? mem[7397] : 
                        (N222)? mem[7470] : 
                        (N224)? mem[7543] : 
                        (N226)? mem[7616] : 
                        (N228)? mem[7689] : 
                        (N230)? mem[7762] : 
                        (N232)? mem[7835] : 
                        (N234)? mem[7908] : 
                        (N236)? mem[7981] : 
                        (N238)? mem[8054] : 
                        (N240)? mem[8127] : 
                        (N242)? mem[8200] : 
                        (N244)? mem[8273] : 
                        (N246)? mem[8346] : 
                        (N248)? mem[8419] : 
                        (N250)? mem[8492] : 
                        (N252)? mem[8565] : 
                        (N254)? mem[8638] : 
                        (N256)? mem[8711] : 
                        (N258)? mem[8784] : 
                        (N260)? mem[8857] : 
                        (N262)? mem[8930] : 
                        (N264)? mem[9003] : 
                        (N266)? mem[9076] : 
                        (N268)? mem[9149] : 
                        (N270)? mem[9222] : 
                        (N272)? mem[9295] : 1'b0;
  assign r_data_o[23] = (N145)? mem[23] : 
                        (N147)? mem[96] : 
                        (N149)? mem[169] : 
                        (N151)? mem[242] : 
                        (N153)? mem[315] : 
                        (N155)? mem[388] : 
                        (N157)? mem[461] : 
                        (N159)? mem[534] : 
                        (N161)? mem[607] : 
                        (N163)? mem[680] : 
                        (N165)? mem[753] : 
                        (N167)? mem[826] : 
                        (N169)? mem[899] : 
                        (N171)? mem[972] : 
                        (N173)? mem[1045] : 
                        (N175)? mem[1118] : 
                        (N177)? mem[1191] : 
                        (N179)? mem[1264] : 
                        (N181)? mem[1337] : 
                        (N183)? mem[1410] : 
                        (N185)? mem[1483] : 
                        (N187)? mem[1556] : 
                        (N189)? mem[1629] : 
                        (N191)? mem[1702] : 
                        (N193)? mem[1775] : 
                        (N195)? mem[1848] : 
                        (N197)? mem[1921] : 
                        (N199)? mem[1994] : 
                        (N201)? mem[2067] : 
                        (N203)? mem[2140] : 
                        (N205)? mem[2213] : 
                        (N207)? mem[2286] : 
                        (N209)? mem[2359] : 
                        (N211)? mem[2432] : 
                        (N213)? mem[2505] : 
                        (N215)? mem[2578] : 
                        (N217)? mem[2651] : 
                        (N219)? mem[2724] : 
                        (N221)? mem[2797] : 
                        (N223)? mem[2870] : 
                        (N225)? mem[2943] : 
                        (N227)? mem[3016] : 
                        (N229)? mem[3089] : 
                        (N231)? mem[3162] : 
                        (N233)? mem[3235] : 
                        (N235)? mem[3308] : 
                        (N237)? mem[3381] : 
                        (N239)? mem[3454] : 
                        (N241)? mem[3527] : 
                        (N243)? mem[3600] : 
                        (N245)? mem[3673] : 
                        (N247)? mem[3746] : 
                        (N249)? mem[3819] : 
                        (N251)? mem[3892] : 
                        (N253)? mem[3965] : 
                        (N255)? mem[4038] : 
                        (N257)? mem[4111] : 
                        (N259)? mem[4184] : 
                        (N261)? mem[4257] : 
                        (N263)? mem[4330] : 
                        (N265)? mem[4403] : 
                        (N267)? mem[4476] : 
                        (N269)? mem[4549] : 
                        (N271)? mem[4622] : 
                        (N146)? mem[4695] : 
                        (N148)? mem[4768] : 
                        (N150)? mem[4841] : 
                        (N152)? mem[4914] : 
                        (N154)? mem[4987] : 
                        (N156)? mem[5060] : 
                        (N158)? mem[5133] : 
                        (N160)? mem[5206] : 
                        (N162)? mem[5279] : 
                        (N164)? mem[5352] : 
                        (N166)? mem[5425] : 
                        (N168)? mem[5498] : 
                        (N170)? mem[5571] : 
                        (N172)? mem[5644] : 
                        (N174)? mem[5717] : 
                        (N176)? mem[5790] : 
                        (N178)? mem[5863] : 
                        (N180)? mem[5936] : 
                        (N182)? mem[6009] : 
                        (N184)? mem[6082] : 
                        (N186)? mem[6155] : 
                        (N188)? mem[6228] : 
                        (N190)? mem[6301] : 
                        (N192)? mem[6374] : 
                        (N194)? mem[6447] : 
                        (N196)? mem[6520] : 
                        (N198)? mem[6593] : 
                        (N200)? mem[6666] : 
                        (N202)? mem[6739] : 
                        (N204)? mem[6812] : 
                        (N206)? mem[6885] : 
                        (N208)? mem[6958] : 
                        (N210)? mem[7031] : 
                        (N212)? mem[7104] : 
                        (N214)? mem[7177] : 
                        (N216)? mem[7250] : 
                        (N218)? mem[7323] : 
                        (N220)? mem[7396] : 
                        (N222)? mem[7469] : 
                        (N224)? mem[7542] : 
                        (N226)? mem[7615] : 
                        (N228)? mem[7688] : 
                        (N230)? mem[7761] : 
                        (N232)? mem[7834] : 
                        (N234)? mem[7907] : 
                        (N236)? mem[7980] : 
                        (N238)? mem[8053] : 
                        (N240)? mem[8126] : 
                        (N242)? mem[8199] : 
                        (N244)? mem[8272] : 
                        (N246)? mem[8345] : 
                        (N248)? mem[8418] : 
                        (N250)? mem[8491] : 
                        (N252)? mem[8564] : 
                        (N254)? mem[8637] : 
                        (N256)? mem[8710] : 
                        (N258)? mem[8783] : 
                        (N260)? mem[8856] : 
                        (N262)? mem[8929] : 
                        (N264)? mem[9002] : 
                        (N266)? mem[9075] : 
                        (N268)? mem[9148] : 
                        (N270)? mem[9221] : 
                        (N272)? mem[9294] : 1'b0;
  assign r_data_o[22] = (N145)? mem[22] : 
                        (N147)? mem[95] : 
                        (N149)? mem[168] : 
                        (N151)? mem[241] : 
                        (N153)? mem[314] : 
                        (N155)? mem[387] : 
                        (N157)? mem[460] : 
                        (N159)? mem[533] : 
                        (N161)? mem[606] : 
                        (N163)? mem[679] : 
                        (N165)? mem[752] : 
                        (N167)? mem[825] : 
                        (N169)? mem[898] : 
                        (N171)? mem[971] : 
                        (N173)? mem[1044] : 
                        (N175)? mem[1117] : 
                        (N177)? mem[1190] : 
                        (N179)? mem[1263] : 
                        (N181)? mem[1336] : 
                        (N183)? mem[1409] : 
                        (N185)? mem[1482] : 
                        (N187)? mem[1555] : 
                        (N189)? mem[1628] : 
                        (N191)? mem[1701] : 
                        (N193)? mem[1774] : 
                        (N195)? mem[1847] : 
                        (N197)? mem[1920] : 
                        (N199)? mem[1993] : 
                        (N201)? mem[2066] : 
                        (N203)? mem[2139] : 
                        (N205)? mem[2212] : 
                        (N207)? mem[2285] : 
                        (N209)? mem[2358] : 
                        (N211)? mem[2431] : 
                        (N213)? mem[2504] : 
                        (N215)? mem[2577] : 
                        (N217)? mem[2650] : 
                        (N219)? mem[2723] : 
                        (N221)? mem[2796] : 
                        (N223)? mem[2869] : 
                        (N225)? mem[2942] : 
                        (N227)? mem[3015] : 
                        (N229)? mem[3088] : 
                        (N231)? mem[3161] : 
                        (N233)? mem[3234] : 
                        (N235)? mem[3307] : 
                        (N237)? mem[3380] : 
                        (N239)? mem[3453] : 
                        (N241)? mem[3526] : 
                        (N243)? mem[3599] : 
                        (N245)? mem[3672] : 
                        (N247)? mem[3745] : 
                        (N249)? mem[3818] : 
                        (N251)? mem[3891] : 
                        (N253)? mem[3964] : 
                        (N255)? mem[4037] : 
                        (N257)? mem[4110] : 
                        (N259)? mem[4183] : 
                        (N261)? mem[4256] : 
                        (N263)? mem[4329] : 
                        (N265)? mem[4402] : 
                        (N267)? mem[4475] : 
                        (N269)? mem[4548] : 
                        (N271)? mem[4621] : 
                        (N146)? mem[4694] : 
                        (N148)? mem[4767] : 
                        (N150)? mem[4840] : 
                        (N152)? mem[4913] : 
                        (N154)? mem[4986] : 
                        (N156)? mem[5059] : 
                        (N158)? mem[5132] : 
                        (N160)? mem[5205] : 
                        (N162)? mem[5278] : 
                        (N164)? mem[5351] : 
                        (N166)? mem[5424] : 
                        (N168)? mem[5497] : 
                        (N170)? mem[5570] : 
                        (N172)? mem[5643] : 
                        (N174)? mem[5716] : 
                        (N176)? mem[5789] : 
                        (N178)? mem[5862] : 
                        (N180)? mem[5935] : 
                        (N182)? mem[6008] : 
                        (N184)? mem[6081] : 
                        (N186)? mem[6154] : 
                        (N188)? mem[6227] : 
                        (N190)? mem[6300] : 
                        (N192)? mem[6373] : 
                        (N194)? mem[6446] : 
                        (N196)? mem[6519] : 
                        (N198)? mem[6592] : 
                        (N200)? mem[6665] : 
                        (N202)? mem[6738] : 
                        (N204)? mem[6811] : 
                        (N206)? mem[6884] : 
                        (N208)? mem[6957] : 
                        (N210)? mem[7030] : 
                        (N212)? mem[7103] : 
                        (N214)? mem[7176] : 
                        (N216)? mem[7249] : 
                        (N218)? mem[7322] : 
                        (N220)? mem[7395] : 
                        (N222)? mem[7468] : 
                        (N224)? mem[7541] : 
                        (N226)? mem[7614] : 
                        (N228)? mem[7687] : 
                        (N230)? mem[7760] : 
                        (N232)? mem[7833] : 
                        (N234)? mem[7906] : 
                        (N236)? mem[7979] : 
                        (N238)? mem[8052] : 
                        (N240)? mem[8125] : 
                        (N242)? mem[8198] : 
                        (N244)? mem[8271] : 
                        (N246)? mem[8344] : 
                        (N248)? mem[8417] : 
                        (N250)? mem[8490] : 
                        (N252)? mem[8563] : 
                        (N254)? mem[8636] : 
                        (N256)? mem[8709] : 
                        (N258)? mem[8782] : 
                        (N260)? mem[8855] : 
                        (N262)? mem[8928] : 
                        (N264)? mem[9001] : 
                        (N266)? mem[9074] : 
                        (N268)? mem[9147] : 
                        (N270)? mem[9220] : 
                        (N272)? mem[9293] : 1'b0;
  assign r_data_o[21] = (N145)? mem[21] : 
                        (N147)? mem[94] : 
                        (N149)? mem[167] : 
                        (N151)? mem[240] : 
                        (N153)? mem[313] : 
                        (N155)? mem[386] : 
                        (N157)? mem[459] : 
                        (N159)? mem[532] : 
                        (N161)? mem[605] : 
                        (N163)? mem[678] : 
                        (N165)? mem[751] : 
                        (N167)? mem[824] : 
                        (N169)? mem[897] : 
                        (N171)? mem[970] : 
                        (N173)? mem[1043] : 
                        (N175)? mem[1116] : 
                        (N177)? mem[1189] : 
                        (N179)? mem[1262] : 
                        (N181)? mem[1335] : 
                        (N183)? mem[1408] : 
                        (N185)? mem[1481] : 
                        (N187)? mem[1554] : 
                        (N189)? mem[1627] : 
                        (N191)? mem[1700] : 
                        (N193)? mem[1773] : 
                        (N195)? mem[1846] : 
                        (N197)? mem[1919] : 
                        (N199)? mem[1992] : 
                        (N201)? mem[2065] : 
                        (N203)? mem[2138] : 
                        (N205)? mem[2211] : 
                        (N207)? mem[2284] : 
                        (N209)? mem[2357] : 
                        (N211)? mem[2430] : 
                        (N213)? mem[2503] : 
                        (N215)? mem[2576] : 
                        (N217)? mem[2649] : 
                        (N219)? mem[2722] : 
                        (N221)? mem[2795] : 
                        (N223)? mem[2868] : 
                        (N225)? mem[2941] : 
                        (N227)? mem[3014] : 
                        (N229)? mem[3087] : 
                        (N231)? mem[3160] : 
                        (N233)? mem[3233] : 
                        (N235)? mem[3306] : 
                        (N237)? mem[3379] : 
                        (N239)? mem[3452] : 
                        (N241)? mem[3525] : 
                        (N243)? mem[3598] : 
                        (N245)? mem[3671] : 
                        (N247)? mem[3744] : 
                        (N249)? mem[3817] : 
                        (N251)? mem[3890] : 
                        (N253)? mem[3963] : 
                        (N255)? mem[4036] : 
                        (N257)? mem[4109] : 
                        (N259)? mem[4182] : 
                        (N261)? mem[4255] : 
                        (N263)? mem[4328] : 
                        (N265)? mem[4401] : 
                        (N267)? mem[4474] : 
                        (N269)? mem[4547] : 
                        (N271)? mem[4620] : 
                        (N146)? mem[4693] : 
                        (N148)? mem[4766] : 
                        (N150)? mem[4839] : 
                        (N152)? mem[4912] : 
                        (N154)? mem[4985] : 
                        (N156)? mem[5058] : 
                        (N158)? mem[5131] : 
                        (N160)? mem[5204] : 
                        (N162)? mem[5277] : 
                        (N164)? mem[5350] : 
                        (N166)? mem[5423] : 
                        (N168)? mem[5496] : 
                        (N170)? mem[5569] : 
                        (N172)? mem[5642] : 
                        (N174)? mem[5715] : 
                        (N176)? mem[5788] : 
                        (N178)? mem[5861] : 
                        (N180)? mem[5934] : 
                        (N182)? mem[6007] : 
                        (N184)? mem[6080] : 
                        (N186)? mem[6153] : 
                        (N188)? mem[6226] : 
                        (N190)? mem[6299] : 
                        (N192)? mem[6372] : 
                        (N194)? mem[6445] : 
                        (N196)? mem[6518] : 
                        (N198)? mem[6591] : 
                        (N200)? mem[6664] : 
                        (N202)? mem[6737] : 
                        (N204)? mem[6810] : 
                        (N206)? mem[6883] : 
                        (N208)? mem[6956] : 
                        (N210)? mem[7029] : 
                        (N212)? mem[7102] : 
                        (N214)? mem[7175] : 
                        (N216)? mem[7248] : 
                        (N218)? mem[7321] : 
                        (N220)? mem[7394] : 
                        (N222)? mem[7467] : 
                        (N224)? mem[7540] : 
                        (N226)? mem[7613] : 
                        (N228)? mem[7686] : 
                        (N230)? mem[7759] : 
                        (N232)? mem[7832] : 
                        (N234)? mem[7905] : 
                        (N236)? mem[7978] : 
                        (N238)? mem[8051] : 
                        (N240)? mem[8124] : 
                        (N242)? mem[8197] : 
                        (N244)? mem[8270] : 
                        (N246)? mem[8343] : 
                        (N248)? mem[8416] : 
                        (N250)? mem[8489] : 
                        (N252)? mem[8562] : 
                        (N254)? mem[8635] : 
                        (N256)? mem[8708] : 
                        (N258)? mem[8781] : 
                        (N260)? mem[8854] : 
                        (N262)? mem[8927] : 
                        (N264)? mem[9000] : 
                        (N266)? mem[9073] : 
                        (N268)? mem[9146] : 
                        (N270)? mem[9219] : 
                        (N272)? mem[9292] : 1'b0;
  assign r_data_o[20] = (N145)? mem[20] : 
                        (N147)? mem[93] : 
                        (N149)? mem[166] : 
                        (N151)? mem[239] : 
                        (N153)? mem[312] : 
                        (N155)? mem[385] : 
                        (N157)? mem[458] : 
                        (N159)? mem[531] : 
                        (N161)? mem[604] : 
                        (N163)? mem[677] : 
                        (N165)? mem[750] : 
                        (N167)? mem[823] : 
                        (N169)? mem[896] : 
                        (N171)? mem[969] : 
                        (N173)? mem[1042] : 
                        (N175)? mem[1115] : 
                        (N177)? mem[1188] : 
                        (N179)? mem[1261] : 
                        (N181)? mem[1334] : 
                        (N183)? mem[1407] : 
                        (N185)? mem[1480] : 
                        (N187)? mem[1553] : 
                        (N189)? mem[1626] : 
                        (N191)? mem[1699] : 
                        (N193)? mem[1772] : 
                        (N195)? mem[1845] : 
                        (N197)? mem[1918] : 
                        (N199)? mem[1991] : 
                        (N201)? mem[2064] : 
                        (N203)? mem[2137] : 
                        (N205)? mem[2210] : 
                        (N207)? mem[2283] : 
                        (N209)? mem[2356] : 
                        (N211)? mem[2429] : 
                        (N213)? mem[2502] : 
                        (N215)? mem[2575] : 
                        (N217)? mem[2648] : 
                        (N219)? mem[2721] : 
                        (N221)? mem[2794] : 
                        (N223)? mem[2867] : 
                        (N225)? mem[2940] : 
                        (N227)? mem[3013] : 
                        (N229)? mem[3086] : 
                        (N231)? mem[3159] : 
                        (N233)? mem[3232] : 
                        (N235)? mem[3305] : 
                        (N237)? mem[3378] : 
                        (N239)? mem[3451] : 
                        (N241)? mem[3524] : 
                        (N243)? mem[3597] : 
                        (N245)? mem[3670] : 
                        (N247)? mem[3743] : 
                        (N249)? mem[3816] : 
                        (N251)? mem[3889] : 
                        (N253)? mem[3962] : 
                        (N255)? mem[4035] : 
                        (N257)? mem[4108] : 
                        (N259)? mem[4181] : 
                        (N261)? mem[4254] : 
                        (N263)? mem[4327] : 
                        (N265)? mem[4400] : 
                        (N267)? mem[4473] : 
                        (N269)? mem[4546] : 
                        (N271)? mem[4619] : 
                        (N146)? mem[4692] : 
                        (N148)? mem[4765] : 
                        (N150)? mem[4838] : 
                        (N152)? mem[4911] : 
                        (N154)? mem[4984] : 
                        (N156)? mem[5057] : 
                        (N158)? mem[5130] : 
                        (N160)? mem[5203] : 
                        (N162)? mem[5276] : 
                        (N164)? mem[5349] : 
                        (N166)? mem[5422] : 
                        (N168)? mem[5495] : 
                        (N170)? mem[5568] : 
                        (N172)? mem[5641] : 
                        (N174)? mem[5714] : 
                        (N176)? mem[5787] : 
                        (N178)? mem[5860] : 
                        (N180)? mem[5933] : 
                        (N182)? mem[6006] : 
                        (N184)? mem[6079] : 
                        (N186)? mem[6152] : 
                        (N188)? mem[6225] : 
                        (N190)? mem[6298] : 
                        (N192)? mem[6371] : 
                        (N194)? mem[6444] : 
                        (N196)? mem[6517] : 
                        (N198)? mem[6590] : 
                        (N200)? mem[6663] : 
                        (N202)? mem[6736] : 
                        (N204)? mem[6809] : 
                        (N206)? mem[6882] : 
                        (N208)? mem[6955] : 
                        (N210)? mem[7028] : 
                        (N212)? mem[7101] : 
                        (N214)? mem[7174] : 
                        (N216)? mem[7247] : 
                        (N218)? mem[7320] : 
                        (N220)? mem[7393] : 
                        (N222)? mem[7466] : 
                        (N224)? mem[7539] : 
                        (N226)? mem[7612] : 
                        (N228)? mem[7685] : 
                        (N230)? mem[7758] : 
                        (N232)? mem[7831] : 
                        (N234)? mem[7904] : 
                        (N236)? mem[7977] : 
                        (N238)? mem[8050] : 
                        (N240)? mem[8123] : 
                        (N242)? mem[8196] : 
                        (N244)? mem[8269] : 
                        (N246)? mem[8342] : 
                        (N248)? mem[8415] : 
                        (N250)? mem[8488] : 
                        (N252)? mem[8561] : 
                        (N254)? mem[8634] : 
                        (N256)? mem[8707] : 
                        (N258)? mem[8780] : 
                        (N260)? mem[8853] : 
                        (N262)? mem[8926] : 
                        (N264)? mem[8999] : 
                        (N266)? mem[9072] : 
                        (N268)? mem[9145] : 
                        (N270)? mem[9218] : 
                        (N272)? mem[9291] : 1'b0;
  assign r_data_o[19] = (N145)? mem[19] : 
                        (N147)? mem[92] : 
                        (N149)? mem[165] : 
                        (N151)? mem[238] : 
                        (N153)? mem[311] : 
                        (N155)? mem[384] : 
                        (N157)? mem[457] : 
                        (N159)? mem[530] : 
                        (N161)? mem[603] : 
                        (N163)? mem[676] : 
                        (N165)? mem[749] : 
                        (N167)? mem[822] : 
                        (N169)? mem[895] : 
                        (N171)? mem[968] : 
                        (N173)? mem[1041] : 
                        (N175)? mem[1114] : 
                        (N177)? mem[1187] : 
                        (N179)? mem[1260] : 
                        (N181)? mem[1333] : 
                        (N183)? mem[1406] : 
                        (N185)? mem[1479] : 
                        (N187)? mem[1552] : 
                        (N189)? mem[1625] : 
                        (N191)? mem[1698] : 
                        (N193)? mem[1771] : 
                        (N195)? mem[1844] : 
                        (N197)? mem[1917] : 
                        (N199)? mem[1990] : 
                        (N201)? mem[2063] : 
                        (N203)? mem[2136] : 
                        (N205)? mem[2209] : 
                        (N207)? mem[2282] : 
                        (N209)? mem[2355] : 
                        (N211)? mem[2428] : 
                        (N213)? mem[2501] : 
                        (N215)? mem[2574] : 
                        (N217)? mem[2647] : 
                        (N219)? mem[2720] : 
                        (N221)? mem[2793] : 
                        (N223)? mem[2866] : 
                        (N225)? mem[2939] : 
                        (N227)? mem[3012] : 
                        (N229)? mem[3085] : 
                        (N231)? mem[3158] : 
                        (N233)? mem[3231] : 
                        (N235)? mem[3304] : 
                        (N237)? mem[3377] : 
                        (N239)? mem[3450] : 
                        (N241)? mem[3523] : 
                        (N243)? mem[3596] : 
                        (N245)? mem[3669] : 
                        (N247)? mem[3742] : 
                        (N249)? mem[3815] : 
                        (N251)? mem[3888] : 
                        (N253)? mem[3961] : 
                        (N255)? mem[4034] : 
                        (N257)? mem[4107] : 
                        (N259)? mem[4180] : 
                        (N261)? mem[4253] : 
                        (N263)? mem[4326] : 
                        (N265)? mem[4399] : 
                        (N267)? mem[4472] : 
                        (N269)? mem[4545] : 
                        (N271)? mem[4618] : 
                        (N146)? mem[4691] : 
                        (N148)? mem[4764] : 
                        (N150)? mem[4837] : 
                        (N152)? mem[4910] : 
                        (N154)? mem[4983] : 
                        (N156)? mem[5056] : 
                        (N158)? mem[5129] : 
                        (N160)? mem[5202] : 
                        (N162)? mem[5275] : 
                        (N164)? mem[5348] : 
                        (N166)? mem[5421] : 
                        (N168)? mem[5494] : 
                        (N170)? mem[5567] : 
                        (N172)? mem[5640] : 
                        (N174)? mem[5713] : 
                        (N176)? mem[5786] : 
                        (N178)? mem[5859] : 
                        (N180)? mem[5932] : 
                        (N182)? mem[6005] : 
                        (N184)? mem[6078] : 
                        (N186)? mem[6151] : 
                        (N188)? mem[6224] : 
                        (N190)? mem[6297] : 
                        (N192)? mem[6370] : 
                        (N194)? mem[6443] : 
                        (N196)? mem[6516] : 
                        (N198)? mem[6589] : 
                        (N200)? mem[6662] : 
                        (N202)? mem[6735] : 
                        (N204)? mem[6808] : 
                        (N206)? mem[6881] : 
                        (N208)? mem[6954] : 
                        (N210)? mem[7027] : 
                        (N212)? mem[7100] : 
                        (N214)? mem[7173] : 
                        (N216)? mem[7246] : 
                        (N218)? mem[7319] : 
                        (N220)? mem[7392] : 
                        (N222)? mem[7465] : 
                        (N224)? mem[7538] : 
                        (N226)? mem[7611] : 
                        (N228)? mem[7684] : 
                        (N230)? mem[7757] : 
                        (N232)? mem[7830] : 
                        (N234)? mem[7903] : 
                        (N236)? mem[7976] : 
                        (N238)? mem[8049] : 
                        (N240)? mem[8122] : 
                        (N242)? mem[8195] : 
                        (N244)? mem[8268] : 
                        (N246)? mem[8341] : 
                        (N248)? mem[8414] : 
                        (N250)? mem[8487] : 
                        (N252)? mem[8560] : 
                        (N254)? mem[8633] : 
                        (N256)? mem[8706] : 
                        (N258)? mem[8779] : 
                        (N260)? mem[8852] : 
                        (N262)? mem[8925] : 
                        (N264)? mem[8998] : 
                        (N266)? mem[9071] : 
                        (N268)? mem[9144] : 
                        (N270)? mem[9217] : 
                        (N272)? mem[9290] : 1'b0;
  assign r_data_o[18] = (N145)? mem[18] : 
                        (N147)? mem[91] : 
                        (N149)? mem[164] : 
                        (N151)? mem[237] : 
                        (N153)? mem[310] : 
                        (N155)? mem[383] : 
                        (N157)? mem[456] : 
                        (N159)? mem[529] : 
                        (N161)? mem[602] : 
                        (N163)? mem[675] : 
                        (N165)? mem[748] : 
                        (N167)? mem[821] : 
                        (N169)? mem[894] : 
                        (N171)? mem[967] : 
                        (N173)? mem[1040] : 
                        (N175)? mem[1113] : 
                        (N177)? mem[1186] : 
                        (N179)? mem[1259] : 
                        (N181)? mem[1332] : 
                        (N183)? mem[1405] : 
                        (N185)? mem[1478] : 
                        (N187)? mem[1551] : 
                        (N189)? mem[1624] : 
                        (N191)? mem[1697] : 
                        (N193)? mem[1770] : 
                        (N195)? mem[1843] : 
                        (N197)? mem[1916] : 
                        (N199)? mem[1989] : 
                        (N201)? mem[2062] : 
                        (N203)? mem[2135] : 
                        (N205)? mem[2208] : 
                        (N207)? mem[2281] : 
                        (N209)? mem[2354] : 
                        (N211)? mem[2427] : 
                        (N213)? mem[2500] : 
                        (N215)? mem[2573] : 
                        (N217)? mem[2646] : 
                        (N219)? mem[2719] : 
                        (N221)? mem[2792] : 
                        (N223)? mem[2865] : 
                        (N225)? mem[2938] : 
                        (N227)? mem[3011] : 
                        (N229)? mem[3084] : 
                        (N231)? mem[3157] : 
                        (N233)? mem[3230] : 
                        (N235)? mem[3303] : 
                        (N237)? mem[3376] : 
                        (N239)? mem[3449] : 
                        (N241)? mem[3522] : 
                        (N243)? mem[3595] : 
                        (N245)? mem[3668] : 
                        (N247)? mem[3741] : 
                        (N249)? mem[3814] : 
                        (N251)? mem[3887] : 
                        (N253)? mem[3960] : 
                        (N255)? mem[4033] : 
                        (N257)? mem[4106] : 
                        (N259)? mem[4179] : 
                        (N261)? mem[4252] : 
                        (N263)? mem[4325] : 
                        (N265)? mem[4398] : 
                        (N267)? mem[4471] : 
                        (N269)? mem[4544] : 
                        (N271)? mem[4617] : 
                        (N146)? mem[4690] : 
                        (N148)? mem[4763] : 
                        (N150)? mem[4836] : 
                        (N152)? mem[4909] : 
                        (N154)? mem[4982] : 
                        (N156)? mem[5055] : 
                        (N158)? mem[5128] : 
                        (N160)? mem[5201] : 
                        (N162)? mem[5274] : 
                        (N164)? mem[5347] : 
                        (N166)? mem[5420] : 
                        (N168)? mem[5493] : 
                        (N170)? mem[5566] : 
                        (N172)? mem[5639] : 
                        (N174)? mem[5712] : 
                        (N176)? mem[5785] : 
                        (N178)? mem[5858] : 
                        (N180)? mem[5931] : 
                        (N182)? mem[6004] : 
                        (N184)? mem[6077] : 
                        (N186)? mem[6150] : 
                        (N188)? mem[6223] : 
                        (N190)? mem[6296] : 
                        (N192)? mem[6369] : 
                        (N194)? mem[6442] : 
                        (N196)? mem[6515] : 
                        (N198)? mem[6588] : 
                        (N200)? mem[6661] : 
                        (N202)? mem[6734] : 
                        (N204)? mem[6807] : 
                        (N206)? mem[6880] : 
                        (N208)? mem[6953] : 
                        (N210)? mem[7026] : 
                        (N212)? mem[7099] : 
                        (N214)? mem[7172] : 
                        (N216)? mem[7245] : 
                        (N218)? mem[7318] : 
                        (N220)? mem[7391] : 
                        (N222)? mem[7464] : 
                        (N224)? mem[7537] : 
                        (N226)? mem[7610] : 
                        (N228)? mem[7683] : 
                        (N230)? mem[7756] : 
                        (N232)? mem[7829] : 
                        (N234)? mem[7902] : 
                        (N236)? mem[7975] : 
                        (N238)? mem[8048] : 
                        (N240)? mem[8121] : 
                        (N242)? mem[8194] : 
                        (N244)? mem[8267] : 
                        (N246)? mem[8340] : 
                        (N248)? mem[8413] : 
                        (N250)? mem[8486] : 
                        (N252)? mem[8559] : 
                        (N254)? mem[8632] : 
                        (N256)? mem[8705] : 
                        (N258)? mem[8778] : 
                        (N260)? mem[8851] : 
                        (N262)? mem[8924] : 
                        (N264)? mem[8997] : 
                        (N266)? mem[9070] : 
                        (N268)? mem[9143] : 
                        (N270)? mem[9216] : 
                        (N272)? mem[9289] : 1'b0;
  assign r_data_o[17] = (N145)? mem[17] : 
                        (N147)? mem[90] : 
                        (N149)? mem[163] : 
                        (N151)? mem[236] : 
                        (N153)? mem[309] : 
                        (N155)? mem[382] : 
                        (N157)? mem[455] : 
                        (N159)? mem[528] : 
                        (N161)? mem[601] : 
                        (N163)? mem[674] : 
                        (N165)? mem[747] : 
                        (N167)? mem[820] : 
                        (N169)? mem[893] : 
                        (N171)? mem[966] : 
                        (N173)? mem[1039] : 
                        (N175)? mem[1112] : 
                        (N177)? mem[1185] : 
                        (N179)? mem[1258] : 
                        (N181)? mem[1331] : 
                        (N183)? mem[1404] : 
                        (N185)? mem[1477] : 
                        (N187)? mem[1550] : 
                        (N189)? mem[1623] : 
                        (N191)? mem[1696] : 
                        (N193)? mem[1769] : 
                        (N195)? mem[1842] : 
                        (N197)? mem[1915] : 
                        (N199)? mem[1988] : 
                        (N201)? mem[2061] : 
                        (N203)? mem[2134] : 
                        (N205)? mem[2207] : 
                        (N207)? mem[2280] : 
                        (N209)? mem[2353] : 
                        (N211)? mem[2426] : 
                        (N213)? mem[2499] : 
                        (N215)? mem[2572] : 
                        (N217)? mem[2645] : 
                        (N219)? mem[2718] : 
                        (N221)? mem[2791] : 
                        (N223)? mem[2864] : 
                        (N225)? mem[2937] : 
                        (N227)? mem[3010] : 
                        (N229)? mem[3083] : 
                        (N231)? mem[3156] : 
                        (N233)? mem[3229] : 
                        (N235)? mem[3302] : 
                        (N237)? mem[3375] : 
                        (N239)? mem[3448] : 
                        (N241)? mem[3521] : 
                        (N243)? mem[3594] : 
                        (N245)? mem[3667] : 
                        (N247)? mem[3740] : 
                        (N249)? mem[3813] : 
                        (N251)? mem[3886] : 
                        (N253)? mem[3959] : 
                        (N255)? mem[4032] : 
                        (N257)? mem[4105] : 
                        (N259)? mem[4178] : 
                        (N261)? mem[4251] : 
                        (N263)? mem[4324] : 
                        (N265)? mem[4397] : 
                        (N267)? mem[4470] : 
                        (N269)? mem[4543] : 
                        (N271)? mem[4616] : 
                        (N146)? mem[4689] : 
                        (N148)? mem[4762] : 
                        (N150)? mem[4835] : 
                        (N152)? mem[4908] : 
                        (N154)? mem[4981] : 
                        (N156)? mem[5054] : 
                        (N158)? mem[5127] : 
                        (N160)? mem[5200] : 
                        (N162)? mem[5273] : 
                        (N164)? mem[5346] : 
                        (N166)? mem[5419] : 
                        (N168)? mem[5492] : 
                        (N170)? mem[5565] : 
                        (N172)? mem[5638] : 
                        (N174)? mem[5711] : 
                        (N176)? mem[5784] : 
                        (N178)? mem[5857] : 
                        (N180)? mem[5930] : 
                        (N182)? mem[6003] : 
                        (N184)? mem[6076] : 
                        (N186)? mem[6149] : 
                        (N188)? mem[6222] : 
                        (N190)? mem[6295] : 
                        (N192)? mem[6368] : 
                        (N194)? mem[6441] : 
                        (N196)? mem[6514] : 
                        (N198)? mem[6587] : 
                        (N200)? mem[6660] : 
                        (N202)? mem[6733] : 
                        (N204)? mem[6806] : 
                        (N206)? mem[6879] : 
                        (N208)? mem[6952] : 
                        (N210)? mem[7025] : 
                        (N212)? mem[7098] : 
                        (N214)? mem[7171] : 
                        (N216)? mem[7244] : 
                        (N218)? mem[7317] : 
                        (N220)? mem[7390] : 
                        (N222)? mem[7463] : 
                        (N224)? mem[7536] : 
                        (N226)? mem[7609] : 
                        (N228)? mem[7682] : 
                        (N230)? mem[7755] : 
                        (N232)? mem[7828] : 
                        (N234)? mem[7901] : 
                        (N236)? mem[7974] : 
                        (N238)? mem[8047] : 
                        (N240)? mem[8120] : 
                        (N242)? mem[8193] : 
                        (N244)? mem[8266] : 
                        (N246)? mem[8339] : 
                        (N248)? mem[8412] : 
                        (N250)? mem[8485] : 
                        (N252)? mem[8558] : 
                        (N254)? mem[8631] : 
                        (N256)? mem[8704] : 
                        (N258)? mem[8777] : 
                        (N260)? mem[8850] : 
                        (N262)? mem[8923] : 
                        (N264)? mem[8996] : 
                        (N266)? mem[9069] : 
                        (N268)? mem[9142] : 
                        (N270)? mem[9215] : 
                        (N272)? mem[9288] : 1'b0;
  assign r_data_o[16] = (N145)? mem[16] : 
                        (N147)? mem[89] : 
                        (N149)? mem[162] : 
                        (N151)? mem[235] : 
                        (N153)? mem[308] : 
                        (N155)? mem[381] : 
                        (N157)? mem[454] : 
                        (N159)? mem[527] : 
                        (N161)? mem[600] : 
                        (N163)? mem[673] : 
                        (N165)? mem[746] : 
                        (N167)? mem[819] : 
                        (N169)? mem[892] : 
                        (N171)? mem[965] : 
                        (N173)? mem[1038] : 
                        (N175)? mem[1111] : 
                        (N177)? mem[1184] : 
                        (N179)? mem[1257] : 
                        (N181)? mem[1330] : 
                        (N183)? mem[1403] : 
                        (N185)? mem[1476] : 
                        (N187)? mem[1549] : 
                        (N189)? mem[1622] : 
                        (N191)? mem[1695] : 
                        (N193)? mem[1768] : 
                        (N195)? mem[1841] : 
                        (N197)? mem[1914] : 
                        (N199)? mem[1987] : 
                        (N201)? mem[2060] : 
                        (N203)? mem[2133] : 
                        (N205)? mem[2206] : 
                        (N207)? mem[2279] : 
                        (N209)? mem[2352] : 
                        (N211)? mem[2425] : 
                        (N213)? mem[2498] : 
                        (N215)? mem[2571] : 
                        (N217)? mem[2644] : 
                        (N219)? mem[2717] : 
                        (N221)? mem[2790] : 
                        (N223)? mem[2863] : 
                        (N225)? mem[2936] : 
                        (N227)? mem[3009] : 
                        (N229)? mem[3082] : 
                        (N231)? mem[3155] : 
                        (N233)? mem[3228] : 
                        (N235)? mem[3301] : 
                        (N237)? mem[3374] : 
                        (N239)? mem[3447] : 
                        (N241)? mem[3520] : 
                        (N243)? mem[3593] : 
                        (N245)? mem[3666] : 
                        (N247)? mem[3739] : 
                        (N249)? mem[3812] : 
                        (N251)? mem[3885] : 
                        (N253)? mem[3958] : 
                        (N255)? mem[4031] : 
                        (N257)? mem[4104] : 
                        (N259)? mem[4177] : 
                        (N261)? mem[4250] : 
                        (N263)? mem[4323] : 
                        (N265)? mem[4396] : 
                        (N267)? mem[4469] : 
                        (N269)? mem[4542] : 
                        (N271)? mem[4615] : 
                        (N146)? mem[4688] : 
                        (N148)? mem[4761] : 
                        (N150)? mem[4834] : 
                        (N152)? mem[4907] : 
                        (N154)? mem[4980] : 
                        (N156)? mem[5053] : 
                        (N158)? mem[5126] : 
                        (N160)? mem[5199] : 
                        (N162)? mem[5272] : 
                        (N164)? mem[5345] : 
                        (N166)? mem[5418] : 
                        (N168)? mem[5491] : 
                        (N170)? mem[5564] : 
                        (N172)? mem[5637] : 
                        (N174)? mem[5710] : 
                        (N176)? mem[5783] : 
                        (N178)? mem[5856] : 
                        (N180)? mem[5929] : 
                        (N182)? mem[6002] : 
                        (N184)? mem[6075] : 
                        (N186)? mem[6148] : 
                        (N188)? mem[6221] : 
                        (N190)? mem[6294] : 
                        (N192)? mem[6367] : 
                        (N194)? mem[6440] : 
                        (N196)? mem[6513] : 
                        (N198)? mem[6586] : 
                        (N200)? mem[6659] : 
                        (N202)? mem[6732] : 
                        (N204)? mem[6805] : 
                        (N206)? mem[6878] : 
                        (N208)? mem[6951] : 
                        (N210)? mem[7024] : 
                        (N212)? mem[7097] : 
                        (N214)? mem[7170] : 
                        (N216)? mem[7243] : 
                        (N218)? mem[7316] : 
                        (N220)? mem[7389] : 
                        (N222)? mem[7462] : 
                        (N224)? mem[7535] : 
                        (N226)? mem[7608] : 
                        (N228)? mem[7681] : 
                        (N230)? mem[7754] : 
                        (N232)? mem[7827] : 
                        (N234)? mem[7900] : 
                        (N236)? mem[7973] : 
                        (N238)? mem[8046] : 
                        (N240)? mem[8119] : 
                        (N242)? mem[8192] : 
                        (N244)? mem[8265] : 
                        (N246)? mem[8338] : 
                        (N248)? mem[8411] : 
                        (N250)? mem[8484] : 
                        (N252)? mem[8557] : 
                        (N254)? mem[8630] : 
                        (N256)? mem[8703] : 
                        (N258)? mem[8776] : 
                        (N260)? mem[8849] : 
                        (N262)? mem[8922] : 
                        (N264)? mem[8995] : 
                        (N266)? mem[9068] : 
                        (N268)? mem[9141] : 
                        (N270)? mem[9214] : 
                        (N272)? mem[9287] : 1'b0;
  assign r_data_o[15] = (N145)? mem[15] : 
                        (N147)? mem[88] : 
                        (N149)? mem[161] : 
                        (N151)? mem[234] : 
                        (N153)? mem[307] : 
                        (N155)? mem[380] : 
                        (N157)? mem[453] : 
                        (N159)? mem[526] : 
                        (N161)? mem[599] : 
                        (N163)? mem[672] : 
                        (N165)? mem[745] : 
                        (N167)? mem[818] : 
                        (N169)? mem[891] : 
                        (N171)? mem[964] : 
                        (N173)? mem[1037] : 
                        (N175)? mem[1110] : 
                        (N177)? mem[1183] : 
                        (N179)? mem[1256] : 
                        (N181)? mem[1329] : 
                        (N183)? mem[1402] : 
                        (N185)? mem[1475] : 
                        (N187)? mem[1548] : 
                        (N189)? mem[1621] : 
                        (N191)? mem[1694] : 
                        (N193)? mem[1767] : 
                        (N195)? mem[1840] : 
                        (N197)? mem[1913] : 
                        (N199)? mem[1986] : 
                        (N201)? mem[2059] : 
                        (N203)? mem[2132] : 
                        (N205)? mem[2205] : 
                        (N207)? mem[2278] : 
                        (N209)? mem[2351] : 
                        (N211)? mem[2424] : 
                        (N213)? mem[2497] : 
                        (N215)? mem[2570] : 
                        (N217)? mem[2643] : 
                        (N219)? mem[2716] : 
                        (N221)? mem[2789] : 
                        (N223)? mem[2862] : 
                        (N225)? mem[2935] : 
                        (N227)? mem[3008] : 
                        (N229)? mem[3081] : 
                        (N231)? mem[3154] : 
                        (N233)? mem[3227] : 
                        (N235)? mem[3300] : 
                        (N237)? mem[3373] : 
                        (N239)? mem[3446] : 
                        (N241)? mem[3519] : 
                        (N243)? mem[3592] : 
                        (N245)? mem[3665] : 
                        (N247)? mem[3738] : 
                        (N249)? mem[3811] : 
                        (N251)? mem[3884] : 
                        (N253)? mem[3957] : 
                        (N255)? mem[4030] : 
                        (N257)? mem[4103] : 
                        (N259)? mem[4176] : 
                        (N261)? mem[4249] : 
                        (N263)? mem[4322] : 
                        (N265)? mem[4395] : 
                        (N267)? mem[4468] : 
                        (N269)? mem[4541] : 
                        (N271)? mem[4614] : 
                        (N146)? mem[4687] : 
                        (N148)? mem[4760] : 
                        (N150)? mem[4833] : 
                        (N152)? mem[4906] : 
                        (N154)? mem[4979] : 
                        (N156)? mem[5052] : 
                        (N158)? mem[5125] : 
                        (N160)? mem[5198] : 
                        (N162)? mem[5271] : 
                        (N164)? mem[5344] : 
                        (N166)? mem[5417] : 
                        (N168)? mem[5490] : 
                        (N170)? mem[5563] : 
                        (N172)? mem[5636] : 
                        (N174)? mem[5709] : 
                        (N176)? mem[5782] : 
                        (N178)? mem[5855] : 
                        (N180)? mem[5928] : 
                        (N182)? mem[6001] : 
                        (N184)? mem[6074] : 
                        (N186)? mem[6147] : 
                        (N188)? mem[6220] : 
                        (N190)? mem[6293] : 
                        (N192)? mem[6366] : 
                        (N194)? mem[6439] : 
                        (N196)? mem[6512] : 
                        (N198)? mem[6585] : 
                        (N200)? mem[6658] : 
                        (N202)? mem[6731] : 
                        (N204)? mem[6804] : 
                        (N206)? mem[6877] : 
                        (N208)? mem[6950] : 
                        (N210)? mem[7023] : 
                        (N212)? mem[7096] : 
                        (N214)? mem[7169] : 
                        (N216)? mem[7242] : 
                        (N218)? mem[7315] : 
                        (N220)? mem[7388] : 
                        (N222)? mem[7461] : 
                        (N224)? mem[7534] : 
                        (N226)? mem[7607] : 
                        (N228)? mem[7680] : 
                        (N230)? mem[7753] : 
                        (N232)? mem[7826] : 
                        (N234)? mem[7899] : 
                        (N236)? mem[7972] : 
                        (N238)? mem[8045] : 
                        (N240)? mem[8118] : 
                        (N242)? mem[8191] : 
                        (N244)? mem[8264] : 
                        (N246)? mem[8337] : 
                        (N248)? mem[8410] : 
                        (N250)? mem[8483] : 
                        (N252)? mem[8556] : 
                        (N254)? mem[8629] : 
                        (N256)? mem[8702] : 
                        (N258)? mem[8775] : 
                        (N260)? mem[8848] : 
                        (N262)? mem[8921] : 
                        (N264)? mem[8994] : 
                        (N266)? mem[9067] : 
                        (N268)? mem[9140] : 
                        (N270)? mem[9213] : 
                        (N272)? mem[9286] : 1'b0;
  assign r_data_o[14] = (N145)? mem[14] : 
                        (N147)? mem[87] : 
                        (N149)? mem[160] : 
                        (N151)? mem[233] : 
                        (N153)? mem[306] : 
                        (N155)? mem[379] : 
                        (N157)? mem[452] : 
                        (N159)? mem[525] : 
                        (N161)? mem[598] : 
                        (N163)? mem[671] : 
                        (N165)? mem[744] : 
                        (N167)? mem[817] : 
                        (N169)? mem[890] : 
                        (N171)? mem[963] : 
                        (N173)? mem[1036] : 
                        (N175)? mem[1109] : 
                        (N177)? mem[1182] : 
                        (N179)? mem[1255] : 
                        (N181)? mem[1328] : 
                        (N183)? mem[1401] : 
                        (N185)? mem[1474] : 
                        (N187)? mem[1547] : 
                        (N189)? mem[1620] : 
                        (N191)? mem[1693] : 
                        (N193)? mem[1766] : 
                        (N195)? mem[1839] : 
                        (N197)? mem[1912] : 
                        (N199)? mem[1985] : 
                        (N201)? mem[2058] : 
                        (N203)? mem[2131] : 
                        (N205)? mem[2204] : 
                        (N207)? mem[2277] : 
                        (N209)? mem[2350] : 
                        (N211)? mem[2423] : 
                        (N213)? mem[2496] : 
                        (N215)? mem[2569] : 
                        (N217)? mem[2642] : 
                        (N219)? mem[2715] : 
                        (N221)? mem[2788] : 
                        (N223)? mem[2861] : 
                        (N225)? mem[2934] : 
                        (N227)? mem[3007] : 
                        (N229)? mem[3080] : 
                        (N231)? mem[3153] : 
                        (N233)? mem[3226] : 
                        (N235)? mem[3299] : 
                        (N237)? mem[3372] : 
                        (N239)? mem[3445] : 
                        (N241)? mem[3518] : 
                        (N243)? mem[3591] : 
                        (N245)? mem[3664] : 
                        (N247)? mem[3737] : 
                        (N249)? mem[3810] : 
                        (N251)? mem[3883] : 
                        (N253)? mem[3956] : 
                        (N255)? mem[4029] : 
                        (N257)? mem[4102] : 
                        (N259)? mem[4175] : 
                        (N261)? mem[4248] : 
                        (N263)? mem[4321] : 
                        (N265)? mem[4394] : 
                        (N267)? mem[4467] : 
                        (N269)? mem[4540] : 
                        (N271)? mem[4613] : 
                        (N146)? mem[4686] : 
                        (N148)? mem[4759] : 
                        (N150)? mem[4832] : 
                        (N152)? mem[4905] : 
                        (N154)? mem[4978] : 
                        (N156)? mem[5051] : 
                        (N158)? mem[5124] : 
                        (N160)? mem[5197] : 
                        (N162)? mem[5270] : 
                        (N164)? mem[5343] : 
                        (N166)? mem[5416] : 
                        (N168)? mem[5489] : 
                        (N170)? mem[5562] : 
                        (N172)? mem[5635] : 
                        (N174)? mem[5708] : 
                        (N176)? mem[5781] : 
                        (N178)? mem[5854] : 
                        (N180)? mem[5927] : 
                        (N182)? mem[6000] : 
                        (N184)? mem[6073] : 
                        (N186)? mem[6146] : 
                        (N188)? mem[6219] : 
                        (N190)? mem[6292] : 
                        (N192)? mem[6365] : 
                        (N194)? mem[6438] : 
                        (N196)? mem[6511] : 
                        (N198)? mem[6584] : 
                        (N200)? mem[6657] : 
                        (N202)? mem[6730] : 
                        (N204)? mem[6803] : 
                        (N206)? mem[6876] : 
                        (N208)? mem[6949] : 
                        (N210)? mem[7022] : 
                        (N212)? mem[7095] : 
                        (N214)? mem[7168] : 
                        (N216)? mem[7241] : 
                        (N218)? mem[7314] : 
                        (N220)? mem[7387] : 
                        (N222)? mem[7460] : 
                        (N224)? mem[7533] : 
                        (N226)? mem[7606] : 
                        (N228)? mem[7679] : 
                        (N230)? mem[7752] : 
                        (N232)? mem[7825] : 
                        (N234)? mem[7898] : 
                        (N236)? mem[7971] : 
                        (N238)? mem[8044] : 
                        (N240)? mem[8117] : 
                        (N242)? mem[8190] : 
                        (N244)? mem[8263] : 
                        (N246)? mem[8336] : 
                        (N248)? mem[8409] : 
                        (N250)? mem[8482] : 
                        (N252)? mem[8555] : 
                        (N254)? mem[8628] : 
                        (N256)? mem[8701] : 
                        (N258)? mem[8774] : 
                        (N260)? mem[8847] : 
                        (N262)? mem[8920] : 
                        (N264)? mem[8993] : 
                        (N266)? mem[9066] : 
                        (N268)? mem[9139] : 
                        (N270)? mem[9212] : 
                        (N272)? mem[9285] : 1'b0;
  assign r_data_o[13] = (N145)? mem[13] : 
                        (N147)? mem[86] : 
                        (N149)? mem[159] : 
                        (N151)? mem[232] : 
                        (N153)? mem[305] : 
                        (N155)? mem[378] : 
                        (N157)? mem[451] : 
                        (N159)? mem[524] : 
                        (N161)? mem[597] : 
                        (N163)? mem[670] : 
                        (N165)? mem[743] : 
                        (N167)? mem[816] : 
                        (N169)? mem[889] : 
                        (N171)? mem[962] : 
                        (N173)? mem[1035] : 
                        (N175)? mem[1108] : 
                        (N177)? mem[1181] : 
                        (N179)? mem[1254] : 
                        (N181)? mem[1327] : 
                        (N183)? mem[1400] : 
                        (N185)? mem[1473] : 
                        (N187)? mem[1546] : 
                        (N189)? mem[1619] : 
                        (N191)? mem[1692] : 
                        (N193)? mem[1765] : 
                        (N195)? mem[1838] : 
                        (N197)? mem[1911] : 
                        (N199)? mem[1984] : 
                        (N201)? mem[2057] : 
                        (N203)? mem[2130] : 
                        (N205)? mem[2203] : 
                        (N207)? mem[2276] : 
                        (N209)? mem[2349] : 
                        (N211)? mem[2422] : 
                        (N213)? mem[2495] : 
                        (N215)? mem[2568] : 
                        (N217)? mem[2641] : 
                        (N219)? mem[2714] : 
                        (N221)? mem[2787] : 
                        (N223)? mem[2860] : 
                        (N225)? mem[2933] : 
                        (N227)? mem[3006] : 
                        (N229)? mem[3079] : 
                        (N231)? mem[3152] : 
                        (N233)? mem[3225] : 
                        (N235)? mem[3298] : 
                        (N237)? mem[3371] : 
                        (N239)? mem[3444] : 
                        (N241)? mem[3517] : 
                        (N243)? mem[3590] : 
                        (N245)? mem[3663] : 
                        (N247)? mem[3736] : 
                        (N249)? mem[3809] : 
                        (N251)? mem[3882] : 
                        (N253)? mem[3955] : 
                        (N255)? mem[4028] : 
                        (N257)? mem[4101] : 
                        (N259)? mem[4174] : 
                        (N261)? mem[4247] : 
                        (N263)? mem[4320] : 
                        (N265)? mem[4393] : 
                        (N267)? mem[4466] : 
                        (N269)? mem[4539] : 
                        (N271)? mem[4612] : 
                        (N146)? mem[4685] : 
                        (N148)? mem[4758] : 
                        (N150)? mem[4831] : 
                        (N152)? mem[4904] : 
                        (N154)? mem[4977] : 
                        (N156)? mem[5050] : 
                        (N158)? mem[5123] : 
                        (N160)? mem[5196] : 
                        (N162)? mem[5269] : 
                        (N164)? mem[5342] : 
                        (N166)? mem[5415] : 
                        (N168)? mem[5488] : 
                        (N170)? mem[5561] : 
                        (N172)? mem[5634] : 
                        (N174)? mem[5707] : 
                        (N176)? mem[5780] : 
                        (N178)? mem[5853] : 
                        (N180)? mem[5926] : 
                        (N182)? mem[5999] : 
                        (N184)? mem[6072] : 
                        (N186)? mem[6145] : 
                        (N188)? mem[6218] : 
                        (N190)? mem[6291] : 
                        (N192)? mem[6364] : 
                        (N194)? mem[6437] : 
                        (N196)? mem[6510] : 
                        (N198)? mem[6583] : 
                        (N200)? mem[6656] : 
                        (N202)? mem[6729] : 
                        (N204)? mem[6802] : 
                        (N206)? mem[6875] : 
                        (N208)? mem[6948] : 
                        (N210)? mem[7021] : 
                        (N212)? mem[7094] : 
                        (N214)? mem[7167] : 
                        (N216)? mem[7240] : 
                        (N218)? mem[7313] : 
                        (N220)? mem[7386] : 
                        (N222)? mem[7459] : 
                        (N224)? mem[7532] : 
                        (N226)? mem[7605] : 
                        (N228)? mem[7678] : 
                        (N230)? mem[7751] : 
                        (N232)? mem[7824] : 
                        (N234)? mem[7897] : 
                        (N236)? mem[7970] : 
                        (N238)? mem[8043] : 
                        (N240)? mem[8116] : 
                        (N242)? mem[8189] : 
                        (N244)? mem[8262] : 
                        (N246)? mem[8335] : 
                        (N248)? mem[8408] : 
                        (N250)? mem[8481] : 
                        (N252)? mem[8554] : 
                        (N254)? mem[8627] : 
                        (N256)? mem[8700] : 
                        (N258)? mem[8773] : 
                        (N260)? mem[8846] : 
                        (N262)? mem[8919] : 
                        (N264)? mem[8992] : 
                        (N266)? mem[9065] : 
                        (N268)? mem[9138] : 
                        (N270)? mem[9211] : 
                        (N272)? mem[9284] : 1'b0;
  assign r_data_o[12] = (N145)? mem[12] : 
                        (N147)? mem[85] : 
                        (N149)? mem[158] : 
                        (N151)? mem[231] : 
                        (N153)? mem[304] : 
                        (N155)? mem[377] : 
                        (N157)? mem[450] : 
                        (N159)? mem[523] : 
                        (N161)? mem[596] : 
                        (N163)? mem[669] : 
                        (N165)? mem[742] : 
                        (N167)? mem[815] : 
                        (N169)? mem[888] : 
                        (N171)? mem[961] : 
                        (N173)? mem[1034] : 
                        (N175)? mem[1107] : 
                        (N177)? mem[1180] : 
                        (N179)? mem[1253] : 
                        (N181)? mem[1326] : 
                        (N183)? mem[1399] : 
                        (N185)? mem[1472] : 
                        (N187)? mem[1545] : 
                        (N189)? mem[1618] : 
                        (N191)? mem[1691] : 
                        (N193)? mem[1764] : 
                        (N195)? mem[1837] : 
                        (N197)? mem[1910] : 
                        (N199)? mem[1983] : 
                        (N201)? mem[2056] : 
                        (N203)? mem[2129] : 
                        (N205)? mem[2202] : 
                        (N207)? mem[2275] : 
                        (N209)? mem[2348] : 
                        (N211)? mem[2421] : 
                        (N213)? mem[2494] : 
                        (N215)? mem[2567] : 
                        (N217)? mem[2640] : 
                        (N219)? mem[2713] : 
                        (N221)? mem[2786] : 
                        (N223)? mem[2859] : 
                        (N225)? mem[2932] : 
                        (N227)? mem[3005] : 
                        (N229)? mem[3078] : 
                        (N231)? mem[3151] : 
                        (N233)? mem[3224] : 
                        (N235)? mem[3297] : 
                        (N237)? mem[3370] : 
                        (N239)? mem[3443] : 
                        (N241)? mem[3516] : 
                        (N243)? mem[3589] : 
                        (N245)? mem[3662] : 
                        (N247)? mem[3735] : 
                        (N249)? mem[3808] : 
                        (N251)? mem[3881] : 
                        (N253)? mem[3954] : 
                        (N255)? mem[4027] : 
                        (N257)? mem[4100] : 
                        (N259)? mem[4173] : 
                        (N261)? mem[4246] : 
                        (N263)? mem[4319] : 
                        (N265)? mem[4392] : 
                        (N267)? mem[4465] : 
                        (N269)? mem[4538] : 
                        (N271)? mem[4611] : 
                        (N146)? mem[4684] : 
                        (N148)? mem[4757] : 
                        (N150)? mem[4830] : 
                        (N152)? mem[4903] : 
                        (N154)? mem[4976] : 
                        (N156)? mem[5049] : 
                        (N158)? mem[5122] : 
                        (N160)? mem[5195] : 
                        (N162)? mem[5268] : 
                        (N164)? mem[5341] : 
                        (N166)? mem[5414] : 
                        (N168)? mem[5487] : 
                        (N170)? mem[5560] : 
                        (N172)? mem[5633] : 
                        (N174)? mem[5706] : 
                        (N176)? mem[5779] : 
                        (N178)? mem[5852] : 
                        (N180)? mem[5925] : 
                        (N182)? mem[5998] : 
                        (N184)? mem[6071] : 
                        (N186)? mem[6144] : 
                        (N188)? mem[6217] : 
                        (N190)? mem[6290] : 
                        (N192)? mem[6363] : 
                        (N194)? mem[6436] : 
                        (N196)? mem[6509] : 
                        (N198)? mem[6582] : 
                        (N200)? mem[6655] : 
                        (N202)? mem[6728] : 
                        (N204)? mem[6801] : 
                        (N206)? mem[6874] : 
                        (N208)? mem[6947] : 
                        (N210)? mem[7020] : 
                        (N212)? mem[7093] : 
                        (N214)? mem[7166] : 
                        (N216)? mem[7239] : 
                        (N218)? mem[7312] : 
                        (N220)? mem[7385] : 
                        (N222)? mem[7458] : 
                        (N224)? mem[7531] : 
                        (N226)? mem[7604] : 
                        (N228)? mem[7677] : 
                        (N230)? mem[7750] : 
                        (N232)? mem[7823] : 
                        (N234)? mem[7896] : 
                        (N236)? mem[7969] : 
                        (N238)? mem[8042] : 
                        (N240)? mem[8115] : 
                        (N242)? mem[8188] : 
                        (N244)? mem[8261] : 
                        (N246)? mem[8334] : 
                        (N248)? mem[8407] : 
                        (N250)? mem[8480] : 
                        (N252)? mem[8553] : 
                        (N254)? mem[8626] : 
                        (N256)? mem[8699] : 
                        (N258)? mem[8772] : 
                        (N260)? mem[8845] : 
                        (N262)? mem[8918] : 
                        (N264)? mem[8991] : 
                        (N266)? mem[9064] : 
                        (N268)? mem[9137] : 
                        (N270)? mem[9210] : 
                        (N272)? mem[9283] : 1'b0;
  assign r_data_o[11] = (N145)? mem[11] : 
                        (N147)? mem[84] : 
                        (N149)? mem[157] : 
                        (N151)? mem[230] : 
                        (N153)? mem[303] : 
                        (N155)? mem[376] : 
                        (N157)? mem[449] : 
                        (N159)? mem[522] : 
                        (N161)? mem[595] : 
                        (N163)? mem[668] : 
                        (N165)? mem[741] : 
                        (N167)? mem[814] : 
                        (N169)? mem[887] : 
                        (N171)? mem[960] : 
                        (N173)? mem[1033] : 
                        (N175)? mem[1106] : 
                        (N177)? mem[1179] : 
                        (N179)? mem[1252] : 
                        (N181)? mem[1325] : 
                        (N183)? mem[1398] : 
                        (N185)? mem[1471] : 
                        (N187)? mem[1544] : 
                        (N189)? mem[1617] : 
                        (N191)? mem[1690] : 
                        (N193)? mem[1763] : 
                        (N195)? mem[1836] : 
                        (N197)? mem[1909] : 
                        (N199)? mem[1982] : 
                        (N201)? mem[2055] : 
                        (N203)? mem[2128] : 
                        (N205)? mem[2201] : 
                        (N207)? mem[2274] : 
                        (N209)? mem[2347] : 
                        (N211)? mem[2420] : 
                        (N213)? mem[2493] : 
                        (N215)? mem[2566] : 
                        (N217)? mem[2639] : 
                        (N219)? mem[2712] : 
                        (N221)? mem[2785] : 
                        (N223)? mem[2858] : 
                        (N225)? mem[2931] : 
                        (N227)? mem[3004] : 
                        (N229)? mem[3077] : 
                        (N231)? mem[3150] : 
                        (N233)? mem[3223] : 
                        (N235)? mem[3296] : 
                        (N237)? mem[3369] : 
                        (N239)? mem[3442] : 
                        (N241)? mem[3515] : 
                        (N243)? mem[3588] : 
                        (N245)? mem[3661] : 
                        (N247)? mem[3734] : 
                        (N249)? mem[3807] : 
                        (N251)? mem[3880] : 
                        (N253)? mem[3953] : 
                        (N255)? mem[4026] : 
                        (N257)? mem[4099] : 
                        (N259)? mem[4172] : 
                        (N261)? mem[4245] : 
                        (N263)? mem[4318] : 
                        (N265)? mem[4391] : 
                        (N267)? mem[4464] : 
                        (N269)? mem[4537] : 
                        (N271)? mem[4610] : 
                        (N146)? mem[4683] : 
                        (N148)? mem[4756] : 
                        (N150)? mem[4829] : 
                        (N152)? mem[4902] : 
                        (N154)? mem[4975] : 
                        (N156)? mem[5048] : 
                        (N158)? mem[5121] : 
                        (N160)? mem[5194] : 
                        (N162)? mem[5267] : 
                        (N164)? mem[5340] : 
                        (N166)? mem[5413] : 
                        (N168)? mem[5486] : 
                        (N170)? mem[5559] : 
                        (N172)? mem[5632] : 
                        (N174)? mem[5705] : 
                        (N176)? mem[5778] : 
                        (N178)? mem[5851] : 
                        (N180)? mem[5924] : 
                        (N182)? mem[5997] : 
                        (N184)? mem[6070] : 
                        (N186)? mem[6143] : 
                        (N188)? mem[6216] : 
                        (N190)? mem[6289] : 
                        (N192)? mem[6362] : 
                        (N194)? mem[6435] : 
                        (N196)? mem[6508] : 
                        (N198)? mem[6581] : 
                        (N200)? mem[6654] : 
                        (N202)? mem[6727] : 
                        (N204)? mem[6800] : 
                        (N206)? mem[6873] : 
                        (N208)? mem[6946] : 
                        (N210)? mem[7019] : 
                        (N212)? mem[7092] : 
                        (N214)? mem[7165] : 
                        (N216)? mem[7238] : 
                        (N218)? mem[7311] : 
                        (N220)? mem[7384] : 
                        (N222)? mem[7457] : 
                        (N224)? mem[7530] : 
                        (N226)? mem[7603] : 
                        (N228)? mem[7676] : 
                        (N230)? mem[7749] : 
                        (N232)? mem[7822] : 
                        (N234)? mem[7895] : 
                        (N236)? mem[7968] : 
                        (N238)? mem[8041] : 
                        (N240)? mem[8114] : 
                        (N242)? mem[8187] : 
                        (N244)? mem[8260] : 
                        (N246)? mem[8333] : 
                        (N248)? mem[8406] : 
                        (N250)? mem[8479] : 
                        (N252)? mem[8552] : 
                        (N254)? mem[8625] : 
                        (N256)? mem[8698] : 
                        (N258)? mem[8771] : 
                        (N260)? mem[8844] : 
                        (N262)? mem[8917] : 
                        (N264)? mem[8990] : 
                        (N266)? mem[9063] : 
                        (N268)? mem[9136] : 
                        (N270)? mem[9209] : 
                        (N272)? mem[9282] : 1'b0;
  assign r_data_o[10] = (N145)? mem[10] : 
                        (N147)? mem[83] : 
                        (N149)? mem[156] : 
                        (N151)? mem[229] : 
                        (N153)? mem[302] : 
                        (N155)? mem[375] : 
                        (N157)? mem[448] : 
                        (N159)? mem[521] : 
                        (N161)? mem[594] : 
                        (N163)? mem[667] : 
                        (N165)? mem[740] : 
                        (N167)? mem[813] : 
                        (N169)? mem[886] : 
                        (N171)? mem[959] : 
                        (N173)? mem[1032] : 
                        (N175)? mem[1105] : 
                        (N177)? mem[1178] : 
                        (N179)? mem[1251] : 
                        (N181)? mem[1324] : 
                        (N183)? mem[1397] : 
                        (N185)? mem[1470] : 
                        (N187)? mem[1543] : 
                        (N189)? mem[1616] : 
                        (N191)? mem[1689] : 
                        (N193)? mem[1762] : 
                        (N195)? mem[1835] : 
                        (N197)? mem[1908] : 
                        (N199)? mem[1981] : 
                        (N201)? mem[2054] : 
                        (N203)? mem[2127] : 
                        (N205)? mem[2200] : 
                        (N207)? mem[2273] : 
                        (N209)? mem[2346] : 
                        (N211)? mem[2419] : 
                        (N213)? mem[2492] : 
                        (N215)? mem[2565] : 
                        (N217)? mem[2638] : 
                        (N219)? mem[2711] : 
                        (N221)? mem[2784] : 
                        (N223)? mem[2857] : 
                        (N225)? mem[2930] : 
                        (N227)? mem[3003] : 
                        (N229)? mem[3076] : 
                        (N231)? mem[3149] : 
                        (N233)? mem[3222] : 
                        (N235)? mem[3295] : 
                        (N237)? mem[3368] : 
                        (N239)? mem[3441] : 
                        (N241)? mem[3514] : 
                        (N243)? mem[3587] : 
                        (N245)? mem[3660] : 
                        (N247)? mem[3733] : 
                        (N249)? mem[3806] : 
                        (N251)? mem[3879] : 
                        (N253)? mem[3952] : 
                        (N255)? mem[4025] : 
                        (N257)? mem[4098] : 
                        (N259)? mem[4171] : 
                        (N261)? mem[4244] : 
                        (N263)? mem[4317] : 
                        (N265)? mem[4390] : 
                        (N267)? mem[4463] : 
                        (N269)? mem[4536] : 
                        (N271)? mem[4609] : 
                        (N146)? mem[4682] : 
                        (N148)? mem[4755] : 
                        (N150)? mem[4828] : 
                        (N152)? mem[4901] : 
                        (N154)? mem[4974] : 
                        (N156)? mem[5047] : 
                        (N158)? mem[5120] : 
                        (N160)? mem[5193] : 
                        (N162)? mem[5266] : 
                        (N164)? mem[5339] : 
                        (N166)? mem[5412] : 
                        (N168)? mem[5485] : 
                        (N170)? mem[5558] : 
                        (N172)? mem[5631] : 
                        (N174)? mem[5704] : 
                        (N176)? mem[5777] : 
                        (N178)? mem[5850] : 
                        (N180)? mem[5923] : 
                        (N182)? mem[5996] : 
                        (N184)? mem[6069] : 
                        (N186)? mem[6142] : 
                        (N188)? mem[6215] : 
                        (N190)? mem[6288] : 
                        (N192)? mem[6361] : 
                        (N194)? mem[6434] : 
                        (N196)? mem[6507] : 
                        (N198)? mem[6580] : 
                        (N200)? mem[6653] : 
                        (N202)? mem[6726] : 
                        (N204)? mem[6799] : 
                        (N206)? mem[6872] : 
                        (N208)? mem[6945] : 
                        (N210)? mem[7018] : 
                        (N212)? mem[7091] : 
                        (N214)? mem[7164] : 
                        (N216)? mem[7237] : 
                        (N218)? mem[7310] : 
                        (N220)? mem[7383] : 
                        (N222)? mem[7456] : 
                        (N224)? mem[7529] : 
                        (N226)? mem[7602] : 
                        (N228)? mem[7675] : 
                        (N230)? mem[7748] : 
                        (N232)? mem[7821] : 
                        (N234)? mem[7894] : 
                        (N236)? mem[7967] : 
                        (N238)? mem[8040] : 
                        (N240)? mem[8113] : 
                        (N242)? mem[8186] : 
                        (N244)? mem[8259] : 
                        (N246)? mem[8332] : 
                        (N248)? mem[8405] : 
                        (N250)? mem[8478] : 
                        (N252)? mem[8551] : 
                        (N254)? mem[8624] : 
                        (N256)? mem[8697] : 
                        (N258)? mem[8770] : 
                        (N260)? mem[8843] : 
                        (N262)? mem[8916] : 
                        (N264)? mem[8989] : 
                        (N266)? mem[9062] : 
                        (N268)? mem[9135] : 
                        (N270)? mem[9208] : 
                        (N272)? mem[9281] : 1'b0;
  assign r_data_o[9] = (N145)? mem[9] : 
                       (N147)? mem[82] : 
                       (N149)? mem[155] : 
                       (N151)? mem[228] : 
                       (N153)? mem[301] : 
                       (N155)? mem[374] : 
                       (N157)? mem[447] : 
                       (N159)? mem[520] : 
                       (N161)? mem[593] : 
                       (N163)? mem[666] : 
                       (N165)? mem[739] : 
                       (N167)? mem[812] : 
                       (N169)? mem[885] : 
                       (N171)? mem[958] : 
                       (N173)? mem[1031] : 
                       (N175)? mem[1104] : 
                       (N177)? mem[1177] : 
                       (N179)? mem[1250] : 
                       (N181)? mem[1323] : 
                       (N183)? mem[1396] : 
                       (N185)? mem[1469] : 
                       (N187)? mem[1542] : 
                       (N189)? mem[1615] : 
                       (N191)? mem[1688] : 
                       (N193)? mem[1761] : 
                       (N195)? mem[1834] : 
                       (N197)? mem[1907] : 
                       (N199)? mem[1980] : 
                       (N201)? mem[2053] : 
                       (N203)? mem[2126] : 
                       (N205)? mem[2199] : 
                       (N207)? mem[2272] : 
                       (N209)? mem[2345] : 
                       (N211)? mem[2418] : 
                       (N213)? mem[2491] : 
                       (N215)? mem[2564] : 
                       (N217)? mem[2637] : 
                       (N219)? mem[2710] : 
                       (N221)? mem[2783] : 
                       (N223)? mem[2856] : 
                       (N225)? mem[2929] : 
                       (N227)? mem[3002] : 
                       (N229)? mem[3075] : 
                       (N231)? mem[3148] : 
                       (N233)? mem[3221] : 
                       (N235)? mem[3294] : 
                       (N237)? mem[3367] : 
                       (N239)? mem[3440] : 
                       (N241)? mem[3513] : 
                       (N243)? mem[3586] : 
                       (N245)? mem[3659] : 
                       (N247)? mem[3732] : 
                       (N249)? mem[3805] : 
                       (N251)? mem[3878] : 
                       (N253)? mem[3951] : 
                       (N255)? mem[4024] : 
                       (N257)? mem[4097] : 
                       (N259)? mem[4170] : 
                       (N261)? mem[4243] : 
                       (N263)? mem[4316] : 
                       (N265)? mem[4389] : 
                       (N267)? mem[4462] : 
                       (N269)? mem[4535] : 
                       (N271)? mem[4608] : 
                       (N146)? mem[4681] : 
                       (N148)? mem[4754] : 
                       (N150)? mem[4827] : 
                       (N152)? mem[4900] : 
                       (N154)? mem[4973] : 
                       (N156)? mem[5046] : 
                       (N158)? mem[5119] : 
                       (N160)? mem[5192] : 
                       (N162)? mem[5265] : 
                       (N164)? mem[5338] : 
                       (N166)? mem[5411] : 
                       (N168)? mem[5484] : 
                       (N170)? mem[5557] : 
                       (N172)? mem[5630] : 
                       (N174)? mem[5703] : 
                       (N176)? mem[5776] : 
                       (N178)? mem[5849] : 
                       (N180)? mem[5922] : 
                       (N182)? mem[5995] : 
                       (N184)? mem[6068] : 
                       (N186)? mem[6141] : 
                       (N188)? mem[6214] : 
                       (N190)? mem[6287] : 
                       (N192)? mem[6360] : 
                       (N194)? mem[6433] : 
                       (N196)? mem[6506] : 
                       (N198)? mem[6579] : 
                       (N200)? mem[6652] : 
                       (N202)? mem[6725] : 
                       (N204)? mem[6798] : 
                       (N206)? mem[6871] : 
                       (N208)? mem[6944] : 
                       (N210)? mem[7017] : 
                       (N212)? mem[7090] : 
                       (N214)? mem[7163] : 
                       (N216)? mem[7236] : 
                       (N218)? mem[7309] : 
                       (N220)? mem[7382] : 
                       (N222)? mem[7455] : 
                       (N224)? mem[7528] : 
                       (N226)? mem[7601] : 
                       (N228)? mem[7674] : 
                       (N230)? mem[7747] : 
                       (N232)? mem[7820] : 
                       (N234)? mem[7893] : 
                       (N236)? mem[7966] : 
                       (N238)? mem[8039] : 
                       (N240)? mem[8112] : 
                       (N242)? mem[8185] : 
                       (N244)? mem[8258] : 
                       (N246)? mem[8331] : 
                       (N248)? mem[8404] : 
                       (N250)? mem[8477] : 
                       (N252)? mem[8550] : 
                       (N254)? mem[8623] : 
                       (N256)? mem[8696] : 
                       (N258)? mem[8769] : 
                       (N260)? mem[8842] : 
                       (N262)? mem[8915] : 
                       (N264)? mem[8988] : 
                       (N266)? mem[9061] : 
                       (N268)? mem[9134] : 
                       (N270)? mem[9207] : 
                       (N272)? mem[9280] : 1'b0;
  assign r_data_o[8] = (N145)? mem[8] : 
                       (N147)? mem[81] : 
                       (N149)? mem[154] : 
                       (N151)? mem[227] : 
                       (N153)? mem[300] : 
                       (N155)? mem[373] : 
                       (N157)? mem[446] : 
                       (N159)? mem[519] : 
                       (N161)? mem[592] : 
                       (N163)? mem[665] : 
                       (N165)? mem[738] : 
                       (N167)? mem[811] : 
                       (N169)? mem[884] : 
                       (N171)? mem[957] : 
                       (N173)? mem[1030] : 
                       (N175)? mem[1103] : 
                       (N177)? mem[1176] : 
                       (N179)? mem[1249] : 
                       (N181)? mem[1322] : 
                       (N183)? mem[1395] : 
                       (N185)? mem[1468] : 
                       (N187)? mem[1541] : 
                       (N189)? mem[1614] : 
                       (N191)? mem[1687] : 
                       (N193)? mem[1760] : 
                       (N195)? mem[1833] : 
                       (N197)? mem[1906] : 
                       (N199)? mem[1979] : 
                       (N201)? mem[2052] : 
                       (N203)? mem[2125] : 
                       (N205)? mem[2198] : 
                       (N207)? mem[2271] : 
                       (N209)? mem[2344] : 
                       (N211)? mem[2417] : 
                       (N213)? mem[2490] : 
                       (N215)? mem[2563] : 
                       (N217)? mem[2636] : 
                       (N219)? mem[2709] : 
                       (N221)? mem[2782] : 
                       (N223)? mem[2855] : 
                       (N225)? mem[2928] : 
                       (N227)? mem[3001] : 
                       (N229)? mem[3074] : 
                       (N231)? mem[3147] : 
                       (N233)? mem[3220] : 
                       (N235)? mem[3293] : 
                       (N237)? mem[3366] : 
                       (N239)? mem[3439] : 
                       (N241)? mem[3512] : 
                       (N243)? mem[3585] : 
                       (N245)? mem[3658] : 
                       (N247)? mem[3731] : 
                       (N249)? mem[3804] : 
                       (N251)? mem[3877] : 
                       (N253)? mem[3950] : 
                       (N255)? mem[4023] : 
                       (N257)? mem[4096] : 
                       (N259)? mem[4169] : 
                       (N261)? mem[4242] : 
                       (N263)? mem[4315] : 
                       (N265)? mem[4388] : 
                       (N267)? mem[4461] : 
                       (N269)? mem[4534] : 
                       (N271)? mem[4607] : 
                       (N146)? mem[4680] : 
                       (N148)? mem[4753] : 
                       (N150)? mem[4826] : 
                       (N152)? mem[4899] : 
                       (N154)? mem[4972] : 
                       (N156)? mem[5045] : 
                       (N158)? mem[5118] : 
                       (N160)? mem[5191] : 
                       (N162)? mem[5264] : 
                       (N164)? mem[5337] : 
                       (N166)? mem[5410] : 
                       (N168)? mem[5483] : 
                       (N170)? mem[5556] : 
                       (N172)? mem[5629] : 
                       (N174)? mem[5702] : 
                       (N176)? mem[5775] : 
                       (N178)? mem[5848] : 
                       (N180)? mem[5921] : 
                       (N182)? mem[5994] : 
                       (N184)? mem[6067] : 
                       (N186)? mem[6140] : 
                       (N188)? mem[6213] : 
                       (N190)? mem[6286] : 
                       (N192)? mem[6359] : 
                       (N194)? mem[6432] : 
                       (N196)? mem[6505] : 
                       (N198)? mem[6578] : 
                       (N200)? mem[6651] : 
                       (N202)? mem[6724] : 
                       (N204)? mem[6797] : 
                       (N206)? mem[6870] : 
                       (N208)? mem[6943] : 
                       (N210)? mem[7016] : 
                       (N212)? mem[7089] : 
                       (N214)? mem[7162] : 
                       (N216)? mem[7235] : 
                       (N218)? mem[7308] : 
                       (N220)? mem[7381] : 
                       (N222)? mem[7454] : 
                       (N224)? mem[7527] : 
                       (N226)? mem[7600] : 
                       (N228)? mem[7673] : 
                       (N230)? mem[7746] : 
                       (N232)? mem[7819] : 
                       (N234)? mem[7892] : 
                       (N236)? mem[7965] : 
                       (N238)? mem[8038] : 
                       (N240)? mem[8111] : 
                       (N242)? mem[8184] : 
                       (N244)? mem[8257] : 
                       (N246)? mem[8330] : 
                       (N248)? mem[8403] : 
                       (N250)? mem[8476] : 
                       (N252)? mem[8549] : 
                       (N254)? mem[8622] : 
                       (N256)? mem[8695] : 
                       (N258)? mem[8768] : 
                       (N260)? mem[8841] : 
                       (N262)? mem[8914] : 
                       (N264)? mem[8987] : 
                       (N266)? mem[9060] : 
                       (N268)? mem[9133] : 
                       (N270)? mem[9206] : 
                       (N272)? mem[9279] : 1'b0;
  assign r_data_o[7] = (N145)? mem[7] : 
                       (N147)? mem[80] : 
                       (N149)? mem[153] : 
                       (N151)? mem[226] : 
                       (N153)? mem[299] : 
                       (N155)? mem[372] : 
                       (N157)? mem[445] : 
                       (N159)? mem[518] : 
                       (N161)? mem[591] : 
                       (N163)? mem[664] : 
                       (N165)? mem[737] : 
                       (N167)? mem[810] : 
                       (N169)? mem[883] : 
                       (N171)? mem[956] : 
                       (N173)? mem[1029] : 
                       (N175)? mem[1102] : 
                       (N177)? mem[1175] : 
                       (N179)? mem[1248] : 
                       (N181)? mem[1321] : 
                       (N183)? mem[1394] : 
                       (N185)? mem[1467] : 
                       (N187)? mem[1540] : 
                       (N189)? mem[1613] : 
                       (N191)? mem[1686] : 
                       (N193)? mem[1759] : 
                       (N195)? mem[1832] : 
                       (N197)? mem[1905] : 
                       (N199)? mem[1978] : 
                       (N201)? mem[2051] : 
                       (N203)? mem[2124] : 
                       (N205)? mem[2197] : 
                       (N207)? mem[2270] : 
                       (N209)? mem[2343] : 
                       (N211)? mem[2416] : 
                       (N213)? mem[2489] : 
                       (N215)? mem[2562] : 
                       (N217)? mem[2635] : 
                       (N219)? mem[2708] : 
                       (N221)? mem[2781] : 
                       (N223)? mem[2854] : 
                       (N225)? mem[2927] : 
                       (N227)? mem[3000] : 
                       (N229)? mem[3073] : 
                       (N231)? mem[3146] : 
                       (N233)? mem[3219] : 
                       (N235)? mem[3292] : 
                       (N237)? mem[3365] : 
                       (N239)? mem[3438] : 
                       (N241)? mem[3511] : 
                       (N243)? mem[3584] : 
                       (N245)? mem[3657] : 
                       (N247)? mem[3730] : 
                       (N249)? mem[3803] : 
                       (N251)? mem[3876] : 
                       (N253)? mem[3949] : 
                       (N255)? mem[4022] : 
                       (N257)? mem[4095] : 
                       (N259)? mem[4168] : 
                       (N261)? mem[4241] : 
                       (N263)? mem[4314] : 
                       (N265)? mem[4387] : 
                       (N267)? mem[4460] : 
                       (N269)? mem[4533] : 
                       (N271)? mem[4606] : 
                       (N146)? mem[4679] : 
                       (N148)? mem[4752] : 
                       (N150)? mem[4825] : 
                       (N152)? mem[4898] : 
                       (N154)? mem[4971] : 
                       (N156)? mem[5044] : 
                       (N158)? mem[5117] : 
                       (N160)? mem[5190] : 
                       (N162)? mem[5263] : 
                       (N164)? mem[5336] : 
                       (N166)? mem[5409] : 
                       (N168)? mem[5482] : 
                       (N170)? mem[5555] : 
                       (N172)? mem[5628] : 
                       (N174)? mem[5701] : 
                       (N176)? mem[5774] : 
                       (N178)? mem[5847] : 
                       (N180)? mem[5920] : 
                       (N182)? mem[5993] : 
                       (N184)? mem[6066] : 
                       (N186)? mem[6139] : 
                       (N188)? mem[6212] : 
                       (N190)? mem[6285] : 
                       (N192)? mem[6358] : 
                       (N194)? mem[6431] : 
                       (N196)? mem[6504] : 
                       (N198)? mem[6577] : 
                       (N200)? mem[6650] : 
                       (N202)? mem[6723] : 
                       (N204)? mem[6796] : 
                       (N206)? mem[6869] : 
                       (N208)? mem[6942] : 
                       (N210)? mem[7015] : 
                       (N212)? mem[7088] : 
                       (N214)? mem[7161] : 
                       (N216)? mem[7234] : 
                       (N218)? mem[7307] : 
                       (N220)? mem[7380] : 
                       (N222)? mem[7453] : 
                       (N224)? mem[7526] : 
                       (N226)? mem[7599] : 
                       (N228)? mem[7672] : 
                       (N230)? mem[7745] : 
                       (N232)? mem[7818] : 
                       (N234)? mem[7891] : 
                       (N236)? mem[7964] : 
                       (N238)? mem[8037] : 
                       (N240)? mem[8110] : 
                       (N242)? mem[8183] : 
                       (N244)? mem[8256] : 
                       (N246)? mem[8329] : 
                       (N248)? mem[8402] : 
                       (N250)? mem[8475] : 
                       (N252)? mem[8548] : 
                       (N254)? mem[8621] : 
                       (N256)? mem[8694] : 
                       (N258)? mem[8767] : 
                       (N260)? mem[8840] : 
                       (N262)? mem[8913] : 
                       (N264)? mem[8986] : 
                       (N266)? mem[9059] : 
                       (N268)? mem[9132] : 
                       (N270)? mem[9205] : 
                       (N272)? mem[9278] : 1'b0;
  assign r_data_o[6] = (N145)? mem[6] : 
                       (N147)? mem[79] : 
                       (N149)? mem[152] : 
                       (N151)? mem[225] : 
                       (N153)? mem[298] : 
                       (N155)? mem[371] : 
                       (N157)? mem[444] : 
                       (N159)? mem[517] : 
                       (N161)? mem[590] : 
                       (N163)? mem[663] : 
                       (N165)? mem[736] : 
                       (N167)? mem[809] : 
                       (N169)? mem[882] : 
                       (N171)? mem[955] : 
                       (N173)? mem[1028] : 
                       (N175)? mem[1101] : 
                       (N177)? mem[1174] : 
                       (N179)? mem[1247] : 
                       (N181)? mem[1320] : 
                       (N183)? mem[1393] : 
                       (N185)? mem[1466] : 
                       (N187)? mem[1539] : 
                       (N189)? mem[1612] : 
                       (N191)? mem[1685] : 
                       (N193)? mem[1758] : 
                       (N195)? mem[1831] : 
                       (N197)? mem[1904] : 
                       (N199)? mem[1977] : 
                       (N201)? mem[2050] : 
                       (N203)? mem[2123] : 
                       (N205)? mem[2196] : 
                       (N207)? mem[2269] : 
                       (N209)? mem[2342] : 
                       (N211)? mem[2415] : 
                       (N213)? mem[2488] : 
                       (N215)? mem[2561] : 
                       (N217)? mem[2634] : 
                       (N219)? mem[2707] : 
                       (N221)? mem[2780] : 
                       (N223)? mem[2853] : 
                       (N225)? mem[2926] : 
                       (N227)? mem[2999] : 
                       (N229)? mem[3072] : 
                       (N231)? mem[3145] : 
                       (N233)? mem[3218] : 
                       (N235)? mem[3291] : 
                       (N237)? mem[3364] : 
                       (N239)? mem[3437] : 
                       (N241)? mem[3510] : 
                       (N243)? mem[3583] : 
                       (N245)? mem[3656] : 
                       (N247)? mem[3729] : 
                       (N249)? mem[3802] : 
                       (N251)? mem[3875] : 
                       (N253)? mem[3948] : 
                       (N255)? mem[4021] : 
                       (N257)? mem[4094] : 
                       (N259)? mem[4167] : 
                       (N261)? mem[4240] : 
                       (N263)? mem[4313] : 
                       (N265)? mem[4386] : 
                       (N267)? mem[4459] : 
                       (N269)? mem[4532] : 
                       (N271)? mem[4605] : 
                       (N146)? mem[4678] : 
                       (N148)? mem[4751] : 
                       (N150)? mem[4824] : 
                       (N152)? mem[4897] : 
                       (N154)? mem[4970] : 
                       (N156)? mem[5043] : 
                       (N158)? mem[5116] : 
                       (N160)? mem[5189] : 
                       (N162)? mem[5262] : 
                       (N164)? mem[5335] : 
                       (N166)? mem[5408] : 
                       (N168)? mem[5481] : 
                       (N170)? mem[5554] : 
                       (N172)? mem[5627] : 
                       (N174)? mem[5700] : 
                       (N176)? mem[5773] : 
                       (N178)? mem[5846] : 
                       (N180)? mem[5919] : 
                       (N182)? mem[5992] : 
                       (N184)? mem[6065] : 
                       (N186)? mem[6138] : 
                       (N188)? mem[6211] : 
                       (N190)? mem[6284] : 
                       (N192)? mem[6357] : 
                       (N194)? mem[6430] : 
                       (N196)? mem[6503] : 
                       (N198)? mem[6576] : 
                       (N200)? mem[6649] : 
                       (N202)? mem[6722] : 
                       (N204)? mem[6795] : 
                       (N206)? mem[6868] : 
                       (N208)? mem[6941] : 
                       (N210)? mem[7014] : 
                       (N212)? mem[7087] : 
                       (N214)? mem[7160] : 
                       (N216)? mem[7233] : 
                       (N218)? mem[7306] : 
                       (N220)? mem[7379] : 
                       (N222)? mem[7452] : 
                       (N224)? mem[7525] : 
                       (N226)? mem[7598] : 
                       (N228)? mem[7671] : 
                       (N230)? mem[7744] : 
                       (N232)? mem[7817] : 
                       (N234)? mem[7890] : 
                       (N236)? mem[7963] : 
                       (N238)? mem[8036] : 
                       (N240)? mem[8109] : 
                       (N242)? mem[8182] : 
                       (N244)? mem[8255] : 
                       (N246)? mem[8328] : 
                       (N248)? mem[8401] : 
                       (N250)? mem[8474] : 
                       (N252)? mem[8547] : 
                       (N254)? mem[8620] : 
                       (N256)? mem[8693] : 
                       (N258)? mem[8766] : 
                       (N260)? mem[8839] : 
                       (N262)? mem[8912] : 
                       (N264)? mem[8985] : 
                       (N266)? mem[9058] : 
                       (N268)? mem[9131] : 
                       (N270)? mem[9204] : 
                       (N272)? mem[9277] : 1'b0;
  assign r_data_o[5] = (N145)? mem[5] : 
                       (N147)? mem[78] : 
                       (N149)? mem[151] : 
                       (N151)? mem[224] : 
                       (N153)? mem[297] : 
                       (N155)? mem[370] : 
                       (N157)? mem[443] : 
                       (N159)? mem[516] : 
                       (N161)? mem[589] : 
                       (N163)? mem[662] : 
                       (N165)? mem[735] : 
                       (N167)? mem[808] : 
                       (N169)? mem[881] : 
                       (N171)? mem[954] : 
                       (N173)? mem[1027] : 
                       (N175)? mem[1100] : 
                       (N177)? mem[1173] : 
                       (N179)? mem[1246] : 
                       (N181)? mem[1319] : 
                       (N183)? mem[1392] : 
                       (N185)? mem[1465] : 
                       (N187)? mem[1538] : 
                       (N189)? mem[1611] : 
                       (N191)? mem[1684] : 
                       (N193)? mem[1757] : 
                       (N195)? mem[1830] : 
                       (N197)? mem[1903] : 
                       (N199)? mem[1976] : 
                       (N201)? mem[2049] : 
                       (N203)? mem[2122] : 
                       (N205)? mem[2195] : 
                       (N207)? mem[2268] : 
                       (N209)? mem[2341] : 
                       (N211)? mem[2414] : 
                       (N213)? mem[2487] : 
                       (N215)? mem[2560] : 
                       (N217)? mem[2633] : 
                       (N219)? mem[2706] : 
                       (N221)? mem[2779] : 
                       (N223)? mem[2852] : 
                       (N225)? mem[2925] : 
                       (N227)? mem[2998] : 
                       (N229)? mem[3071] : 
                       (N231)? mem[3144] : 
                       (N233)? mem[3217] : 
                       (N235)? mem[3290] : 
                       (N237)? mem[3363] : 
                       (N239)? mem[3436] : 
                       (N241)? mem[3509] : 
                       (N243)? mem[3582] : 
                       (N245)? mem[3655] : 
                       (N247)? mem[3728] : 
                       (N249)? mem[3801] : 
                       (N251)? mem[3874] : 
                       (N253)? mem[3947] : 
                       (N255)? mem[4020] : 
                       (N257)? mem[4093] : 
                       (N259)? mem[4166] : 
                       (N261)? mem[4239] : 
                       (N263)? mem[4312] : 
                       (N265)? mem[4385] : 
                       (N267)? mem[4458] : 
                       (N269)? mem[4531] : 
                       (N271)? mem[4604] : 
                       (N146)? mem[4677] : 
                       (N148)? mem[4750] : 
                       (N150)? mem[4823] : 
                       (N152)? mem[4896] : 
                       (N154)? mem[4969] : 
                       (N156)? mem[5042] : 
                       (N158)? mem[5115] : 
                       (N160)? mem[5188] : 
                       (N162)? mem[5261] : 
                       (N164)? mem[5334] : 
                       (N166)? mem[5407] : 
                       (N168)? mem[5480] : 
                       (N170)? mem[5553] : 
                       (N172)? mem[5626] : 
                       (N174)? mem[5699] : 
                       (N176)? mem[5772] : 
                       (N178)? mem[5845] : 
                       (N180)? mem[5918] : 
                       (N182)? mem[5991] : 
                       (N184)? mem[6064] : 
                       (N186)? mem[6137] : 
                       (N188)? mem[6210] : 
                       (N190)? mem[6283] : 
                       (N192)? mem[6356] : 
                       (N194)? mem[6429] : 
                       (N196)? mem[6502] : 
                       (N198)? mem[6575] : 
                       (N200)? mem[6648] : 
                       (N202)? mem[6721] : 
                       (N204)? mem[6794] : 
                       (N206)? mem[6867] : 
                       (N208)? mem[6940] : 
                       (N210)? mem[7013] : 
                       (N212)? mem[7086] : 
                       (N214)? mem[7159] : 
                       (N216)? mem[7232] : 
                       (N218)? mem[7305] : 
                       (N220)? mem[7378] : 
                       (N222)? mem[7451] : 
                       (N224)? mem[7524] : 
                       (N226)? mem[7597] : 
                       (N228)? mem[7670] : 
                       (N230)? mem[7743] : 
                       (N232)? mem[7816] : 
                       (N234)? mem[7889] : 
                       (N236)? mem[7962] : 
                       (N238)? mem[8035] : 
                       (N240)? mem[8108] : 
                       (N242)? mem[8181] : 
                       (N244)? mem[8254] : 
                       (N246)? mem[8327] : 
                       (N248)? mem[8400] : 
                       (N250)? mem[8473] : 
                       (N252)? mem[8546] : 
                       (N254)? mem[8619] : 
                       (N256)? mem[8692] : 
                       (N258)? mem[8765] : 
                       (N260)? mem[8838] : 
                       (N262)? mem[8911] : 
                       (N264)? mem[8984] : 
                       (N266)? mem[9057] : 
                       (N268)? mem[9130] : 
                       (N270)? mem[9203] : 
                       (N272)? mem[9276] : 1'b0;
  assign r_data_o[4] = (N145)? mem[4] : 
                       (N147)? mem[77] : 
                       (N149)? mem[150] : 
                       (N151)? mem[223] : 
                       (N153)? mem[296] : 
                       (N155)? mem[369] : 
                       (N157)? mem[442] : 
                       (N159)? mem[515] : 
                       (N161)? mem[588] : 
                       (N163)? mem[661] : 
                       (N165)? mem[734] : 
                       (N167)? mem[807] : 
                       (N169)? mem[880] : 
                       (N171)? mem[953] : 
                       (N173)? mem[1026] : 
                       (N175)? mem[1099] : 
                       (N177)? mem[1172] : 
                       (N179)? mem[1245] : 
                       (N181)? mem[1318] : 
                       (N183)? mem[1391] : 
                       (N185)? mem[1464] : 
                       (N187)? mem[1537] : 
                       (N189)? mem[1610] : 
                       (N191)? mem[1683] : 
                       (N193)? mem[1756] : 
                       (N195)? mem[1829] : 
                       (N197)? mem[1902] : 
                       (N199)? mem[1975] : 
                       (N201)? mem[2048] : 
                       (N203)? mem[2121] : 
                       (N205)? mem[2194] : 
                       (N207)? mem[2267] : 
                       (N209)? mem[2340] : 
                       (N211)? mem[2413] : 
                       (N213)? mem[2486] : 
                       (N215)? mem[2559] : 
                       (N217)? mem[2632] : 
                       (N219)? mem[2705] : 
                       (N221)? mem[2778] : 
                       (N223)? mem[2851] : 
                       (N225)? mem[2924] : 
                       (N227)? mem[2997] : 
                       (N229)? mem[3070] : 
                       (N231)? mem[3143] : 
                       (N233)? mem[3216] : 
                       (N235)? mem[3289] : 
                       (N237)? mem[3362] : 
                       (N239)? mem[3435] : 
                       (N241)? mem[3508] : 
                       (N243)? mem[3581] : 
                       (N245)? mem[3654] : 
                       (N247)? mem[3727] : 
                       (N249)? mem[3800] : 
                       (N251)? mem[3873] : 
                       (N253)? mem[3946] : 
                       (N255)? mem[4019] : 
                       (N257)? mem[4092] : 
                       (N259)? mem[4165] : 
                       (N261)? mem[4238] : 
                       (N263)? mem[4311] : 
                       (N265)? mem[4384] : 
                       (N267)? mem[4457] : 
                       (N269)? mem[4530] : 
                       (N271)? mem[4603] : 
                       (N146)? mem[4676] : 
                       (N148)? mem[4749] : 
                       (N150)? mem[4822] : 
                       (N152)? mem[4895] : 
                       (N154)? mem[4968] : 
                       (N156)? mem[5041] : 
                       (N158)? mem[5114] : 
                       (N160)? mem[5187] : 
                       (N162)? mem[5260] : 
                       (N164)? mem[5333] : 
                       (N166)? mem[5406] : 
                       (N168)? mem[5479] : 
                       (N170)? mem[5552] : 
                       (N172)? mem[5625] : 
                       (N174)? mem[5698] : 
                       (N176)? mem[5771] : 
                       (N178)? mem[5844] : 
                       (N180)? mem[5917] : 
                       (N182)? mem[5990] : 
                       (N184)? mem[6063] : 
                       (N186)? mem[6136] : 
                       (N188)? mem[6209] : 
                       (N190)? mem[6282] : 
                       (N192)? mem[6355] : 
                       (N194)? mem[6428] : 
                       (N196)? mem[6501] : 
                       (N198)? mem[6574] : 
                       (N200)? mem[6647] : 
                       (N202)? mem[6720] : 
                       (N204)? mem[6793] : 
                       (N206)? mem[6866] : 
                       (N208)? mem[6939] : 
                       (N210)? mem[7012] : 
                       (N212)? mem[7085] : 
                       (N214)? mem[7158] : 
                       (N216)? mem[7231] : 
                       (N218)? mem[7304] : 
                       (N220)? mem[7377] : 
                       (N222)? mem[7450] : 
                       (N224)? mem[7523] : 
                       (N226)? mem[7596] : 
                       (N228)? mem[7669] : 
                       (N230)? mem[7742] : 
                       (N232)? mem[7815] : 
                       (N234)? mem[7888] : 
                       (N236)? mem[7961] : 
                       (N238)? mem[8034] : 
                       (N240)? mem[8107] : 
                       (N242)? mem[8180] : 
                       (N244)? mem[8253] : 
                       (N246)? mem[8326] : 
                       (N248)? mem[8399] : 
                       (N250)? mem[8472] : 
                       (N252)? mem[8545] : 
                       (N254)? mem[8618] : 
                       (N256)? mem[8691] : 
                       (N258)? mem[8764] : 
                       (N260)? mem[8837] : 
                       (N262)? mem[8910] : 
                       (N264)? mem[8983] : 
                       (N266)? mem[9056] : 
                       (N268)? mem[9129] : 
                       (N270)? mem[9202] : 
                       (N272)? mem[9275] : 1'b0;
  assign r_data_o[3] = (N145)? mem[3] : 
                       (N147)? mem[76] : 
                       (N149)? mem[149] : 
                       (N151)? mem[222] : 
                       (N153)? mem[295] : 
                       (N155)? mem[368] : 
                       (N157)? mem[441] : 
                       (N159)? mem[514] : 
                       (N161)? mem[587] : 
                       (N163)? mem[660] : 
                       (N165)? mem[733] : 
                       (N167)? mem[806] : 
                       (N169)? mem[879] : 
                       (N171)? mem[952] : 
                       (N173)? mem[1025] : 
                       (N175)? mem[1098] : 
                       (N177)? mem[1171] : 
                       (N179)? mem[1244] : 
                       (N181)? mem[1317] : 
                       (N183)? mem[1390] : 
                       (N185)? mem[1463] : 
                       (N187)? mem[1536] : 
                       (N189)? mem[1609] : 
                       (N191)? mem[1682] : 
                       (N193)? mem[1755] : 
                       (N195)? mem[1828] : 
                       (N197)? mem[1901] : 
                       (N199)? mem[1974] : 
                       (N201)? mem[2047] : 
                       (N203)? mem[2120] : 
                       (N205)? mem[2193] : 
                       (N207)? mem[2266] : 
                       (N209)? mem[2339] : 
                       (N211)? mem[2412] : 
                       (N213)? mem[2485] : 
                       (N215)? mem[2558] : 
                       (N217)? mem[2631] : 
                       (N219)? mem[2704] : 
                       (N221)? mem[2777] : 
                       (N223)? mem[2850] : 
                       (N225)? mem[2923] : 
                       (N227)? mem[2996] : 
                       (N229)? mem[3069] : 
                       (N231)? mem[3142] : 
                       (N233)? mem[3215] : 
                       (N235)? mem[3288] : 
                       (N237)? mem[3361] : 
                       (N239)? mem[3434] : 
                       (N241)? mem[3507] : 
                       (N243)? mem[3580] : 
                       (N245)? mem[3653] : 
                       (N247)? mem[3726] : 
                       (N249)? mem[3799] : 
                       (N251)? mem[3872] : 
                       (N253)? mem[3945] : 
                       (N255)? mem[4018] : 
                       (N257)? mem[4091] : 
                       (N259)? mem[4164] : 
                       (N261)? mem[4237] : 
                       (N263)? mem[4310] : 
                       (N265)? mem[4383] : 
                       (N267)? mem[4456] : 
                       (N269)? mem[4529] : 
                       (N271)? mem[4602] : 
                       (N146)? mem[4675] : 
                       (N148)? mem[4748] : 
                       (N150)? mem[4821] : 
                       (N152)? mem[4894] : 
                       (N154)? mem[4967] : 
                       (N156)? mem[5040] : 
                       (N158)? mem[5113] : 
                       (N160)? mem[5186] : 
                       (N162)? mem[5259] : 
                       (N164)? mem[5332] : 
                       (N166)? mem[5405] : 
                       (N168)? mem[5478] : 
                       (N170)? mem[5551] : 
                       (N172)? mem[5624] : 
                       (N174)? mem[5697] : 
                       (N176)? mem[5770] : 
                       (N178)? mem[5843] : 
                       (N180)? mem[5916] : 
                       (N182)? mem[5989] : 
                       (N184)? mem[6062] : 
                       (N186)? mem[6135] : 
                       (N188)? mem[6208] : 
                       (N190)? mem[6281] : 
                       (N192)? mem[6354] : 
                       (N194)? mem[6427] : 
                       (N196)? mem[6500] : 
                       (N198)? mem[6573] : 
                       (N200)? mem[6646] : 
                       (N202)? mem[6719] : 
                       (N204)? mem[6792] : 
                       (N206)? mem[6865] : 
                       (N208)? mem[6938] : 
                       (N210)? mem[7011] : 
                       (N212)? mem[7084] : 
                       (N214)? mem[7157] : 
                       (N216)? mem[7230] : 
                       (N218)? mem[7303] : 
                       (N220)? mem[7376] : 
                       (N222)? mem[7449] : 
                       (N224)? mem[7522] : 
                       (N226)? mem[7595] : 
                       (N228)? mem[7668] : 
                       (N230)? mem[7741] : 
                       (N232)? mem[7814] : 
                       (N234)? mem[7887] : 
                       (N236)? mem[7960] : 
                       (N238)? mem[8033] : 
                       (N240)? mem[8106] : 
                       (N242)? mem[8179] : 
                       (N244)? mem[8252] : 
                       (N246)? mem[8325] : 
                       (N248)? mem[8398] : 
                       (N250)? mem[8471] : 
                       (N252)? mem[8544] : 
                       (N254)? mem[8617] : 
                       (N256)? mem[8690] : 
                       (N258)? mem[8763] : 
                       (N260)? mem[8836] : 
                       (N262)? mem[8909] : 
                       (N264)? mem[8982] : 
                       (N266)? mem[9055] : 
                       (N268)? mem[9128] : 
                       (N270)? mem[9201] : 
                       (N272)? mem[9274] : 1'b0;
  assign r_data_o[2] = (N145)? mem[2] : 
                       (N147)? mem[75] : 
                       (N149)? mem[148] : 
                       (N151)? mem[221] : 
                       (N153)? mem[294] : 
                       (N155)? mem[367] : 
                       (N157)? mem[440] : 
                       (N159)? mem[513] : 
                       (N161)? mem[586] : 
                       (N163)? mem[659] : 
                       (N165)? mem[732] : 
                       (N167)? mem[805] : 
                       (N169)? mem[878] : 
                       (N171)? mem[951] : 
                       (N173)? mem[1024] : 
                       (N175)? mem[1097] : 
                       (N177)? mem[1170] : 
                       (N179)? mem[1243] : 
                       (N181)? mem[1316] : 
                       (N183)? mem[1389] : 
                       (N185)? mem[1462] : 
                       (N187)? mem[1535] : 
                       (N189)? mem[1608] : 
                       (N191)? mem[1681] : 
                       (N193)? mem[1754] : 
                       (N195)? mem[1827] : 
                       (N197)? mem[1900] : 
                       (N199)? mem[1973] : 
                       (N201)? mem[2046] : 
                       (N203)? mem[2119] : 
                       (N205)? mem[2192] : 
                       (N207)? mem[2265] : 
                       (N209)? mem[2338] : 
                       (N211)? mem[2411] : 
                       (N213)? mem[2484] : 
                       (N215)? mem[2557] : 
                       (N217)? mem[2630] : 
                       (N219)? mem[2703] : 
                       (N221)? mem[2776] : 
                       (N223)? mem[2849] : 
                       (N225)? mem[2922] : 
                       (N227)? mem[2995] : 
                       (N229)? mem[3068] : 
                       (N231)? mem[3141] : 
                       (N233)? mem[3214] : 
                       (N235)? mem[3287] : 
                       (N237)? mem[3360] : 
                       (N239)? mem[3433] : 
                       (N241)? mem[3506] : 
                       (N243)? mem[3579] : 
                       (N245)? mem[3652] : 
                       (N247)? mem[3725] : 
                       (N249)? mem[3798] : 
                       (N251)? mem[3871] : 
                       (N253)? mem[3944] : 
                       (N255)? mem[4017] : 
                       (N257)? mem[4090] : 
                       (N259)? mem[4163] : 
                       (N261)? mem[4236] : 
                       (N263)? mem[4309] : 
                       (N265)? mem[4382] : 
                       (N267)? mem[4455] : 
                       (N269)? mem[4528] : 
                       (N271)? mem[4601] : 
                       (N146)? mem[4674] : 
                       (N148)? mem[4747] : 
                       (N150)? mem[4820] : 
                       (N152)? mem[4893] : 
                       (N154)? mem[4966] : 
                       (N156)? mem[5039] : 
                       (N158)? mem[5112] : 
                       (N160)? mem[5185] : 
                       (N162)? mem[5258] : 
                       (N164)? mem[5331] : 
                       (N166)? mem[5404] : 
                       (N168)? mem[5477] : 
                       (N170)? mem[5550] : 
                       (N172)? mem[5623] : 
                       (N174)? mem[5696] : 
                       (N176)? mem[5769] : 
                       (N178)? mem[5842] : 
                       (N180)? mem[5915] : 
                       (N182)? mem[5988] : 
                       (N184)? mem[6061] : 
                       (N186)? mem[6134] : 
                       (N188)? mem[6207] : 
                       (N190)? mem[6280] : 
                       (N192)? mem[6353] : 
                       (N194)? mem[6426] : 
                       (N196)? mem[6499] : 
                       (N198)? mem[6572] : 
                       (N200)? mem[6645] : 
                       (N202)? mem[6718] : 
                       (N204)? mem[6791] : 
                       (N206)? mem[6864] : 
                       (N208)? mem[6937] : 
                       (N210)? mem[7010] : 
                       (N212)? mem[7083] : 
                       (N214)? mem[7156] : 
                       (N216)? mem[7229] : 
                       (N218)? mem[7302] : 
                       (N220)? mem[7375] : 
                       (N222)? mem[7448] : 
                       (N224)? mem[7521] : 
                       (N226)? mem[7594] : 
                       (N228)? mem[7667] : 
                       (N230)? mem[7740] : 
                       (N232)? mem[7813] : 
                       (N234)? mem[7886] : 
                       (N236)? mem[7959] : 
                       (N238)? mem[8032] : 
                       (N240)? mem[8105] : 
                       (N242)? mem[8178] : 
                       (N244)? mem[8251] : 
                       (N246)? mem[8324] : 
                       (N248)? mem[8397] : 
                       (N250)? mem[8470] : 
                       (N252)? mem[8543] : 
                       (N254)? mem[8616] : 
                       (N256)? mem[8689] : 
                       (N258)? mem[8762] : 
                       (N260)? mem[8835] : 
                       (N262)? mem[8908] : 
                       (N264)? mem[8981] : 
                       (N266)? mem[9054] : 
                       (N268)? mem[9127] : 
                       (N270)? mem[9200] : 
                       (N272)? mem[9273] : 1'b0;
  assign r_data_o[1] = (N145)? mem[1] : 
                       (N147)? mem[74] : 
                       (N149)? mem[147] : 
                       (N151)? mem[220] : 
                       (N153)? mem[293] : 
                       (N155)? mem[366] : 
                       (N157)? mem[439] : 
                       (N159)? mem[512] : 
                       (N161)? mem[585] : 
                       (N163)? mem[658] : 
                       (N165)? mem[731] : 
                       (N167)? mem[804] : 
                       (N169)? mem[877] : 
                       (N171)? mem[950] : 
                       (N173)? mem[1023] : 
                       (N175)? mem[1096] : 
                       (N177)? mem[1169] : 
                       (N179)? mem[1242] : 
                       (N181)? mem[1315] : 
                       (N183)? mem[1388] : 
                       (N185)? mem[1461] : 
                       (N187)? mem[1534] : 
                       (N189)? mem[1607] : 
                       (N191)? mem[1680] : 
                       (N193)? mem[1753] : 
                       (N195)? mem[1826] : 
                       (N197)? mem[1899] : 
                       (N199)? mem[1972] : 
                       (N201)? mem[2045] : 
                       (N203)? mem[2118] : 
                       (N205)? mem[2191] : 
                       (N207)? mem[2264] : 
                       (N209)? mem[2337] : 
                       (N211)? mem[2410] : 
                       (N213)? mem[2483] : 
                       (N215)? mem[2556] : 
                       (N217)? mem[2629] : 
                       (N219)? mem[2702] : 
                       (N221)? mem[2775] : 
                       (N223)? mem[2848] : 
                       (N225)? mem[2921] : 
                       (N227)? mem[2994] : 
                       (N229)? mem[3067] : 
                       (N231)? mem[3140] : 
                       (N233)? mem[3213] : 
                       (N235)? mem[3286] : 
                       (N237)? mem[3359] : 
                       (N239)? mem[3432] : 
                       (N241)? mem[3505] : 
                       (N243)? mem[3578] : 
                       (N245)? mem[3651] : 
                       (N247)? mem[3724] : 
                       (N249)? mem[3797] : 
                       (N251)? mem[3870] : 
                       (N253)? mem[3943] : 
                       (N255)? mem[4016] : 
                       (N257)? mem[4089] : 
                       (N259)? mem[4162] : 
                       (N261)? mem[4235] : 
                       (N263)? mem[4308] : 
                       (N265)? mem[4381] : 
                       (N267)? mem[4454] : 
                       (N269)? mem[4527] : 
                       (N271)? mem[4600] : 
                       (N146)? mem[4673] : 
                       (N148)? mem[4746] : 
                       (N150)? mem[4819] : 
                       (N152)? mem[4892] : 
                       (N154)? mem[4965] : 
                       (N156)? mem[5038] : 
                       (N158)? mem[5111] : 
                       (N160)? mem[5184] : 
                       (N162)? mem[5257] : 
                       (N164)? mem[5330] : 
                       (N166)? mem[5403] : 
                       (N168)? mem[5476] : 
                       (N170)? mem[5549] : 
                       (N172)? mem[5622] : 
                       (N174)? mem[5695] : 
                       (N176)? mem[5768] : 
                       (N178)? mem[5841] : 
                       (N180)? mem[5914] : 
                       (N182)? mem[5987] : 
                       (N184)? mem[6060] : 
                       (N186)? mem[6133] : 
                       (N188)? mem[6206] : 
                       (N190)? mem[6279] : 
                       (N192)? mem[6352] : 
                       (N194)? mem[6425] : 
                       (N196)? mem[6498] : 
                       (N198)? mem[6571] : 
                       (N200)? mem[6644] : 
                       (N202)? mem[6717] : 
                       (N204)? mem[6790] : 
                       (N206)? mem[6863] : 
                       (N208)? mem[6936] : 
                       (N210)? mem[7009] : 
                       (N212)? mem[7082] : 
                       (N214)? mem[7155] : 
                       (N216)? mem[7228] : 
                       (N218)? mem[7301] : 
                       (N220)? mem[7374] : 
                       (N222)? mem[7447] : 
                       (N224)? mem[7520] : 
                       (N226)? mem[7593] : 
                       (N228)? mem[7666] : 
                       (N230)? mem[7739] : 
                       (N232)? mem[7812] : 
                       (N234)? mem[7885] : 
                       (N236)? mem[7958] : 
                       (N238)? mem[8031] : 
                       (N240)? mem[8104] : 
                       (N242)? mem[8177] : 
                       (N244)? mem[8250] : 
                       (N246)? mem[8323] : 
                       (N248)? mem[8396] : 
                       (N250)? mem[8469] : 
                       (N252)? mem[8542] : 
                       (N254)? mem[8615] : 
                       (N256)? mem[8688] : 
                       (N258)? mem[8761] : 
                       (N260)? mem[8834] : 
                       (N262)? mem[8907] : 
                       (N264)? mem[8980] : 
                       (N266)? mem[9053] : 
                       (N268)? mem[9126] : 
                       (N270)? mem[9199] : 
                       (N272)? mem[9272] : 1'b0;
  assign r_data_o[0] = (N145)? mem[0] : 
                       (N147)? mem[73] : 
                       (N149)? mem[146] : 
                       (N151)? mem[219] : 
                       (N153)? mem[292] : 
                       (N155)? mem[365] : 
                       (N157)? mem[438] : 
                       (N159)? mem[511] : 
                       (N161)? mem[584] : 
                       (N163)? mem[657] : 
                       (N165)? mem[730] : 
                       (N167)? mem[803] : 
                       (N169)? mem[876] : 
                       (N171)? mem[949] : 
                       (N173)? mem[1022] : 
                       (N175)? mem[1095] : 
                       (N177)? mem[1168] : 
                       (N179)? mem[1241] : 
                       (N181)? mem[1314] : 
                       (N183)? mem[1387] : 
                       (N185)? mem[1460] : 
                       (N187)? mem[1533] : 
                       (N189)? mem[1606] : 
                       (N191)? mem[1679] : 
                       (N193)? mem[1752] : 
                       (N195)? mem[1825] : 
                       (N197)? mem[1898] : 
                       (N199)? mem[1971] : 
                       (N201)? mem[2044] : 
                       (N203)? mem[2117] : 
                       (N205)? mem[2190] : 
                       (N207)? mem[2263] : 
                       (N209)? mem[2336] : 
                       (N211)? mem[2409] : 
                       (N213)? mem[2482] : 
                       (N215)? mem[2555] : 
                       (N217)? mem[2628] : 
                       (N219)? mem[2701] : 
                       (N221)? mem[2774] : 
                       (N223)? mem[2847] : 
                       (N225)? mem[2920] : 
                       (N227)? mem[2993] : 
                       (N229)? mem[3066] : 
                       (N231)? mem[3139] : 
                       (N233)? mem[3212] : 
                       (N235)? mem[3285] : 
                       (N237)? mem[3358] : 
                       (N239)? mem[3431] : 
                       (N241)? mem[3504] : 
                       (N243)? mem[3577] : 
                       (N245)? mem[3650] : 
                       (N247)? mem[3723] : 
                       (N249)? mem[3796] : 
                       (N251)? mem[3869] : 
                       (N253)? mem[3942] : 
                       (N255)? mem[4015] : 
                       (N257)? mem[4088] : 
                       (N259)? mem[4161] : 
                       (N261)? mem[4234] : 
                       (N263)? mem[4307] : 
                       (N265)? mem[4380] : 
                       (N267)? mem[4453] : 
                       (N269)? mem[4526] : 
                       (N271)? mem[4599] : 
                       (N146)? mem[4672] : 
                       (N148)? mem[4745] : 
                       (N150)? mem[4818] : 
                       (N152)? mem[4891] : 
                       (N154)? mem[4964] : 
                       (N156)? mem[5037] : 
                       (N158)? mem[5110] : 
                       (N160)? mem[5183] : 
                       (N162)? mem[5256] : 
                       (N164)? mem[5329] : 
                       (N166)? mem[5402] : 
                       (N168)? mem[5475] : 
                       (N170)? mem[5548] : 
                       (N172)? mem[5621] : 
                       (N174)? mem[5694] : 
                       (N176)? mem[5767] : 
                       (N178)? mem[5840] : 
                       (N180)? mem[5913] : 
                       (N182)? mem[5986] : 
                       (N184)? mem[6059] : 
                       (N186)? mem[6132] : 
                       (N188)? mem[6205] : 
                       (N190)? mem[6278] : 
                       (N192)? mem[6351] : 
                       (N194)? mem[6424] : 
                       (N196)? mem[6497] : 
                       (N198)? mem[6570] : 
                       (N200)? mem[6643] : 
                       (N202)? mem[6716] : 
                       (N204)? mem[6789] : 
                       (N206)? mem[6862] : 
                       (N208)? mem[6935] : 
                       (N210)? mem[7008] : 
                       (N212)? mem[7081] : 
                       (N214)? mem[7154] : 
                       (N216)? mem[7227] : 
                       (N218)? mem[7300] : 
                       (N220)? mem[7373] : 
                       (N222)? mem[7446] : 
                       (N224)? mem[7519] : 
                       (N226)? mem[7592] : 
                       (N228)? mem[7665] : 
                       (N230)? mem[7738] : 
                       (N232)? mem[7811] : 
                       (N234)? mem[7884] : 
                       (N236)? mem[7957] : 
                       (N238)? mem[8030] : 
                       (N240)? mem[8103] : 
                       (N242)? mem[8176] : 
                       (N244)? mem[8249] : 
                       (N246)? mem[8322] : 
                       (N248)? mem[8395] : 
                       (N250)? mem[8468] : 
                       (N252)? mem[8541] : 
                       (N254)? mem[8614] : 
                       (N256)? mem[8687] : 
                       (N258)? mem[8760] : 
                       (N260)? mem[8833] : 
                       (N262)? mem[8906] : 
                       (N264)? mem[8979] : 
                       (N266)? mem[9052] : 
                       (N268)? mem[9125] : 
                       (N270)? mem[9198] : 
                       (N272)? mem[9271] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9343] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9342] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9341] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9340] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9339] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9338] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9337] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9336] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9335] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9334] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9333] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9332] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9331] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9330] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9329] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9328] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9327] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9326] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9325] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9324] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9323] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9322] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9321] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9320] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9319] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9318] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9317] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9316] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9315] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9314] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9313] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9312] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9311] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9310] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9309] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9308] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9307] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9306] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9305] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9304] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9303] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9302] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9301] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9300] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9299] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9298] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9297] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9296] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9295] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9294] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9293] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9292] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9291] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9290] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9289] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9288] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9287] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9286] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9285] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9284] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9283] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9282] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9281] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9280] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9279] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9278] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9277] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9276] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9275] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9274] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9273] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9272] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N529) begin
      mem[9271] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9270] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9269] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9268] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9267] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9266] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9265] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9264] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9263] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9262] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9261] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9260] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9259] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9258] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9257] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9256] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9255] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9254] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9253] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9252] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9251] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9250] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9249] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9248] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9247] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9246] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9245] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9244] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9243] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9242] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9241] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9240] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9239] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9238] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9237] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9236] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9235] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9234] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9233] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9232] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9231] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9230] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9229] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9228] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9227] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9226] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9225] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9224] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9223] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9222] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9221] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9220] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9219] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9218] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9217] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9216] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9215] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9214] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9213] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9212] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9211] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9210] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9209] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9208] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9207] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9206] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9205] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9204] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9203] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9202] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9201] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9200] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9199] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N528) begin
      mem[9198] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9197] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9196] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9195] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9194] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9193] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9192] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9191] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9190] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9189] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9188] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9187] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9186] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9185] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9184] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9183] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9182] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9181] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9180] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9179] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9178] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9177] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9176] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9175] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9174] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9173] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9172] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9171] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9170] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9169] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9168] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9167] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9166] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9165] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9164] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9163] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9162] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9161] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9160] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9159] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9158] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9157] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9156] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9155] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9154] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9153] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9152] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9151] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9150] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9149] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9148] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9147] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9146] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9145] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9144] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9143] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9142] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9141] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9140] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9139] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9138] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9137] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9136] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9135] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9134] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9133] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9132] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9131] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9130] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9129] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9128] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9127] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9126] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N527) begin
      mem[9125] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9124] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9123] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9122] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9121] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9120] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9119] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9118] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9117] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9116] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9115] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9114] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9113] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9112] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9111] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9110] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9109] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9108] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9107] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9106] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9105] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9104] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9103] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9102] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9101] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9100] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9099] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9098] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9097] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9096] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9095] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9094] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9093] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9092] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9091] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9090] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9089] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9088] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9087] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9086] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9085] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9084] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9083] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9082] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9081] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9080] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9079] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9078] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9077] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9076] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9075] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9074] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9073] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9072] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9071] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9070] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9069] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9068] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9067] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9066] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9065] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9064] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9063] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9062] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9061] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9060] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9059] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9058] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9057] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9056] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9055] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9054] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9053] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N526) begin
      mem[9052] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9051] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9050] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9049] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9048] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9047] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9046] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9045] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9044] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9043] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9042] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9041] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9040] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9039] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9038] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9037] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9036] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9035] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9034] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9033] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9032] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9031] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9030] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9029] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9028] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9027] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9026] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9025] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9024] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9023] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9022] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9021] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9020] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9019] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9018] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9017] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9016] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9015] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9014] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9013] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9012] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9011] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9010] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9009] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9008] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9007] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9006] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9005] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9004] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9003] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9002] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9001] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[9000] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8999] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8998] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8997] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8996] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8995] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8994] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8993] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8992] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8991] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8990] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8989] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8988] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8987] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8986] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8985] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8984] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8983] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8982] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8981] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8980] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N525) begin
      mem[8979] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8978] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8977] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8976] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8975] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8974] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8973] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8972] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8971] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8970] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8969] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8968] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8967] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8966] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8965] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8964] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8963] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8962] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8961] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8960] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8959] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8958] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8957] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8956] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8955] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8954] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8953] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8952] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8951] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8950] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8949] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8948] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8947] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8946] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8945] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8944] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8943] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8942] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8941] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8940] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8939] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8938] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8937] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8936] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8935] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8934] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8933] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8932] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8931] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8930] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8929] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8928] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8927] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8926] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8925] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8924] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8923] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8922] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8921] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8920] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8919] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8918] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8917] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8916] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8915] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8914] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8913] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8912] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8911] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8910] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8909] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8908] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8907] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N524) begin
      mem[8906] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8905] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8904] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8903] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8902] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8901] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8900] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8899] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8898] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8897] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8896] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8895] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8894] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8893] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8892] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8891] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8890] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8889] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8888] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8887] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8886] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8885] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8884] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8883] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8882] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8881] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8880] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8879] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8878] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8877] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8876] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8875] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8874] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8873] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8872] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8871] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8870] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8869] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8868] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8867] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8866] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8865] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8864] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8863] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8862] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8861] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8860] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8859] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8858] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8857] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8856] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8855] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8854] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8853] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8852] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8851] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8850] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8849] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8848] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8847] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8846] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8845] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8844] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8843] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8842] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8841] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8840] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8839] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8838] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8837] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8836] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8835] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8834] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N523) begin
      mem[8833] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8832] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8831] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8830] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8829] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8828] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8827] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8826] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8825] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8824] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8823] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8822] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8821] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8820] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8819] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8818] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8817] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8816] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8815] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8814] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8813] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8812] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8811] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8810] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8809] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8808] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8807] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8806] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8805] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8804] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8803] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8802] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8801] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8800] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8799] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8798] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8797] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8796] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8795] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8794] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8793] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8792] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8791] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8790] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8789] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8788] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8787] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8786] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8785] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8784] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8783] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8782] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8781] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8780] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8779] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8778] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8777] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8776] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8775] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8774] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8773] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8772] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8771] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8770] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8769] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8768] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8767] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8766] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8765] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8764] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8763] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8762] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8761] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N522) begin
      mem[8760] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8759] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8758] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8757] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8756] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8755] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8754] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8753] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8752] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8751] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8750] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8749] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8748] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8747] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8746] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8745] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8744] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8743] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8742] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8741] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8740] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8739] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8738] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8737] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8736] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8735] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8734] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8733] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8732] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8731] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8730] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8729] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8728] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8727] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8726] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8725] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8724] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8723] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8722] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8721] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8720] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8719] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8718] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8717] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8716] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8715] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8714] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8713] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8712] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8711] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8710] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8709] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8708] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8707] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8706] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8705] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8704] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8703] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8702] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8701] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8700] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8699] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8698] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8697] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8696] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8695] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8694] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8693] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8692] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8691] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8690] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8689] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8688] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N521) begin
      mem[8687] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8686] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8685] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8684] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8683] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8682] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8681] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8680] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8679] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8678] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8677] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8676] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8675] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8674] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8673] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8672] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8671] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8670] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8669] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8668] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8667] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8666] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8665] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8664] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8663] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8662] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8661] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8660] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8659] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8658] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8657] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8656] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8655] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8654] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8653] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8652] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8651] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8650] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8649] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8648] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8647] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8646] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8645] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8644] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8643] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8642] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8641] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8640] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8639] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8638] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8637] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8636] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8635] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8634] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8633] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8632] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8631] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8630] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8629] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8628] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8627] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8626] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8625] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8624] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8623] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8622] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8621] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8620] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8619] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8618] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8617] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8616] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8615] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N520) begin
      mem[8614] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8613] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8612] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8611] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8610] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8609] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8608] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8607] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8606] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8605] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8604] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8603] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8602] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8601] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8600] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8599] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8598] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8597] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8596] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8595] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8594] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8593] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8592] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8591] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8590] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8589] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8588] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8587] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8586] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8585] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8584] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8583] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8582] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8581] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8580] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8579] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8578] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8577] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8576] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8575] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8574] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8573] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8572] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8571] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8570] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8569] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8568] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8567] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8566] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8565] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8564] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8563] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8562] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8561] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8560] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8559] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8558] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8557] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8556] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8555] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8554] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8553] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8552] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8551] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8550] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8549] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8548] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8547] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8546] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8545] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8544] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8543] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8542] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N519) begin
      mem[8541] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8540] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8539] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8538] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8537] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8536] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8535] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8534] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8533] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8532] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8531] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8530] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8529] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8528] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8527] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8526] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8525] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8524] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8523] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8522] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8521] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8520] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8519] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8518] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8517] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8516] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8515] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8514] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8513] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8512] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8511] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8510] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8509] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8508] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8507] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8506] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8505] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8504] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8503] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8502] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8501] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8500] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8499] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8498] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8497] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8496] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8495] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8494] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8493] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8492] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8491] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8490] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8489] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8488] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8487] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8486] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8485] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8484] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8483] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8482] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8481] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8480] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8479] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8478] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8477] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8476] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8475] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8474] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8473] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8472] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8471] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8470] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8469] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N518) begin
      mem[8468] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8467] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8466] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8465] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8464] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8463] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8462] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8461] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8460] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8459] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8458] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8457] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8456] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8455] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8454] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8453] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8452] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8451] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8450] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8449] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8448] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8447] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8446] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8445] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8444] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8443] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8442] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8441] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8440] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8439] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8438] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8437] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8436] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8435] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8434] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8433] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8432] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8431] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8430] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8429] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8428] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8427] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8426] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8425] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8424] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8423] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8422] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8421] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8420] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8419] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8418] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8417] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8416] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8415] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8414] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8413] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8412] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8411] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8410] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8409] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8408] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8407] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8406] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8405] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8404] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8403] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8402] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8401] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8400] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8399] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8398] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8397] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8396] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N517) begin
      mem[8395] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8394] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8393] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8392] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8391] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8390] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8389] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8388] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8387] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8386] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8385] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8384] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8383] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8382] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8381] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8380] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8379] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8378] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8377] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8376] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8375] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8374] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8373] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8372] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8371] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8370] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8369] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8368] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8367] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8366] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8365] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8364] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8363] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8362] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8361] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8360] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8359] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8358] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8357] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8356] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8355] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8354] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8353] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8352] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8351] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8350] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8349] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8348] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8347] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8346] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8345] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8344] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8343] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8342] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8341] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8340] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8339] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8338] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8337] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8336] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8335] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8334] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8333] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8332] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8331] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8330] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8329] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8328] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8327] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8326] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8325] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8324] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8323] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N516) begin
      mem[8322] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8321] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8320] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8319] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8318] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8317] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8316] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8315] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8314] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8313] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8312] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8311] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8310] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8309] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8308] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8307] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8306] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8305] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8304] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8303] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8302] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8301] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8300] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8299] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8298] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8297] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8296] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8295] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8294] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8293] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8292] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8291] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8290] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8289] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8288] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8287] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8286] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8285] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8284] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8283] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8282] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8281] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8280] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8279] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8278] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8277] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8276] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8275] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8274] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8273] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8272] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8271] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8270] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8269] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8268] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8267] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8266] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8265] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8264] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8263] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8262] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8261] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8260] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8259] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8258] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8257] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8256] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8255] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8254] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8253] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8252] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8251] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8250] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N515) begin
      mem[8249] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8248] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8247] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8246] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8245] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8244] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8243] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8242] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8241] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8240] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8239] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8238] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8237] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8236] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8235] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8234] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8233] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8232] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8231] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8230] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8229] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8228] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8227] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8226] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8225] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8224] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8223] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8222] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8221] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8220] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8219] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8218] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8217] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8216] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8215] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8214] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8213] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8212] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8211] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8210] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8209] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8208] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8207] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8206] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8205] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8204] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8203] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8202] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8201] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8200] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8199] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8198] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8197] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8196] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8195] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8194] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8193] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8192] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8191] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8190] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8189] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8188] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8187] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8186] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8185] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8184] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8183] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8182] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8181] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8180] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8179] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8178] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8177] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N514) begin
      mem[8176] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8175] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8174] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8173] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8172] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8171] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8170] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8169] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8168] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8167] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8166] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8165] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8164] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8163] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8162] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8161] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8160] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8159] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8158] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8157] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8156] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8155] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8154] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8153] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8152] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8151] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8150] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8149] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8148] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8147] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8146] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8145] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8144] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8143] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8142] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8141] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8140] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8139] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8138] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8137] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8136] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8135] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8134] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8133] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8132] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8131] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8130] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8129] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8128] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8127] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8126] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8125] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8124] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8123] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8122] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8121] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8120] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8119] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8118] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8117] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8116] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8115] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8114] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8113] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8112] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8111] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8110] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8109] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8108] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8107] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8106] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8105] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8104] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N513) begin
      mem[8103] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8102] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8101] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8100] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8099] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8098] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8097] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8096] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8095] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8094] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8093] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8092] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8091] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8090] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8089] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8088] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8087] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8086] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8085] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8084] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8083] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8082] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8081] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8080] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8079] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8078] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8077] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8076] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8075] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8074] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8073] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8072] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8071] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8070] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8069] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8068] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8067] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8066] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8065] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8064] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8063] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8062] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8061] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8060] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8059] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8058] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8057] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8056] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8055] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8054] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8053] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8052] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8051] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8050] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8049] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8048] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8047] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8046] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8045] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8044] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8043] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8042] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8041] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8040] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8039] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8038] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8037] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8036] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8035] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8034] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8033] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8032] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8031] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N512) begin
      mem[8030] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8029] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8028] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8027] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8026] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8025] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8024] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8023] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8022] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8021] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8020] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8019] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8018] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8017] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8016] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8015] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8014] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8013] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8012] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8011] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8010] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8009] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8008] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8007] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8006] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8005] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8004] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8003] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8002] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8001] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[8000] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7999] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7998] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7997] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7996] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7995] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7994] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7993] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7992] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7991] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7990] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7989] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7988] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7987] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7986] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7985] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7984] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7983] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7982] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7981] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7980] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7979] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7978] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7977] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7976] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7975] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7974] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7973] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7972] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7971] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7970] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7969] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7968] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7967] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7966] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7965] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7964] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7963] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7962] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7961] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7960] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7959] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7958] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N511) begin
      mem[7957] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7956] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7955] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7954] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7953] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7952] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7951] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7950] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7949] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7948] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7947] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7946] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7945] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7944] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7943] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7942] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7941] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7940] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7939] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7938] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7937] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7936] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7935] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7934] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7933] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7932] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7931] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7930] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7929] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7928] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7927] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7926] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7925] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7924] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7923] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7922] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7921] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7920] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7919] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7918] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7917] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7916] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7915] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7914] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7913] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7912] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7911] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7910] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7909] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7908] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7907] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7906] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7905] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7904] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7903] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7902] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7901] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7900] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7899] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7898] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7897] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7896] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7895] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7894] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7893] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7892] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7891] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7890] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7889] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7888] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7887] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7886] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7885] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N510) begin
      mem[7884] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7883] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7882] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7881] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7880] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7879] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7878] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7877] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7876] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7875] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7874] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7873] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7872] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7871] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7870] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7869] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7868] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7867] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7866] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7865] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7864] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7863] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7862] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7861] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7860] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7859] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7858] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7857] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7856] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7855] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7854] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7853] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7852] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7851] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7850] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7849] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7848] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7847] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7846] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7845] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7844] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7843] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7842] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7841] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7840] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7839] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7838] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7837] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7836] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7835] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7834] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7833] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7832] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7831] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7830] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7829] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7828] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7827] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7826] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7825] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7824] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7823] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7822] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7821] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7820] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7819] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7818] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7817] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7816] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7815] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7814] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7813] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7812] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N509) begin
      mem[7811] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7810] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7809] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7808] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7807] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7806] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7805] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7804] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7803] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7802] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7801] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7800] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7799] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7798] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7797] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7796] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7795] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7794] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7793] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7792] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7791] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7790] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7789] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7788] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7787] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7786] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7785] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7784] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7783] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7782] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7781] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7780] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7779] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7778] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7777] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7776] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7775] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7774] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7773] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7772] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7771] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7770] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7769] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7768] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7767] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7766] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7765] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7764] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7763] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7762] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7761] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7760] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7759] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7758] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7757] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7756] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7755] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7754] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7753] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7752] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7751] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7750] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7749] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7748] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7747] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7746] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7745] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7744] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7743] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7742] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7741] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7740] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7739] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N508) begin
      mem[7738] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7737] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7736] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7735] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7734] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7733] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7732] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7731] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7730] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7729] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7728] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7727] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7726] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7725] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7724] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7723] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7722] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7721] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7720] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7719] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7718] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7717] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7716] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7715] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7714] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7713] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7712] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7711] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7710] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7709] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7708] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7707] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7706] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7705] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7704] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7703] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7702] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7701] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7700] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7699] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7698] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7697] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7696] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7695] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7694] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7693] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7692] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7691] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7690] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7689] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7688] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7687] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7686] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7685] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7684] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7683] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7682] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7681] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7680] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7679] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7678] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7677] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7676] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7675] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7674] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7673] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7672] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7671] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7670] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7669] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7668] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7667] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7666] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N507) begin
      mem[7665] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7664] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7663] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7662] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7661] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7660] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7659] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7658] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7657] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7656] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7655] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7654] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7653] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7652] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7651] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7650] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7649] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7648] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7647] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7646] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7645] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7644] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7643] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7642] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7641] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7640] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7639] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7638] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7637] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7636] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7635] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7634] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7633] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7632] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7631] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7630] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7629] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7628] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7627] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7626] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7625] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7624] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7623] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7622] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7621] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7620] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7619] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7618] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7617] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7616] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7615] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7614] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7613] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7612] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7611] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7610] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7609] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7608] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7607] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7606] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7605] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7604] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7603] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7602] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7601] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7600] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7599] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7598] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7597] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7596] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7595] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7594] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7593] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N506) begin
      mem[7592] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7591] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7590] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7589] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7588] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7587] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7586] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7585] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7584] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7583] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7582] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7581] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7580] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7579] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7578] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7577] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7576] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7575] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7574] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7573] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7572] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7571] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7570] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7569] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7568] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7567] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7566] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7565] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7564] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7563] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7562] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7561] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7560] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7559] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7558] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7557] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7556] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7555] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7554] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7553] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7552] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7551] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7550] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7549] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7548] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7547] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7546] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7545] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7544] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7543] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7542] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7541] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7540] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7539] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7538] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7537] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7536] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7535] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7534] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7533] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7532] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7531] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7530] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7529] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7528] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7527] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7526] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7525] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7524] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7523] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7522] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7521] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7520] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N505) begin
      mem[7519] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7518] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7517] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7516] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7515] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7514] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7513] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7512] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7511] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7510] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7509] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7508] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7507] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7506] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7505] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7504] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7503] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7502] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7501] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7500] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7499] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7498] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7497] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7496] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7495] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7494] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7493] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7492] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7491] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7490] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7489] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7488] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7487] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7486] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7485] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7484] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7483] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7482] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7481] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7480] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7479] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7478] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7477] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7476] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7475] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7474] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7473] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7472] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7471] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7470] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7469] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7468] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7467] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7466] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7465] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7464] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7463] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7462] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7461] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7460] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7459] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7458] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7457] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7456] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7455] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7454] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7453] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7452] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7451] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7450] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7449] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7448] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7447] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N504) begin
      mem[7446] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7445] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7444] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7443] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7442] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7441] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7440] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7439] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7438] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7437] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7436] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7435] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7434] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7433] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7432] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7431] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7430] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7429] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7428] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7427] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7426] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7425] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7424] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7423] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7422] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7421] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7420] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7419] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7418] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7417] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7416] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7415] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7414] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7413] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7412] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7411] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7410] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7409] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7408] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7407] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7406] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7405] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7404] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7403] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7402] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7401] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7400] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7399] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7398] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7397] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7396] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7395] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7394] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7393] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7392] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7391] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7390] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7389] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7388] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7387] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7386] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7385] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7384] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7383] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7382] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7381] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7380] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7379] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7378] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7377] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7376] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7375] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7374] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N503) begin
      mem[7373] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7372] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7371] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7370] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7369] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7368] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7367] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7366] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7365] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7364] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7363] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7362] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7361] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7360] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7359] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7358] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7357] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7356] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7355] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7354] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7353] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7352] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7351] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7350] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7349] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7348] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7347] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7346] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7345] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7344] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7343] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7342] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7341] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7340] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7339] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7338] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7337] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7336] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7335] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7334] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7333] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7332] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7331] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7330] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7329] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7328] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7327] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7326] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7325] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7324] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7323] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7322] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7321] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7320] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7319] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7318] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7317] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7316] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7315] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7314] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7313] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7312] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7311] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7310] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7309] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7308] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7307] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7306] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7305] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7304] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7303] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7302] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7301] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N502) begin
      mem[7300] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7299] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7298] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7297] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7296] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7295] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7294] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7293] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7292] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7291] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7290] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7289] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7288] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7287] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7286] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7285] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7284] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7283] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7282] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7281] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7280] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7279] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7278] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7277] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7276] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7275] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7274] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7273] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7272] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7271] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7270] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7269] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7268] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7267] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7266] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7265] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7264] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7263] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7262] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7261] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7260] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7259] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7258] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7257] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7256] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7255] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7254] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7253] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7252] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7251] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7250] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7249] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7248] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7247] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7246] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7245] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7244] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7243] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7242] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7241] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7240] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7239] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7238] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7237] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7236] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7235] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7234] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7233] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7232] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7231] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7230] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7229] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7228] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N501) begin
      mem[7227] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7226] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7225] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7224] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7223] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7222] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7221] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7220] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7219] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7218] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7217] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7216] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7215] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7214] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7213] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7212] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7211] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7210] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7209] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7208] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7207] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7206] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7205] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7204] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7203] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7202] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7201] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7200] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7199] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7198] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7197] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7196] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7195] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7194] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7193] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7192] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7191] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7190] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7189] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7188] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7187] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7186] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7185] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7184] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7183] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7182] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7181] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7180] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7179] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7178] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7177] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7176] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7175] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7174] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7173] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7172] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7171] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7170] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7169] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7168] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7167] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7166] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7165] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7164] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7163] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7162] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7161] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7160] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7159] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7158] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7157] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7156] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7155] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N500) begin
      mem[7154] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7153] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7152] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7151] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7150] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7149] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7148] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7147] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7146] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7145] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7144] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7143] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7142] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7141] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7140] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7139] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7138] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7137] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7136] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7135] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7134] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7133] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7132] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7131] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7130] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7129] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7128] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7127] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7126] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7125] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7124] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7123] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7122] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7121] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7120] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7119] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7118] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7117] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7116] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7115] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7114] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7113] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7112] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7111] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7110] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7109] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7108] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7107] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7106] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7105] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7104] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7103] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7102] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7101] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7100] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7099] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7098] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7097] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7096] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7095] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7094] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7093] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7092] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7091] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7090] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7089] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7088] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7087] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7086] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7085] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7084] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7083] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7082] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N499) begin
      mem[7081] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7080] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7079] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7078] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7077] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7076] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7075] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7074] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7073] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7072] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7071] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7070] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7069] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7068] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7067] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7066] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7065] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7064] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7063] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7062] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7061] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7060] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7059] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7058] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7057] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7056] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7055] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7054] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7053] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7052] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7051] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7050] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7049] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7048] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7047] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7046] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7045] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7044] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7043] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7042] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7041] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7040] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7039] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7038] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7037] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7036] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7035] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7034] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7033] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7032] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7031] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7030] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7029] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7028] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7027] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7026] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7025] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7024] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7023] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7022] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7021] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7020] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7019] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7018] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7017] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7016] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7015] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7014] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7013] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7012] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7011] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7010] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7009] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N498) begin
      mem[7008] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7007] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7006] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7005] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7004] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7003] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7002] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7001] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[7000] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6999] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6998] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6997] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6996] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6995] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6994] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6993] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6992] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6991] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6990] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6989] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6988] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6987] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6986] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6985] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6984] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6983] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6982] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6981] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6980] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6979] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6978] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6977] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6976] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6975] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6974] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6973] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6972] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6971] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6970] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6969] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6968] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6967] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6966] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6965] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6964] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6963] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6962] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6961] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6960] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6959] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6958] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6957] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6956] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6955] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6954] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6953] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6952] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6951] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6950] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6949] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6948] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6947] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6946] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6945] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6944] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6943] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6942] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6941] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6940] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6939] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6938] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6937] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6936] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N497) begin
      mem[6935] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6934] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6933] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6932] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6931] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6930] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6929] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6928] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6927] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6926] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6925] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6924] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6923] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6922] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6921] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6920] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6919] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6918] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6917] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6916] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6915] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6914] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6913] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6912] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6911] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6910] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6909] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6908] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6907] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6906] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6905] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6904] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6903] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6902] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6901] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6900] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6899] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6898] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6897] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6896] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6895] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6894] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6893] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6892] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6891] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6890] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6889] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6888] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6887] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6886] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6885] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6884] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6883] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6882] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6881] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6880] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6879] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6878] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6877] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6876] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6875] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6874] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6873] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6872] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6871] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6870] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6869] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6868] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6867] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6866] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6865] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6864] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6863] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N496) begin
      mem[6862] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6861] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6860] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6859] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6858] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6857] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6856] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6855] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6854] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6853] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6852] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6851] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6850] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6849] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6848] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6847] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6846] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6845] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6844] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6843] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6842] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6841] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6840] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6839] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6838] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6837] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6836] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6835] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6834] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6833] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6832] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6831] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6830] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6829] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6828] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6827] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6826] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6825] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6824] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6823] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6822] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6821] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6820] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6819] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6818] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6817] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6816] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6815] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6814] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6813] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6812] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6811] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6810] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6809] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6808] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6807] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6806] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6805] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6804] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6803] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6802] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6801] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6800] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6799] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6798] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6797] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6796] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6795] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6794] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6793] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6792] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6791] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6790] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N495) begin
      mem[6789] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6788] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6787] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6786] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6785] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6784] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6783] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6782] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6781] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6780] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6779] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6778] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6777] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6776] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6775] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6774] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6773] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6772] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6771] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6770] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6769] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6768] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6767] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6766] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6765] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6764] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6763] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6762] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6761] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6760] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6759] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6758] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6757] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6756] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6755] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6754] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6753] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6752] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6751] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6750] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6749] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6748] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6747] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6746] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6745] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6744] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6743] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6742] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6741] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6740] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6739] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6738] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6737] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6736] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6735] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6734] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6733] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6732] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6731] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6730] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6729] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6728] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6727] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6726] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6725] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6724] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6723] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6722] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6721] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6720] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6719] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6718] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6717] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N494) begin
      mem[6716] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6715] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6714] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6713] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6712] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6711] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6710] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6709] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6708] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6707] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6706] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6705] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6704] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6703] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6702] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6701] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6700] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6699] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6698] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6697] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6696] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6695] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6694] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6693] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6692] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6691] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6690] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6689] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6688] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6687] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6686] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6685] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6684] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6683] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6682] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6681] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6680] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6679] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6678] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6677] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6676] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6675] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6674] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6673] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6672] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6671] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6670] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6669] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6668] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6667] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6666] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6665] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6664] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6663] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6662] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6661] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6660] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6659] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6658] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6657] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6656] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6655] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6654] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6653] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6652] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6651] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6650] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6649] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6648] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6647] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6646] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6645] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6644] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N493) begin
      mem[6643] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6642] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6641] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6640] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6639] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6638] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6637] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6636] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6635] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6634] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6633] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6632] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6631] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6630] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6629] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6628] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6627] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6626] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6625] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6624] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6623] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6622] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6621] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6620] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6619] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6618] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6617] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6616] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6615] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6614] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6613] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6612] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6611] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6610] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6609] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6608] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6607] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6606] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6605] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6604] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6603] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6602] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6601] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6600] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6599] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6598] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6597] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6596] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6595] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6594] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6593] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6592] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6591] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6590] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6589] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6588] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6587] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6586] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6585] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6584] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6583] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6582] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6581] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6580] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6579] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6578] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6577] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6576] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6575] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6574] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6573] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6572] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6571] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N492) begin
      mem[6570] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6569] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6568] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6567] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6566] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6565] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6564] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6563] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6562] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6561] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6560] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6559] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6558] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6557] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6556] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6555] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6554] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6553] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6552] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6551] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6550] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6549] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6548] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6547] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6546] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6545] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6544] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6543] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6542] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6541] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6540] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6539] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6538] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6537] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6536] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6535] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6534] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6533] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6532] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6531] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6530] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6529] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6528] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6527] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6526] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6525] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6524] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6523] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6522] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6521] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6520] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6519] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6518] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6517] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6516] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6515] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6514] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6513] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6512] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6511] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6510] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6509] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6508] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6507] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6506] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6505] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6504] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6503] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6502] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6501] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6500] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6499] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6498] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N491) begin
      mem[6497] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6496] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6495] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6494] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6493] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6492] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6491] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6490] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6489] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6488] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6487] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6486] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6485] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6484] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6483] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6482] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6481] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6480] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6479] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6478] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6477] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6476] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6475] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6474] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6473] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6472] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6471] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6470] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6469] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6468] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6467] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6466] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6465] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6464] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6463] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6462] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6461] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6460] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6459] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6458] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6457] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6456] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6455] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6454] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6453] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6452] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6451] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6450] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6449] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6448] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6447] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6446] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6445] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6444] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6443] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6442] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6441] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6440] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6439] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6438] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6437] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6436] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6435] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6434] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6433] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6432] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6431] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6430] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6429] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6428] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6427] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6426] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6425] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N490) begin
      mem[6424] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6423] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6422] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6421] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6420] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6419] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6418] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6417] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6416] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6415] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6414] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6413] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6412] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6411] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6410] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6409] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6408] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6407] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6406] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6405] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6404] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6403] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6402] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6401] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6400] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6399] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6398] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6397] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6396] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6395] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6394] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6393] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6392] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6391] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6390] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6389] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6388] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6387] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6386] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6385] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6384] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6383] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6382] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6381] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6380] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6379] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6378] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6377] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6376] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6375] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6374] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6373] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6372] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6371] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6370] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6369] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6368] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6367] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6366] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6365] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6364] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6363] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6362] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6361] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6360] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6359] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6358] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6357] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6356] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6355] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6354] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6353] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6352] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N489) begin
      mem[6351] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6350] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6349] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6348] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6347] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6346] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6345] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6344] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6343] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6342] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6341] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6340] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6339] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6338] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6337] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6336] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6335] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6334] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6333] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6332] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6331] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6330] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6329] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6328] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6327] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6326] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6325] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6324] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6323] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6322] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6321] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6320] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6319] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6318] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6317] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6316] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6315] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6314] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6313] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6312] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6311] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6310] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6309] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6308] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6307] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6306] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6305] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6304] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6303] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6302] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6301] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6300] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6299] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6298] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6297] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6296] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6295] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6294] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6293] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6292] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6291] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6290] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6289] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6288] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6287] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6286] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6285] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6284] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6283] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6282] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6281] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6280] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6279] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N488) begin
      mem[6278] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6277] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6276] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6275] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6274] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6273] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6272] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6271] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6270] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6269] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6268] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6267] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6266] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6265] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6264] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6263] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6262] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6261] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6260] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6259] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6258] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6257] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6256] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6255] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6254] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6253] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6252] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6251] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6250] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6249] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6248] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6247] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6246] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6245] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6244] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6243] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6242] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6241] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6240] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6239] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6238] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6237] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6236] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6235] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6234] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6233] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6232] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6231] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6230] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6229] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6228] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6227] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6226] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6225] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6224] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6223] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6222] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6221] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6220] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6219] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6218] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6217] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6216] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6215] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6214] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6213] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6212] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6211] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6210] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6209] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6208] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6207] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6206] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N487) begin
      mem[6205] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6204] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6203] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6202] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6201] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6200] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6199] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6198] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6197] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6196] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6195] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6194] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6193] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6192] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6191] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6190] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6189] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6188] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6187] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6186] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6185] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6184] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6183] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6182] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6181] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6180] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6179] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6178] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6177] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6176] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6175] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6174] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6173] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6172] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6171] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6170] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6169] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6168] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6167] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6166] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6165] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6164] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6163] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6162] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6161] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6160] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6159] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6158] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6157] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6156] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6155] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6154] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6153] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6152] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6151] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6150] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6149] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6148] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6147] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6146] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6145] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6144] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6143] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6142] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6141] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6140] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6139] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6138] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6137] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6136] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6135] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6134] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6133] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N486) begin
      mem[6132] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6131] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6130] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6129] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6128] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6127] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6126] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6125] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6124] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6123] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6122] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6121] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6120] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6119] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6118] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6117] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6116] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6115] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6114] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6113] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6112] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6111] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6110] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6109] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6108] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6107] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6106] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6105] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6104] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6103] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6102] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6101] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6100] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6099] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6098] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6097] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6096] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6095] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6094] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6093] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6092] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6091] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6090] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6089] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6088] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6087] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6086] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6085] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6084] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6083] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6082] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6081] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6080] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6079] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6078] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6077] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6076] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6075] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6074] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6073] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6072] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6071] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6070] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6069] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6068] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6067] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6066] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6065] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6064] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6063] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6062] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6061] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6060] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N485) begin
      mem[6059] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6058] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6057] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6056] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6055] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6054] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6053] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6052] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6051] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6050] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6049] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6048] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6047] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6046] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6045] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6044] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6043] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6042] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6041] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6040] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6039] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6038] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6037] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6036] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6035] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6034] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6033] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6032] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6031] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6030] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6029] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6028] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6027] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6026] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6025] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6024] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6023] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6022] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6021] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6020] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6019] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6018] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6017] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6016] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6015] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6014] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6013] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6012] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6011] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6010] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6009] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6008] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6007] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6006] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6005] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6004] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6003] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6002] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6001] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[6000] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5999] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5998] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5997] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5996] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5995] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5994] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5993] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5992] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5991] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5990] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5989] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5988] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5987] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N484) begin
      mem[5986] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5985] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5984] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5983] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5982] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5981] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5980] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5979] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5978] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5977] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5976] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5975] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5974] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5973] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5972] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5971] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5970] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5969] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5968] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5967] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5966] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5965] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5964] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5963] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5962] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5961] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5960] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5959] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5958] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5957] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5956] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5955] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5954] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5953] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5952] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5951] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5950] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5949] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5948] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5947] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5946] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5945] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5944] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5943] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5942] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5941] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5940] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5939] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5938] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5937] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5936] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5935] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5934] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5933] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5932] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5931] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5930] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5929] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5928] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5927] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5926] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5925] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5924] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5923] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5922] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5921] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5920] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5919] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5918] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5917] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5916] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5915] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5914] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N483) begin
      mem[5913] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5912] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5911] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5910] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5909] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5908] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5907] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5906] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5905] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5904] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5903] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5902] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5901] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5900] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5899] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5898] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5897] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5896] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5895] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5894] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5893] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5892] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5891] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5890] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5889] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5888] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5887] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5886] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5885] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5884] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5883] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5882] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5881] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5880] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5879] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5878] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5877] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5876] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5875] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5874] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5873] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5872] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5871] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5870] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5869] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5868] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5867] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5866] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5865] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5864] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5863] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5862] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5861] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5860] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5859] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5858] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5857] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5856] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5855] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5854] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5853] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5852] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5851] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5850] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5849] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5848] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5847] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5846] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5845] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5844] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5843] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5842] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5841] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N482) begin
      mem[5840] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5839] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5838] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5837] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5836] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5835] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5834] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5833] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5832] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5831] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5830] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5829] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5828] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5827] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5826] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5825] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5824] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5823] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5822] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5821] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5820] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5819] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5818] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5817] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5816] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5815] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5814] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5813] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5812] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5811] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5810] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5809] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5808] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5807] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5806] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5805] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5804] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5803] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5802] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5801] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5800] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5799] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5798] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5797] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5796] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5795] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5794] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5793] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5792] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5791] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5790] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5789] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5788] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5787] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5786] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5785] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5784] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5783] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5782] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5781] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5780] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5779] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5778] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5777] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5776] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5775] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5774] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5773] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5772] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5771] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5770] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5769] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5768] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N481) begin
      mem[5767] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5766] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5765] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5764] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5763] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5762] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5761] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5760] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5759] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5758] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5757] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5756] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5755] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5754] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5753] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5752] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5751] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5750] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5749] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5748] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5747] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5746] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5745] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5744] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5743] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5742] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5741] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5740] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5739] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5738] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5737] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5736] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5735] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5734] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5733] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5732] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5731] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5730] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5729] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5728] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5727] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5726] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5725] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5724] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5723] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5722] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5721] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5720] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5719] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5718] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5717] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5716] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5715] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5714] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5713] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5712] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5711] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5710] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5709] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5708] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5707] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5706] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5705] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5704] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5703] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5702] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5701] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5700] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5699] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5698] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5697] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5696] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5695] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N480) begin
      mem[5694] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5693] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5692] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5691] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5690] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5689] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5688] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5687] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5686] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5685] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5684] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5683] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5682] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5681] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5680] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5679] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5678] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5677] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5676] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5675] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5674] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5673] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5672] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5671] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5670] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5669] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5668] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5667] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5666] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5665] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5664] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5663] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5662] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5661] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5660] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5659] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5658] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5657] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5656] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5655] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5654] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5653] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5652] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5651] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5650] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5649] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5648] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5647] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5646] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5645] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5644] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5643] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5642] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5641] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5640] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5639] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5638] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5637] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5636] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5635] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5634] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5633] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5632] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5631] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5630] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5629] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5628] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5627] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5626] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5625] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5624] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5623] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5622] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N479) begin
      mem[5621] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5620] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5619] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5618] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5617] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5616] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5615] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5614] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5613] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5612] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5611] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5610] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5609] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5608] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5607] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5606] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5605] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5604] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5603] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5602] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5601] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5600] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5599] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5598] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5597] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5596] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5595] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5594] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5593] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5592] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5591] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5590] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5589] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5588] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5587] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5586] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5585] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5584] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5583] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5582] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5581] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5580] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5579] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5578] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5577] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5576] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5575] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5574] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5573] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5572] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5571] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5570] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5569] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5568] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5567] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5566] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5565] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5564] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5563] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5562] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5561] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5560] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5559] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5558] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5557] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5556] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5555] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5554] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5553] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5552] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5551] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5550] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5549] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N478) begin
      mem[5548] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5547] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5546] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5545] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5544] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5543] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5542] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5541] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5540] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5539] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5538] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5537] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5536] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5535] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5534] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5533] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5532] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5531] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5530] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5529] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5528] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5527] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5526] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5525] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5524] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5523] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5522] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5521] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5520] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5519] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5518] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5517] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5516] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5515] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5514] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5513] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5512] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5511] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5510] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5509] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5508] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5507] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5506] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5505] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5504] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5503] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5502] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5501] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5500] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5499] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5498] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5497] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5496] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5495] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5494] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5493] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5492] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5491] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5490] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5489] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5488] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5487] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5486] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5485] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5484] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5483] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5482] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5481] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5480] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5479] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5478] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5477] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5476] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N477) begin
      mem[5475] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5474] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5473] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5472] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5471] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5470] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5469] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5468] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5467] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5466] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5465] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5464] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5463] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5462] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5461] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5460] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5459] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5458] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5457] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5456] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5455] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5454] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5453] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5452] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5451] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5450] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5449] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5448] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5447] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5446] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5445] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5444] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5443] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5442] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5441] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5440] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5439] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5438] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5437] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5436] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5435] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5434] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5433] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5432] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5431] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5430] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5429] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5428] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5427] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5426] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5425] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5424] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5423] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5422] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5421] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5420] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5419] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5418] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5417] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5416] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5415] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5414] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5413] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5412] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5411] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5410] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5409] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5408] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5407] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5406] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5405] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5404] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5403] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N476) begin
      mem[5402] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5401] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5400] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5399] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5398] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5397] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5396] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5395] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5394] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5393] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5392] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5391] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5390] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5389] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5388] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5387] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5386] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5385] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5384] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5383] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5382] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5381] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5380] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5379] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5378] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5377] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5376] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5375] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5374] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5373] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5372] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5371] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5370] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5369] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5368] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5367] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5366] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5365] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5364] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5363] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5362] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5361] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5360] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5359] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5358] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5357] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5356] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5355] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5354] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5353] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5352] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5351] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5350] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5349] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5348] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5347] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5346] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5345] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5344] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5343] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5342] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5341] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5340] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5339] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5338] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5337] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5336] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5335] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5334] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5333] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5332] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5331] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5330] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N475) begin
      mem[5329] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5328] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5327] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5326] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5325] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5324] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5323] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5322] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5321] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5320] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5319] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5318] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5317] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5316] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5315] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5314] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5313] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5312] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5311] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5310] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5309] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5308] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5307] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5306] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5305] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5304] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5303] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5302] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5301] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5300] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5299] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5298] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5297] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5296] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5295] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5294] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5293] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5292] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5291] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5290] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5289] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5288] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5287] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5286] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5285] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5284] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5283] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5282] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5281] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5280] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5279] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5278] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5277] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5276] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5275] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5274] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5273] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5272] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5271] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5270] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5269] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5268] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5267] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5266] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5265] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5264] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5263] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5262] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5261] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5260] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5259] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5258] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5257] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N474) begin
      mem[5256] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5255] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5254] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5253] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5252] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5251] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5250] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5249] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5248] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5247] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5246] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5245] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5244] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5243] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5242] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5241] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5240] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5239] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5238] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5237] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5236] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5235] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5234] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5233] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5232] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5231] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5230] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5229] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5228] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5227] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5226] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5225] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5224] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5223] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5222] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5221] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5220] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5219] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5218] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5217] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5216] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5215] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5214] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5213] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5212] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5211] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5210] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5209] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5208] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5207] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5206] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5205] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5204] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5203] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5202] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5201] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5200] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5199] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5198] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5197] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5196] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5195] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5194] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5193] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5192] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5191] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5190] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5189] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5188] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5187] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5186] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5185] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5184] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N473) begin
      mem[5183] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5182] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5181] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5180] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5179] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5178] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5177] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5176] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5175] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5174] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5173] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5172] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5171] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5170] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5169] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5168] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5167] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5166] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5165] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5164] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5163] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5162] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5161] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5160] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5159] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5158] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5157] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5156] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5155] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5154] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5153] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5152] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5151] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5150] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5149] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5148] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5147] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5146] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5145] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5144] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5143] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5142] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5141] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5140] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5139] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5138] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5137] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5136] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5135] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5134] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5133] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5132] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5131] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5130] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5129] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5128] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5127] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5126] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5125] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5124] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5123] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5122] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5121] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5120] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5119] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5118] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5117] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5116] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5115] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5114] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5113] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5112] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5111] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N472) begin
      mem[5110] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5109] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5108] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5107] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5106] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5105] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5104] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5103] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5102] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5101] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5100] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5099] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5098] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5097] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5096] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5095] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5094] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5093] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5092] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5091] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5090] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5089] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5088] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5087] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5086] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5085] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5084] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5083] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5082] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5081] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5080] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5079] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5078] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5077] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5076] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5075] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5074] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5073] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5072] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5071] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5070] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5069] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5068] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5067] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5066] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5065] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5064] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5063] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5062] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5061] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5060] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5059] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5058] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5057] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5056] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5055] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5054] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5053] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5052] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5051] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5050] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5049] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5048] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5047] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5046] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5045] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5044] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5043] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5042] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5041] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5040] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5039] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5038] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N471) begin
      mem[5037] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5036] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5035] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5034] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5033] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5032] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5031] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5030] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5029] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5028] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5027] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5026] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5025] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5024] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5023] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5022] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5021] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5020] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5019] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5018] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5017] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5016] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5015] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5014] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5013] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5012] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5011] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5010] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5009] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5008] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5007] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5006] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5005] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5004] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5003] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5002] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5001] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[5000] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4999] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4998] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4997] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4996] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4995] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4994] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4993] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4992] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4991] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4990] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4989] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4988] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4987] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4986] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4985] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4984] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4983] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4982] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4981] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4980] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4979] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4978] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4977] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4976] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4975] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4974] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4973] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4972] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4971] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4970] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4969] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4968] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4967] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4966] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4965] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N470) begin
      mem[4964] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4963] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4962] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4961] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4960] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4959] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4958] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4957] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4956] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4955] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4954] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4953] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4952] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4951] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4950] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4949] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4948] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4947] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4946] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4945] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4944] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4943] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4942] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4941] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4940] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4939] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4938] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4937] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4936] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4935] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4934] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4933] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4932] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4931] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4930] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4929] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4928] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4927] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4926] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4925] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4924] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4923] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4922] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4921] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4920] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4919] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4918] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4917] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4916] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4915] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4914] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4913] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4912] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4911] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4910] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4909] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4908] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4907] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4906] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4905] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4904] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4903] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4902] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4901] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4900] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4899] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4898] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4897] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4896] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4895] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4894] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4893] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4892] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N469) begin
      mem[4891] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4890] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4889] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4888] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4887] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4886] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4885] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4884] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4883] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4882] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4881] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4880] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4879] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4878] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4877] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4876] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4875] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4874] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4873] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4872] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4871] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4870] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4869] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4868] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4867] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4866] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4865] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4864] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4863] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4862] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4861] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4860] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4859] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4858] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4857] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4856] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4855] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4854] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4853] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4852] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4851] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4850] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4849] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4848] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4847] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4846] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4845] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4844] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4843] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4842] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4841] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4840] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4839] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4838] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4837] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4836] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4835] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4834] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4833] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4832] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4831] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4830] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4829] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4828] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4827] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4826] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4825] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4824] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4823] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4822] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4821] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4820] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4819] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N468) begin
      mem[4818] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4817] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4816] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4815] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4814] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4813] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4812] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4811] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4810] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4809] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4808] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4807] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4806] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4805] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4804] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4803] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4802] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4801] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4800] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4799] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4798] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4797] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4796] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4795] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4794] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4793] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4792] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4791] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4790] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4789] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4788] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4787] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4786] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4785] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4784] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4783] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4782] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4781] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4780] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4779] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4778] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4777] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4776] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4775] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4774] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4773] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4772] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4771] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4770] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4769] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4768] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4767] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4766] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4765] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4764] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4763] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4762] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4761] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4760] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4759] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4758] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4757] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4756] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4755] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4754] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4753] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4752] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4751] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4750] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4749] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4748] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4747] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4746] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N467) begin
      mem[4745] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4744] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4743] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4742] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4741] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4740] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4739] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4738] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4737] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4736] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4735] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4734] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4733] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4732] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4731] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4730] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4729] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4728] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4727] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4726] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4725] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4724] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4723] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4722] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4721] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4720] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4719] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4718] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4717] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4716] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4715] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4714] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4713] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4712] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4711] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4710] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4709] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4708] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4707] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4706] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4705] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4704] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4703] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4702] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4701] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4700] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4699] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4698] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4697] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4696] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4695] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4694] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4693] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4692] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4691] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4690] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4689] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4688] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4687] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4686] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4685] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4684] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4683] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4682] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4681] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4680] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4679] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4678] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4677] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4676] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4675] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4674] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4673] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N466) begin
      mem[4672] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4671] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4670] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4669] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4668] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4667] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4666] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4665] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4664] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4663] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4662] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4661] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4660] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4659] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4658] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4657] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4656] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4655] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4654] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4653] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4652] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4651] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4650] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4649] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4648] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4647] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4646] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4645] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4644] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4643] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4642] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4641] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4640] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4639] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4638] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4637] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4636] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4635] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4634] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4633] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4632] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4631] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4630] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4629] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4628] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4627] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4626] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4625] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4624] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4623] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4622] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4621] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4620] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4619] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4618] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4617] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4616] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4615] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4614] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4613] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4612] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4611] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4610] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4609] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4608] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4607] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4606] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4605] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4604] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4603] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4602] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4601] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4600] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N465) begin
      mem[4599] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4598] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4597] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4596] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4595] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4594] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4593] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4592] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4591] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4590] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4589] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4588] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4587] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4586] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4585] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4584] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4583] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4582] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4581] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4580] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4579] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4578] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4577] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4576] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4575] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4574] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4573] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4572] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4571] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4570] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4569] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4568] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4567] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4566] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4565] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4564] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4563] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4562] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4561] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4560] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4559] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4558] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4557] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4556] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4555] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4554] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4553] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4552] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4551] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4550] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4549] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4548] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4547] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4546] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4545] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4544] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4543] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4542] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4541] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4540] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4539] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4538] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4537] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4536] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4535] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4534] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4533] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4532] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4531] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4530] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4529] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4528] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4527] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N464) begin
      mem[4526] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4525] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4524] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4523] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4522] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4521] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4520] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4519] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4518] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4517] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4516] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4515] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4514] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4513] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4512] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4511] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4510] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4509] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4508] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4507] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4506] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4505] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4504] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4503] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4502] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4501] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4500] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4499] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4498] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4497] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4496] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4495] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4494] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4493] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4492] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4491] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4490] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4489] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4488] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4487] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4486] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4485] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4484] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4483] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4482] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4481] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4480] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4479] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4478] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4477] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4476] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4475] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4474] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4473] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4472] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4471] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4470] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4469] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4468] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4467] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4466] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4465] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4464] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4463] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4462] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4461] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4460] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4459] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4458] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4457] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4456] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4455] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4454] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N463) begin
      mem[4453] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4452] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4451] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4450] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4449] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4448] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4447] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4446] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4445] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4444] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4443] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4442] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4441] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4440] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4439] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4438] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4437] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4436] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4435] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4434] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4433] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4432] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4431] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4430] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4429] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4428] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4427] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4426] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4425] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4424] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4423] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4422] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4421] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4420] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4419] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4418] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4417] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4416] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4415] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4414] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4413] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4412] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4411] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4410] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4409] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4408] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4407] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4406] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4405] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4404] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4403] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4402] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4401] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4400] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4399] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4398] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4397] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4396] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4395] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4394] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4393] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4392] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4391] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4390] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4389] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4388] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4387] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4386] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4385] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4384] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4383] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4382] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4381] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N462) begin
      mem[4380] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4379] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4378] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4377] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4376] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4375] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4374] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4373] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4372] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4371] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4370] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4369] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4368] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4367] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4366] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4365] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4364] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4363] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4362] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4361] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4360] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4359] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4358] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4357] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4356] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4355] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4354] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4353] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4352] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4351] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4350] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4349] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4348] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4347] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4346] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4345] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4344] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4343] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4342] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4341] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4340] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4339] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4338] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4337] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4336] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4335] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4334] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4333] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4332] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4331] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4330] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4329] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4328] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4327] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4326] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4325] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4324] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4323] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4322] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4321] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4320] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4319] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4318] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4317] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4316] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4315] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4314] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4313] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4312] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4311] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4310] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4309] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4308] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N461) begin
      mem[4307] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4306] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4305] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4304] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4303] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4302] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4301] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4300] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4299] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4298] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4297] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4296] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4295] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4294] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4293] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4292] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4291] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4290] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4289] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4288] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4287] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4286] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4285] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4284] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4283] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4282] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4281] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4280] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4279] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4278] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4277] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4276] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4275] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4274] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4273] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4272] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4271] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4270] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4269] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4268] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4267] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4266] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4265] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4264] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4263] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4262] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4261] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4260] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4259] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4258] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4257] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4256] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4255] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4254] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4253] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4252] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4251] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4250] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4249] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4248] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4247] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4246] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4245] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4244] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4243] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4242] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4241] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4240] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4239] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4238] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4237] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4236] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4235] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N460) begin
      mem[4234] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4233] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4232] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4231] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4230] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4229] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4228] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4227] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4226] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4225] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4224] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4223] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4222] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4221] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4220] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4219] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4218] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4217] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4216] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4215] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4214] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4213] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4212] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4211] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4210] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4209] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4208] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4207] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4206] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4205] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4204] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4203] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4202] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4201] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4200] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4199] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4198] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4197] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4196] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4195] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4194] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4193] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4192] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4191] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4190] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4189] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4188] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4187] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4186] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4185] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4184] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4183] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4182] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4181] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4180] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4179] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4178] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4177] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4176] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4175] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4174] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4173] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4172] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4171] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4170] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4169] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4168] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4167] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4166] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4165] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4164] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4163] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4162] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N459) begin
      mem[4161] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4160] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4159] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4158] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4157] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4156] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4155] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4154] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4153] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4152] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4151] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4150] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4149] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4148] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4147] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4146] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4145] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4144] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4143] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4142] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4141] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4140] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4139] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4138] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4137] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4136] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4135] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4134] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4133] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4132] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4131] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4130] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4129] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4128] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4127] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4126] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4125] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4124] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4123] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4122] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4121] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4120] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4119] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4118] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4117] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4116] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4115] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4114] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4113] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4112] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4111] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4110] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4109] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4108] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4107] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4106] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4105] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4104] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4103] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4102] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4101] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4100] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4099] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4098] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4097] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4096] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4095] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4094] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4093] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4092] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4091] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4090] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4089] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N458) begin
      mem[4088] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4087] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4086] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4085] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4084] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4083] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4082] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4081] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4080] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4079] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4078] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4077] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4076] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4075] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4074] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4073] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4072] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4071] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4070] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4069] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4068] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4067] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4066] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4065] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4064] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4063] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4062] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4061] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4060] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4059] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4058] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4057] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4056] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4055] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4054] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4053] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4052] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4051] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4050] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4049] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4048] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4047] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4046] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4045] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4044] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4043] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4042] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4041] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4040] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4039] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4038] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4037] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4036] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4035] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4034] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4033] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4032] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4031] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4030] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4029] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4028] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4027] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4026] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4025] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4024] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4023] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4022] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4021] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4020] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4019] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4018] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4017] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4016] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N457) begin
      mem[4015] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4014] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4013] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4012] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4011] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4010] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4009] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4008] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4007] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4006] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4005] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4004] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4003] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4002] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4001] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[4000] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3999] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3998] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3997] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3996] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3995] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3994] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3993] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3992] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3991] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3990] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3989] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3988] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3987] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3986] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3985] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3984] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3983] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3982] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3981] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3980] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3979] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3978] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3977] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3976] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3975] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3974] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3973] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3972] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3971] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3970] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3969] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3968] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3967] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3966] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3965] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3964] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3963] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3962] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3961] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3960] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3959] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3958] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3957] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3956] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3955] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3954] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3953] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3952] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3951] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3950] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3949] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3948] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3947] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3946] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3945] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3944] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3943] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N456) begin
      mem[3942] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3941] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3940] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3939] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3938] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3937] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3936] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3935] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3934] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3933] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3932] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3931] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3930] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3929] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3928] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3927] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3926] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3925] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3924] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3923] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3922] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3921] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3920] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3919] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3918] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3917] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3916] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3915] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3914] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3913] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3912] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3911] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3910] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3909] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3908] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3907] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3906] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3905] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3904] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3903] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3902] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3901] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3900] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3899] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3898] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3897] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3896] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3895] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3894] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3893] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3892] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3891] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3890] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3889] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3888] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3887] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3886] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3885] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3884] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3883] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3882] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3881] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3880] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3879] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3878] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3877] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3876] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3875] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3874] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3873] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3872] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3871] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3870] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N455) begin
      mem[3869] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3868] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3867] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3866] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3865] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3864] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3863] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3862] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3861] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3860] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3859] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3858] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3857] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3856] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3855] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3854] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3853] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3852] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3851] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3850] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3849] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3848] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3847] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3846] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3845] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3844] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3843] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3842] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3841] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3840] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3839] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3838] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3837] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3836] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3835] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3834] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3833] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3832] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3831] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3830] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3829] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3828] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3827] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3826] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3825] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3824] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3823] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3822] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3821] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3820] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3819] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3818] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3817] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3816] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3815] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3814] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3813] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3812] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3811] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3810] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3809] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3808] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3807] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3806] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3805] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3804] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3803] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3802] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3801] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3800] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3799] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3798] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3797] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N454) begin
      mem[3796] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3795] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3794] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3793] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3792] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3791] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3790] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3789] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3788] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3787] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3786] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3785] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3784] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3783] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3782] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3781] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3780] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3779] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3778] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3777] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3776] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3775] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3774] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3773] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3772] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3771] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3770] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3769] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3768] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3767] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3766] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3765] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3764] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3763] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3762] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3761] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3760] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3759] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3758] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3757] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3756] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3755] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3754] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3753] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3752] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3751] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3750] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3749] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3748] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3747] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3746] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3745] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3744] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3743] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3742] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3741] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3740] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3739] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3738] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3737] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3736] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3735] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3734] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3733] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3732] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3731] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3730] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3729] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3728] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3727] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3726] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3725] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3724] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N453) begin
      mem[3723] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3722] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3721] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3720] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3719] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3718] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3717] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3716] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3715] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3714] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3713] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3712] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3711] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3710] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3709] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3708] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3707] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3706] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3705] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3704] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3703] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3702] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3701] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3700] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3699] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3698] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3697] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3696] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3695] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3694] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3693] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3692] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3691] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3690] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3689] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3688] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3687] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3686] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3685] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3684] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3683] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3682] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3681] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3680] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3679] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3678] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3677] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3676] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3675] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3674] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3673] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3672] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3671] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3670] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3669] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3668] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3667] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3666] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3665] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3664] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3663] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3662] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3661] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3660] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3659] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3658] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3657] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3656] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3655] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3654] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3653] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3652] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3651] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N452) begin
      mem[3650] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3649] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3648] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3647] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3646] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3645] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3644] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3643] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3642] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3641] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3640] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3639] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3638] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3637] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3636] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3635] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3634] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3633] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3632] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3631] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3630] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3629] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3628] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3627] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3626] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3625] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3624] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3623] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3622] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3621] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3620] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3619] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3618] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3617] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3616] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3615] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3614] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3613] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3612] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3611] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3610] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3609] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3608] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3607] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3606] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3605] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3604] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3603] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3602] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3601] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3600] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3599] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3598] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3597] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3596] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3595] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3594] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3593] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3592] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3591] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3590] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3589] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3588] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3587] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3586] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3585] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3584] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3583] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3582] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3581] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3580] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3579] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3578] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N451) begin
      mem[3577] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3576] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3575] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3574] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3573] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3572] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3571] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3570] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3569] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3568] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3567] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3566] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3565] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3564] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3563] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3562] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3561] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3560] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3559] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3558] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3557] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3556] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3555] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3554] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3553] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3552] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3551] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3550] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3549] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3548] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3547] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3546] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3545] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3544] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3543] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3542] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3541] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3540] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3539] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3538] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3537] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3536] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3535] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3534] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3533] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3532] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3531] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3530] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3529] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3528] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3527] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3526] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3525] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3524] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3523] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3522] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3521] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3520] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3519] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3518] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3517] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3516] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3515] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3514] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3513] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3512] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3511] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3510] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3509] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3508] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3507] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3506] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3505] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N450) begin
      mem[3504] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3503] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3502] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3501] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3500] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3499] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3498] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3497] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3496] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3495] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3494] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3493] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3492] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3491] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3490] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3489] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3488] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3487] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3486] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3485] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3484] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3483] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3482] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3481] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3480] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3479] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3478] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3477] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3476] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3475] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3474] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3473] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3472] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3471] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3470] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3469] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3468] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3467] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3466] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3465] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3464] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3463] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3462] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3461] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3460] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3459] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3458] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3457] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3456] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3455] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3454] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3453] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3452] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3451] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3450] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3449] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3448] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3447] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3446] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3445] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3444] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3443] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3442] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3441] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3440] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3439] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3438] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3437] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3436] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3435] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3434] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3433] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3432] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N449) begin
      mem[3431] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3430] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3429] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3428] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3427] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3426] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3425] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3424] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3423] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3422] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3421] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3420] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3419] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3418] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3417] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3416] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3415] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3414] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3413] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3412] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3411] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3410] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3409] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3408] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3407] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3406] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3405] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3404] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3403] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3402] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3401] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3400] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3399] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3398] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3397] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3396] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3395] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3394] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3393] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3392] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3391] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3390] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3389] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3388] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3387] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3386] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3385] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3384] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3383] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3382] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3381] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3380] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3379] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3378] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3377] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3376] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3375] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3374] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3373] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3372] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3371] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3370] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3369] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3368] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3367] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3366] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3365] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3364] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3363] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3362] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3361] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3360] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3359] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N448) begin
      mem[3358] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3357] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3356] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3355] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3354] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3353] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3352] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3351] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3350] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3349] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3348] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3347] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3346] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3345] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3344] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3343] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3342] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3341] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3340] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3339] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3338] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3337] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3336] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3335] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3334] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3333] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3332] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3331] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3330] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3329] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3328] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3327] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3326] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3325] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3324] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3323] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3322] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3321] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3320] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3319] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3318] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3317] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3316] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3315] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3314] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3313] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3312] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3311] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3310] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3309] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3308] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3307] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3306] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3305] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3304] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3303] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3302] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3301] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3300] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3299] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3298] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3297] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3296] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3295] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3294] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3293] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3292] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3291] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3290] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3289] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3288] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3287] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3286] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N447) begin
      mem[3285] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3284] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3283] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3282] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3281] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3280] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3279] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3278] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3277] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3276] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3275] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3274] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3273] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3272] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3271] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3270] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3269] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3268] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3267] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3266] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3265] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3264] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3263] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3262] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3261] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3260] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3259] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3258] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3257] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3256] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3255] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3254] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3253] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3252] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3251] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3250] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3249] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3248] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3247] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3246] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3245] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3244] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3243] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3242] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3241] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3240] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3239] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3238] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3237] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3236] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3235] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3234] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3233] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3232] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3231] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3230] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3229] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3228] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3227] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3226] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3225] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3224] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3223] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3222] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3221] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3220] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3219] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3218] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3217] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3216] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3215] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3214] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3213] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N446) begin
      mem[3212] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3211] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3210] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3209] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3208] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3207] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3206] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3205] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3204] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3203] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3202] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3201] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3200] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3199] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3198] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3197] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3196] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3195] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3194] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3193] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3192] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3191] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3190] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3189] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3188] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3187] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3186] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3185] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3184] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3183] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3182] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3181] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3180] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3179] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3178] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3177] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3176] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3175] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3174] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3173] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3172] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3171] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3170] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3169] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3168] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3167] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3166] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3165] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3164] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3163] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3162] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3161] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3160] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3159] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3158] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3157] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3156] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3155] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3154] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3153] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3152] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3151] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3150] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3149] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3148] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3147] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3146] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3145] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3144] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3143] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3142] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3141] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3140] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N445) begin
      mem[3139] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3138] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3137] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3136] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3135] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3134] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3133] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3132] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3131] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3130] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3129] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3128] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3127] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3126] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3125] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3124] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3123] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3122] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3121] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3120] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3119] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3118] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3117] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3116] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3115] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3114] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3113] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3112] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3111] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3110] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3109] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3108] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3107] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3106] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3105] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3104] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3103] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3102] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3101] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3100] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3099] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3098] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3097] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3096] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3095] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3094] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3093] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3092] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3091] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3090] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3089] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3088] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3087] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3086] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3085] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3084] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3083] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3082] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3081] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3080] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3079] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3078] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3077] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3076] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3075] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3074] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3073] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3072] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3071] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3070] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3069] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3068] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3067] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N444) begin
      mem[3066] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3065] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3064] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3063] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3062] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3061] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3060] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3059] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3058] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3057] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3056] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3055] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3054] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3053] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3052] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3051] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3050] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3049] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3048] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3047] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3046] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3045] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3044] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3043] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3042] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3041] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3040] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3039] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3038] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3037] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3036] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3035] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3034] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3033] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3032] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3031] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3030] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3029] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3028] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3027] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3026] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3025] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3024] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3023] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3022] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3021] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3020] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3019] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3018] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3017] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3016] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3015] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3014] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3013] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3012] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3011] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3010] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3009] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3008] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3007] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3006] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3005] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3004] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3003] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3002] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3001] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[3000] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[2999] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[2998] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[2997] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[2996] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[2995] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[2994] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N443) begin
      mem[2993] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2992] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2991] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2990] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2989] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2988] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2987] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2986] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2985] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2984] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2983] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2982] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2981] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2980] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2979] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2978] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2977] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2976] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2975] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2974] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2973] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2972] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2971] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2970] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2969] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2968] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2967] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2966] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2965] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2964] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2963] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2962] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2961] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2960] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2959] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2958] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2957] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2956] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2955] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2954] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2953] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2952] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2951] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2950] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2949] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2948] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2947] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2946] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2945] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2944] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2943] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2942] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2941] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2940] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2939] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2938] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2937] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2936] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2935] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2934] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2933] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2932] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2931] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2930] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2929] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2928] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2927] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2926] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2925] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2924] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2923] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2922] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2921] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N442) begin
      mem[2920] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2919] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2918] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2917] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2916] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2915] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2914] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2913] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2912] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2911] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2910] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2909] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2908] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2907] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2906] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2905] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2904] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2903] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2902] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2901] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2900] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2899] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2898] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2897] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2896] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2895] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2894] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2893] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2892] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2891] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2890] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2889] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2888] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2887] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2886] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2885] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2884] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2883] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2882] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2881] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2880] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2879] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2878] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2877] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2876] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2875] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2874] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2873] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2872] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2871] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2870] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2869] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2868] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2867] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2866] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2865] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2864] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2863] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2862] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2861] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2860] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2859] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2858] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2857] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2856] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2855] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2854] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2853] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2852] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2851] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2850] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2849] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2848] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N441) begin
      mem[2847] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2846] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2845] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2844] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2843] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2842] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2841] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2840] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2839] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2838] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2837] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2836] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2835] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2834] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2833] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2832] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2831] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2830] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2829] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2828] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2827] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2826] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2825] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2824] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2823] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2822] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2821] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2820] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2819] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2818] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2817] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2816] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2815] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2814] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2813] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2812] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2811] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2810] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2809] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2808] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2807] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2806] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2805] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2804] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2803] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2802] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2801] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2800] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2799] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2798] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2797] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2796] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2795] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2794] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2793] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2792] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2791] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2790] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2789] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2788] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2787] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2786] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2785] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2784] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2783] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2782] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2781] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2780] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2779] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2778] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2777] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2776] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2775] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N440) begin
      mem[2774] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2773] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2772] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2771] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2770] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2769] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2768] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2767] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2766] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2765] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2764] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2763] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2762] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2761] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2760] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2759] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2758] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2757] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2756] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2755] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2754] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2753] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2752] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2751] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2750] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2749] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2748] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2747] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2746] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2745] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2744] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2743] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2742] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2741] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2740] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2739] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2738] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2737] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2736] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2735] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2734] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2733] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2732] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2731] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2730] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2729] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2728] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2727] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2726] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2725] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2724] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2723] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2722] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2721] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2720] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2719] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2718] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2717] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2716] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2715] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2714] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2713] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2712] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2711] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2710] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2709] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2708] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2707] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2706] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2705] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2704] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2703] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2702] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N439) begin
      mem[2701] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2700] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2699] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2698] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2697] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2696] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2695] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2694] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2693] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2692] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2691] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2690] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2689] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2688] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2687] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2686] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2685] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2684] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2683] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2682] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2681] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2680] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2679] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2678] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2677] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2676] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2675] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2674] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2673] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2672] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2671] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2670] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2669] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2668] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2667] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2666] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2665] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2664] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2663] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2662] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2661] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2660] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2659] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2658] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2657] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2656] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2655] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2654] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2653] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2652] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2651] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2650] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2649] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2648] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2647] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2646] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2645] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2644] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2643] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2642] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2641] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2640] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2639] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2638] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2637] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2636] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2635] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2634] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2633] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2632] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2631] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2630] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2629] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N438) begin
      mem[2628] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2627] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2626] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2625] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2624] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2623] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2622] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2621] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2620] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2619] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2618] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2617] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2616] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2615] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2614] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2613] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2612] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2611] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2610] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2609] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2608] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2607] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2606] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2605] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2604] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2603] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2602] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2601] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2600] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2599] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2598] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2597] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2596] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2595] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2594] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2593] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2592] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2591] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2590] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2589] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2588] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2587] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2586] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2585] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2584] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2583] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2582] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2581] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2580] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2579] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2578] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2577] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2576] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2575] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2574] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2573] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2572] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2571] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2570] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2569] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2568] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2567] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2566] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2565] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2564] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2563] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2562] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2561] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2560] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2559] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2558] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2557] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2556] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N437) begin
      mem[2555] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2554] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2553] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2552] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2551] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2550] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2549] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2548] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2547] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2546] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2545] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2544] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2543] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2542] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2541] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2540] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2539] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2538] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2537] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2536] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2535] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2534] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2533] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2532] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2531] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2530] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2529] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2528] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2527] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2526] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2525] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2524] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2523] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2522] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2521] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2520] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2519] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2518] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2517] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2516] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2515] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2514] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2513] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2512] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2511] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2510] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2509] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2508] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2507] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2506] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2505] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2504] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2503] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2502] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2501] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2500] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2499] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2498] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2497] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2496] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2495] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2494] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2493] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2492] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2491] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2490] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2489] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2488] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2487] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2486] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2485] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2484] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2483] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N436) begin
      mem[2482] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2481] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2480] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2479] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2478] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2477] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2476] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2475] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2474] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2473] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2472] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2471] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2470] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2469] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2468] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2467] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2466] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2465] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2464] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2463] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2462] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2461] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2460] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2459] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2458] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2457] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2456] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2455] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2454] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2453] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2452] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2451] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2450] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2449] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2448] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2447] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2446] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2445] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2444] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2443] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2442] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2441] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2440] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2439] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2438] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2437] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2436] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2435] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2434] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2433] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2432] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2431] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2430] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2429] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2428] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2427] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2426] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2425] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2424] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2423] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2422] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2421] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2420] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2419] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2418] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2417] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2416] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2415] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2414] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2413] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2412] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2411] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2410] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N435) begin
      mem[2409] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2408] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2407] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2406] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2405] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2404] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2403] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2402] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2401] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2400] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2399] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2398] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2397] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2396] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2395] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2394] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2393] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2392] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2391] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2390] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2389] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2388] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2387] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2386] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2385] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2384] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2383] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2382] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2381] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2380] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2379] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2378] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2377] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2376] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2375] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2374] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2373] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2372] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2371] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2370] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2369] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2368] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2367] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2366] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2365] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2364] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2363] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2362] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2361] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2360] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2359] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2358] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2357] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2356] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2355] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2354] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2353] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2352] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2351] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2350] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2349] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2348] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2347] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2346] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2345] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2344] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2343] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2342] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2341] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2340] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2339] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2338] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2337] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N434) begin
      mem[2336] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2335] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2334] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2333] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2332] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2331] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2330] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2329] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2328] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2327] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2326] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2325] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2324] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2323] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2322] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2321] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2320] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2319] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2318] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2317] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2316] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2315] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2314] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2313] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2312] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2311] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2310] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2309] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2308] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2307] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2306] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2305] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2304] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2303] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2302] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2301] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2300] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2299] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2298] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2297] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2296] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2295] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2294] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2293] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2292] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2291] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2290] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2289] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2288] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2287] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2286] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2285] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2284] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2283] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2282] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2281] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2280] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2279] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2278] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2277] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2276] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2275] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2274] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2273] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2272] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2271] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2270] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2269] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2268] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2267] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2266] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2265] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2264] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N433) begin
      mem[2263] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2262] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2261] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2260] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2259] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2258] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2257] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2256] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2255] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2254] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2253] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2252] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2251] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2250] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2249] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2248] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2247] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2246] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2245] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2244] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2243] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2242] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2241] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2240] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2239] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2238] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2237] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2236] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2235] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2234] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2233] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2232] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2231] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2230] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2229] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2228] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2227] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2226] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2225] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2224] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2223] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2222] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2221] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2220] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2219] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2218] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2217] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2216] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2215] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2214] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2213] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2212] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2211] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2210] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2209] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2208] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2207] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2206] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2205] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2204] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2203] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2202] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2201] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2200] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2199] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2198] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2197] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2196] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2195] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2194] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2193] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2192] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2191] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N432) begin
      mem[2190] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2189] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2188] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2187] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2186] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2185] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2184] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2183] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2182] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2181] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2180] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2179] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2178] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2177] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2176] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2175] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2174] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2173] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2172] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2171] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2170] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2169] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2168] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2167] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2166] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2165] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2164] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2163] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2162] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2161] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2160] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2159] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2158] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2157] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2156] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2155] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2154] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2153] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2152] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2151] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2150] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2149] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2148] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2147] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2146] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2145] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2144] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2143] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2142] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2141] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2140] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2139] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2138] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2137] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2136] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2135] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2134] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2133] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2132] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2131] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2130] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2129] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2128] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2127] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2126] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2125] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2124] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2123] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2122] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2121] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2120] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2119] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2118] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N431) begin
      mem[2117] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2116] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2115] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2114] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2113] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2112] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2111] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2110] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2109] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2108] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2107] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2106] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2105] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2104] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2103] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2102] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2101] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2100] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2099] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2098] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2097] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2096] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2095] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2094] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2093] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2092] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2091] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2090] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2089] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2088] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2087] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2086] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2085] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2084] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2083] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2082] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2081] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2080] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2079] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2078] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2077] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2076] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2075] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2074] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2073] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2072] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2071] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2070] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2069] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2068] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2067] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2066] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2065] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2064] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2063] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2062] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2061] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2060] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2059] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2058] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2057] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2056] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2055] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2054] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2053] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2052] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2051] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2050] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2049] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2048] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2047] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2046] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2045] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N430) begin
      mem[2044] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2043] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2042] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2041] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2040] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2039] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2038] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2037] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2036] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2035] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2034] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2033] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2032] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2031] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2030] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2029] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2028] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2027] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2026] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2025] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2024] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2023] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2022] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2021] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2020] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2019] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2018] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2017] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2016] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2015] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2014] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2013] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2012] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2011] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2010] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2009] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2008] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2007] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2006] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2005] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2004] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2003] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2002] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2001] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[2000] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1999] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1998] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1997] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1996] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1995] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1994] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1993] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1992] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1991] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1990] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1989] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1988] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1987] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1986] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1985] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1984] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1983] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1982] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1981] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1980] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1979] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1978] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1977] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1976] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1975] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1974] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1973] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1972] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N429) begin
      mem[1971] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1970] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1969] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1968] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1967] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1966] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1965] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1964] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1963] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1962] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1961] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1960] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1959] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1958] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1957] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1956] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1955] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1954] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1953] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1952] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1951] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1950] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1949] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1948] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1947] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1946] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1945] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1944] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1943] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1942] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1941] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1940] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1939] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1938] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1937] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1936] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1935] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1934] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1933] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1932] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1931] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1930] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1929] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1928] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1927] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1926] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1925] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1924] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1923] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1922] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1921] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1920] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1919] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1918] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1917] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1916] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1915] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1914] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1913] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1912] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1911] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1910] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1909] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1908] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1907] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1906] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1905] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1904] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1903] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1902] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1901] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1900] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1899] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N428) begin
      mem[1898] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1897] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1896] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1895] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1894] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1893] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1892] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1891] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1890] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1889] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1888] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1887] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1886] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1885] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1884] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1883] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1882] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1881] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1880] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1879] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1878] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1877] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1876] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1875] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1874] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1873] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1872] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1871] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1870] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1869] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1868] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1867] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1866] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1865] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1864] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1863] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1862] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1861] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1860] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1859] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1858] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1857] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1856] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1855] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1854] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1853] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1852] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1851] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1850] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1849] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1848] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1847] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1846] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1845] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1844] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1843] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1842] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1841] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1840] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1839] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1838] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1837] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1836] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1835] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1834] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1833] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1832] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1831] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1830] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1829] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1828] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1827] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1826] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N427) begin
      mem[1825] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1824] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1823] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1822] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1821] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1820] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1819] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1818] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1817] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1816] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1815] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1814] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1813] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1812] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1811] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1810] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1809] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1808] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1807] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1806] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1805] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1804] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1803] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1802] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1801] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1800] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1799] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1798] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1797] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1796] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1795] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1794] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1793] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1792] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1791] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1790] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1789] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1788] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1787] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1786] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1785] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1784] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1783] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1782] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1781] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1780] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1779] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1778] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1777] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1776] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1775] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1774] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1773] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1772] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1771] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1770] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1769] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1768] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1767] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1766] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1765] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1764] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1763] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1762] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1761] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1760] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1759] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1758] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1757] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1756] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1755] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1754] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1753] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N426) begin
      mem[1752] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1751] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1750] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1749] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1748] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1747] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1746] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1745] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1744] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1743] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1742] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1741] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1740] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1739] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1738] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1737] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1736] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1735] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1734] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1733] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1732] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1731] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1730] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1729] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1728] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1727] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1726] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1725] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1724] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1723] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1722] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1721] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1720] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1719] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1718] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1717] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1716] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1715] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1714] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1713] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1712] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1711] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1710] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1709] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1708] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1707] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1706] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1705] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1704] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1703] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1702] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1701] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1700] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1699] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1698] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1697] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1696] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1695] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1694] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1693] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1692] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1691] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1690] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1689] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1688] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1687] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1686] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1685] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1684] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1683] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1682] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1681] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1680] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N425) begin
      mem[1679] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1678] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1677] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1676] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1675] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1674] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1673] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1672] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1671] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1670] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1669] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1668] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1667] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1666] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1665] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1664] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1663] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1662] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1661] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1660] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1659] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1658] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1657] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1656] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1655] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1654] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1653] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1652] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1651] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1650] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1649] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1648] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1647] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1646] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1645] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1644] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1643] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1642] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1641] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1640] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1639] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1638] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1637] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1636] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1635] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1634] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1633] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1632] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1631] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1630] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1629] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1628] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1627] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1626] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1625] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1624] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1623] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1622] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1621] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1620] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1619] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1618] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1617] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1616] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1615] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1614] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1613] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1612] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1611] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1610] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1609] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1608] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1607] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N424) begin
      mem[1606] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1605] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1604] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1603] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1602] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1601] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1600] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1599] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1598] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1597] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1596] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1595] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1594] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1593] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1592] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1591] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1590] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1589] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1588] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1587] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1586] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1585] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1584] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1583] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1582] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1581] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1580] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1579] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1578] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1577] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1576] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1575] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1574] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1573] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1572] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1571] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1570] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1569] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1568] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1567] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1566] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1565] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1564] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1563] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1562] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1561] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1560] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1559] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1558] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1557] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1556] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1555] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1554] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1553] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1552] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1551] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1550] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1549] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1548] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1547] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1546] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1545] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1544] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1543] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1542] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1541] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1540] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1539] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1538] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1537] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1536] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1535] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1534] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N423) begin
      mem[1533] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1532] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1531] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1530] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1529] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1528] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1527] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1526] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1525] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1524] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1523] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1522] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1521] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1520] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1519] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1518] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1517] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1516] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1515] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1514] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1513] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1512] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1511] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1510] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1509] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1508] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1507] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1506] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1505] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1504] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1503] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1502] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1501] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1500] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1499] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1498] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1497] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1496] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1495] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1494] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1493] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1492] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1491] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1490] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1489] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1488] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1487] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1486] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1485] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1484] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1483] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1482] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1481] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1480] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1479] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1478] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1477] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1476] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1475] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1474] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1473] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1472] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1471] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1470] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1469] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1468] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1467] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1466] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1465] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1464] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1463] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1462] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1461] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N422) begin
      mem[1460] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1459] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1458] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1457] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1456] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1455] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1454] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1453] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1452] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1451] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1450] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1449] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1448] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1447] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1446] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1445] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1444] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1443] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1442] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1441] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1440] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1439] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1438] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1437] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1436] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1435] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1434] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1433] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1432] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1431] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1430] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1429] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1428] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1427] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1426] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1425] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1424] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1423] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1422] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1421] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1420] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1419] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1418] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1417] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1416] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1415] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1414] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1413] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1412] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1411] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1410] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1409] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1408] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1407] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1406] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1405] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1404] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1403] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1402] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1401] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1400] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1399] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1398] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1397] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1396] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1395] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1394] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1393] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1392] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1391] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1390] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1389] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1388] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N421) begin
      mem[1387] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1386] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1385] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1384] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1383] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1382] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1381] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1380] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1379] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1378] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1377] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1376] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1375] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1374] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1373] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1372] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1371] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1370] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1369] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1368] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1367] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1366] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1365] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1364] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1363] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1362] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1361] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1360] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1359] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1358] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1357] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1356] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1355] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1354] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1353] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1352] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1351] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1350] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1349] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1348] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1347] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1346] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1345] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1344] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1343] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1342] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1341] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1340] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1339] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1338] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1337] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1336] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1335] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1334] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1333] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1332] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1331] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1330] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1329] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1328] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1327] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1326] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1325] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1324] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1323] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1322] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1321] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1320] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1319] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1318] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1317] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1316] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1315] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N420) begin
      mem[1314] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1313] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1312] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1311] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1310] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1309] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1308] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1307] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1306] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1305] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1304] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1303] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1302] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1301] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1300] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1299] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1298] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1297] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1296] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1295] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1294] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1293] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1292] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1291] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1290] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1289] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1288] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1287] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1286] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1285] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1284] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1283] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1282] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1281] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1280] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1279] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1278] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1277] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1276] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1275] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1274] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1273] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1272] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1271] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1270] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1269] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1268] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1267] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1266] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1265] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1264] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1263] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1262] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1261] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1260] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1259] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1258] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1257] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1256] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1255] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1254] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1253] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1252] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1251] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1250] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1249] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1248] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1247] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1246] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1245] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1244] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1243] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1242] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N419) begin
      mem[1241] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1240] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1239] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1238] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1237] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1236] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1235] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1234] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1233] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1232] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1231] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1230] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1229] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1228] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1227] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1226] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1225] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1224] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1223] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1222] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1221] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1220] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1219] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1218] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1217] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1216] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1215] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1214] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1213] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1212] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1211] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1210] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1209] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1208] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1207] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1206] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1205] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1204] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1203] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1202] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1201] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1200] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1199] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1198] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1197] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1196] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1195] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1194] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1193] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1192] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1191] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1190] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1189] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1188] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1187] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1186] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1185] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1184] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1183] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1182] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1181] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1180] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1179] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1178] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1177] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1176] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1175] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1174] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1173] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1172] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1171] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1170] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1169] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N418) begin
      mem[1168] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1167] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1166] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1165] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1164] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1163] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1162] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1161] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1160] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1159] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1158] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1157] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1156] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1155] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1154] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1153] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1152] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1151] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1150] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1149] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1148] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1147] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1146] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1145] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1144] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1143] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1142] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1141] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1140] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1139] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1138] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1137] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1136] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1135] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1134] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1133] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1132] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1131] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1130] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1129] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1128] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1127] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1126] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1125] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1124] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1123] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1122] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1121] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1120] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1119] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1118] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1117] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1116] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1115] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1114] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1113] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1112] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1111] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1110] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1109] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1108] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1107] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1106] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1105] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1104] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1103] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1102] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1101] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1100] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1099] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1098] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1097] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1096] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N417) begin
      mem[1095] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1094] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1093] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1092] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1091] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1090] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1089] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1088] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1087] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1086] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1085] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1084] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1083] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1082] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1081] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1080] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1079] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1078] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1077] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1076] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1075] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1074] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1073] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1072] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1071] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1070] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1069] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1068] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1067] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1066] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1065] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1064] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1063] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1062] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1061] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1060] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1059] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1058] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1057] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1056] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1055] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1054] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1053] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1052] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1051] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1050] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1049] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1048] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1047] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1046] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1045] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1044] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1043] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1042] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1041] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1040] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1039] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1038] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1037] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1036] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1035] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1034] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1033] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1032] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1031] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1030] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1029] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1028] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1027] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1026] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1025] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1024] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1023] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N416) begin
      mem[1022] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1021] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1020] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1019] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1018] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1017] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1016] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1015] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1014] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1013] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1012] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1011] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1010] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1009] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1008] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1007] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1006] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1005] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1004] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1003] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1002] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1001] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[1000] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[999] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[998] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[997] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[996] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[995] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[994] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[993] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[992] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[991] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[990] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[989] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[988] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[987] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[986] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[985] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[984] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[983] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[982] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[981] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[980] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[979] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[978] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[977] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[976] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[975] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[974] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[973] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[972] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[971] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[970] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[969] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[968] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[967] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[966] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[965] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[964] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[963] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[962] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[961] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[960] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[959] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[958] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[957] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[956] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[955] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[954] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[953] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[952] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[951] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[950] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N415) begin
      mem[949] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[948] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[947] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[946] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[945] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[944] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[943] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[942] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[941] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[940] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[939] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[938] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[937] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[936] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[935] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[934] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[933] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[932] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[931] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[930] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[929] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[928] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[927] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[926] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[925] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[924] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[923] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[922] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[921] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[920] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[919] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[918] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[917] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[916] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[915] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[914] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[913] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[912] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[911] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[910] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[909] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[908] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[907] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[906] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[905] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[904] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[903] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[902] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[901] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[900] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[899] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[898] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[897] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[896] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[895] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[894] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[893] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[892] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[891] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[890] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[889] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[888] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[887] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[886] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[885] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[884] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[883] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[882] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[881] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[880] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[879] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[878] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[877] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N414) begin
      mem[876] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[875] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[874] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[873] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[872] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[871] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[870] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[869] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[868] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[867] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[866] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[865] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[864] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[863] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[862] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[861] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[860] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[859] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[858] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[857] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[856] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[855] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[854] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[853] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[852] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[851] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[850] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[849] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[848] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[847] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[846] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[845] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[844] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[843] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[842] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[841] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[840] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[839] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[838] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[837] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[836] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[835] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[834] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[833] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[832] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[831] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[830] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[829] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[828] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[827] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[826] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[825] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[824] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[823] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[822] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[821] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[820] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[819] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[818] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[817] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[816] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[815] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[814] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[813] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[812] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[811] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[810] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[809] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[808] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[807] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[806] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[805] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[804] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N413) begin
      mem[803] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[802] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[801] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[800] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[799] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[798] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[797] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[796] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[795] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[794] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[793] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[792] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[791] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[790] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[789] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[788] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[787] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[786] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[785] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[784] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[783] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[782] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[781] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[780] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[779] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[778] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[777] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[776] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[775] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[774] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[773] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[772] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[771] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[770] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[769] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[768] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[767] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[766] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[765] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[764] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[763] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[762] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[761] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[760] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[759] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[758] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[757] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[756] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[755] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[754] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[753] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[752] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[751] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[750] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[749] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[748] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[747] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[746] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[745] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[744] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[743] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[742] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[741] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[740] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[739] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[738] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[737] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[736] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[735] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[734] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[733] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[732] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[731] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N412) begin
      mem[730] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[729] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[728] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[727] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[726] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[725] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[724] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[723] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[722] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[721] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[720] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[719] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[718] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[717] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[716] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[715] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[714] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[713] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[712] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[711] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[710] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[709] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[708] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[707] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[706] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[705] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[704] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[703] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[702] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[701] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[700] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[699] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[698] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[697] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[696] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[695] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[694] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[693] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[692] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[691] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[690] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[689] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[688] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[687] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[686] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[685] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[684] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[683] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[682] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[681] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[680] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[679] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[678] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[677] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[676] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[675] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[674] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[673] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[672] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[671] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[670] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[669] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[668] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[667] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[666] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[665] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[664] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[663] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[662] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[661] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[660] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[659] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[658] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N411) begin
      mem[657] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[656] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[655] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[654] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[653] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[652] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[651] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[650] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[649] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[648] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[647] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[646] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[645] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[644] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[643] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[642] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[641] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[640] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[639] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[638] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[637] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[636] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[635] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[634] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[633] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[632] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[631] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[630] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[629] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[628] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[627] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[626] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[625] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[624] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[623] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[622] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[621] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[620] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[619] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[618] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[617] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[616] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[615] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[614] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[613] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[612] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[611] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[610] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[609] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[608] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[607] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[606] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[605] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[604] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[603] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[602] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[601] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[600] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[599] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[598] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[597] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[596] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[595] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[594] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[593] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[592] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[591] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[590] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[589] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[588] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[587] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[586] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[585] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N410) begin
      mem[584] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[583] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[582] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[581] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[580] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[579] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[578] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[577] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[576] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[575] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[574] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[573] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[572] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[571] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[570] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[569] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[568] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[567] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[566] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[565] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[564] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[563] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[562] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[561] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[560] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[559] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[558] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[557] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[556] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[555] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[554] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[553] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[552] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[551] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[550] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[549] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[548] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[547] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[546] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[545] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[544] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[543] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[542] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[541] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[540] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[539] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[538] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[537] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[536] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[535] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[534] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[533] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[532] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[531] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[530] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[529] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[528] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[527] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[526] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[525] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[524] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[523] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[522] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[521] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[520] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[519] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[518] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[517] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[516] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[515] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[514] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[513] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[512] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N409) begin
      mem[511] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[510] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[509] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[508] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[507] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[506] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[505] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[504] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[503] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[502] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[501] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[500] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[499] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[498] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[497] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[496] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[495] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[494] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[493] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[492] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[491] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[490] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[489] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[488] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[487] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[486] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[485] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[484] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[483] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[482] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[481] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[480] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[479] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[478] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[477] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[476] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[475] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[474] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[473] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[472] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[471] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[470] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[469] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[468] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[467] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[466] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[465] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[464] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[463] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[462] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[461] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[460] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[459] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[458] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[457] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[456] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[455] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[454] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[453] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[452] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[451] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[450] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[449] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[448] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[447] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[446] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[445] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[444] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[443] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[442] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[441] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[440] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[439] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N408) begin
      mem[438] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[437] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[436] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[435] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[434] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[433] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[432] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[431] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[430] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[429] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[428] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[427] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[426] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[425] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[424] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[423] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[422] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[421] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[420] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[419] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[418] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[417] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[416] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[415] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[414] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[413] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[412] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[411] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[410] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[409] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[408] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[407] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[406] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[405] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[404] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[403] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[402] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[401] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[400] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[399] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[398] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[397] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[396] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[395] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[394] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[393] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[392] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[391] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[390] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[389] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[388] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[387] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[386] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[385] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[384] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[383] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[382] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[381] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[380] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[379] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[378] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[377] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[376] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[375] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[374] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[373] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[372] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[371] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[370] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[369] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[368] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[367] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[366] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N407) begin
      mem[365] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[364] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[363] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[362] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[361] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[360] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[359] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[358] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[357] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[356] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[355] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[354] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[353] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[352] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[351] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[350] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[349] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[348] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[347] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[346] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[345] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[344] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[343] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[342] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[341] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[340] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[339] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[338] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[337] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[336] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[335] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[334] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[333] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[332] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[331] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[330] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[329] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[328] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[327] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[326] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[325] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[324] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[323] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[322] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[321] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[320] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[319] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[318] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[317] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[316] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[315] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[314] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[313] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[312] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[311] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[310] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[309] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[308] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[307] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[306] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[305] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[304] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[303] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[302] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[301] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[300] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[299] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[298] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[297] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[296] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[295] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[294] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[293] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N406) begin
      mem[292] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[291] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[290] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[289] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[288] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[287] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[286] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[285] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[284] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[283] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[282] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[281] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[280] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[279] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[278] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[277] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[276] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[275] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[274] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[273] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[272] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[271] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[270] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[269] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[268] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[267] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[266] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[265] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[264] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[263] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[262] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[261] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[260] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[259] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[258] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[257] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[256] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[255] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[254] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[253] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[252] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[251] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[250] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[249] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[248] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[247] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[246] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[245] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[244] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[243] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[242] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[241] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[240] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[239] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[238] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[237] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[236] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[235] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[234] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[233] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[232] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[231] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[230] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[229] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[228] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[227] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[226] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[225] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[224] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[223] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[222] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[221] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[220] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N405) begin
      mem[219] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[218] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[217] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[216] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[215] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[214] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[213] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[212] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[211] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[210] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[209] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[208] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[207] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[206] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[205] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[204] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[203] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[202] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[201] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[200] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[199] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[198] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[197] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[196] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[195] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[194] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[193] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[192] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[191] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[190] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[189] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[188] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[187] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[186] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[185] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[184] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[183] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[182] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[181] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[180] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[179] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[178] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[177] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[176] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[175] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[174] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[173] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[172] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[171] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[170] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[169] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[168] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[167] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[166] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[165] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[164] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[163] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[162] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[161] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[160] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[159] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[158] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[157] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[156] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[155] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[154] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[153] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[152] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[151] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[150] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[149] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[148] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[147] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N404) begin
      mem[146] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[145] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[144] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[143] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[142] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[141] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[140] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[139] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[138] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[137] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[136] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[135] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[134] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[133] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[132] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[131] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[130] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[129] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[128] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[127] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[126] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[125] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[124] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[123] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[122] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[121] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[120] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[119] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[118] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[117] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[116] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[115] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[114] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[113] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[112] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[111] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[110] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[109] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[108] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[107] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[106] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[105] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[104] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[103] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[102] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[101] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[100] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[99] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[98] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[97] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[96] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[95] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[94] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[93] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[92] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[91] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[90] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[89] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[88] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[87] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[86] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[85] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[84] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[83] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[82] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[81] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[80] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[79] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[78] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[77] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[76] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[75] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[74] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N403) begin
      mem[73] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[72] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[71] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[70] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[69] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[68] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[67] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[66] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[65] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[64] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[63] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[62] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[61] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[60] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[59] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[58] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[57] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[56] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[55] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[54] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[53] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[52] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[51] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[50] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[49] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[48] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[47] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[46] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[45] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[44] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[43] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[42] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[41] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[40] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[39] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[38] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[37] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[36] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[35] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[34] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[33] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[32] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[31] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[30] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[29] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[28] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[27] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[26] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[25] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[24] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[23] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[22] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[21] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[20] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[19] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[18] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[17] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[16] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[15] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[14] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[13] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[12] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[11] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[10] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[9] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[8] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[7] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[6] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[5] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[4] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[3] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[2] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[1] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N402) begin
      mem[0] <= w_data_i[0];
    end 
  end

  assign N530 = ~w_addr_i[6];
  assign N531 = w_addr_i[4] & w_addr_i[5];
  assign N532 = N0 & w_addr_i[5];
  assign N0 = ~w_addr_i[4];
  assign N533 = w_addr_i[4] & N1;
  assign N1 = ~w_addr_i[5];
  assign N534 = N2 & N3;
  assign N2 = ~w_addr_i[4];
  assign N3 = ~w_addr_i[5];
  assign N535 = w_addr_i[6] & N531;
  assign N536 = w_addr_i[6] & N532;
  assign N537 = w_addr_i[6] & N533;
  assign N538 = w_addr_i[6] & N534;
  assign N539 = N530 & N531;
  assign N540 = N530 & N532;
  assign N541 = N530 & N533;
  assign N542 = N530 & N534;
  assign N543 = w_addr_i[2] & w_addr_i[3];
  assign N544 = N4 & w_addr_i[3];
  assign N4 = ~w_addr_i[2];
  assign N545 = w_addr_i[2] & N5;
  assign N5 = ~w_addr_i[3];
  assign N546 = N6 & N7;
  assign N6 = ~w_addr_i[2];
  assign N7 = ~w_addr_i[3];
  assign N547 = w_addr_i[0] & w_addr_i[1];
  assign N548 = N8 & w_addr_i[1];
  assign N8 = ~w_addr_i[0];
  assign N549 = w_addr_i[0] & N9;
  assign N9 = ~w_addr_i[1];
  assign N550 = N10 & N11;
  assign N10 = ~w_addr_i[0];
  assign N11 = ~w_addr_i[1];
  assign N551 = N543 & N547;
  assign N552 = N543 & N548;
  assign N553 = N543 & N549;
  assign N554 = N543 & N550;
  assign N555 = N544 & N547;
  assign N556 = N544 & N548;
  assign N557 = N544 & N549;
  assign N558 = N544 & N550;
  assign N559 = N545 & N547;
  assign N560 = N545 & N548;
  assign N561 = N545 & N549;
  assign N562 = N545 & N550;
  assign N563 = N546 & N547;
  assign N564 = N546 & N548;
  assign N565 = N546 & N549;
  assign N566 = N546 & N550;
  assign N401 = N535 & N551;
  assign N400 = N535 & N552;
  assign N399 = N535 & N553;
  assign N398 = N535 & N554;
  assign N397 = N535 & N555;
  assign N396 = N535 & N556;
  assign N395 = N535 & N557;
  assign N394 = N535 & N558;
  assign N393 = N535 & N559;
  assign N392 = N535 & N560;
  assign N391 = N535 & N561;
  assign N390 = N535 & N562;
  assign N389 = N535 & N563;
  assign N388 = N535 & N564;
  assign N387 = N535 & N565;
  assign N386 = N535 & N566;
  assign N385 = N536 & N551;
  assign N384 = N536 & N552;
  assign N383 = N536 & N553;
  assign N382 = N536 & N554;
  assign N381 = N536 & N555;
  assign N380 = N536 & N556;
  assign N379 = N536 & N557;
  assign N378 = N536 & N558;
  assign N377 = N536 & N559;
  assign N376 = N536 & N560;
  assign N375 = N536 & N561;
  assign N374 = N536 & N562;
  assign N373 = N536 & N563;
  assign N372 = N536 & N564;
  assign N371 = N536 & N565;
  assign N370 = N536 & N566;
  assign N369 = N537 & N551;
  assign N368 = N537 & N552;
  assign N367 = N537 & N553;
  assign N366 = N537 & N554;
  assign N365 = N537 & N555;
  assign N364 = N537 & N556;
  assign N363 = N537 & N557;
  assign N362 = N537 & N558;
  assign N361 = N537 & N559;
  assign N360 = N537 & N560;
  assign N359 = N537 & N561;
  assign N358 = N537 & N562;
  assign N357 = N537 & N563;
  assign N356 = N537 & N564;
  assign N355 = N537 & N565;
  assign N354 = N537 & N566;
  assign N353 = N538 & N551;
  assign N352 = N538 & N552;
  assign N351 = N538 & N553;
  assign N350 = N538 & N554;
  assign N349 = N538 & N555;
  assign N348 = N538 & N556;
  assign N347 = N538 & N557;
  assign N346 = N538 & N558;
  assign N345 = N538 & N559;
  assign N344 = N538 & N560;
  assign N343 = N538 & N561;
  assign N342 = N538 & N562;
  assign N341 = N538 & N563;
  assign N340 = N538 & N564;
  assign N339 = N538 & N565;
  assign N338 = N538 & N566;
  assign N337 = N539 & N551;
  assign N336 = N539 & N552;
  assign N335 = N539 & N553;
  assign N334 = N539 & N554;
  assign N333 = N539 & N555;
  assign N332 = N539 & N556;
  assign N331 = N539 & N557;
  assign N330 = N539 & N558;
  assign N329 = N539 & N559;
  assign N328 = N539 & N560;
  assign N327 = N539 & N561;
  assign N326 = N539 & N562;
  assign N325 = N539 & N563;
  assign N324 = N539 & N564;
  assign N323 = N539 & N565;
  assign N322 = N539 & N566;
  assign N321 = N540 & N551;
  assign N320 = N540 & N552;
  assign N319 = N540 & N553;
  assign N318 = N540 & N554;
  assign N317 = N540 & N555;
  assign N316 = N540 & N556;
  assign N315 = N540 & N557;
  assign N314 = N540 & N558;
  assign N313 = N540 & N559;
  assign N312 = N540 & N560;
  assign N311 = N540 & N561;
  assign N310 = N540 & N562;
  assign N309 = N540 & N563;
  assign N308 = N540 & N564;
  assign N307 = N540 & N565;
  assign N306 = N540 & N566;
  assign N305 = N541 & N551;
  assign N304 = N541 & N552;
  assign N303 = N541 & N553;
  assign N302 = N541 & N554;
  assign N301 = N541 & N555;
  assign N300 = N541 & N556;
  assign N299 = N541 & N557;
  assign N298 = N541 & N558;
  assign N297 = N541 & N559;
  assign N296 = N541 & N560;
  assign N295 = N541 & N561;
  assign N294 = N541 & N562;
  assign N293 = N541 & N563;
  assign N292 = N541 & N564;
  assign N291 = N541 & N565;
  assign N290 = N541 & N566;
  assign N289 = N542 & N551;
  assign N288 = N542 & N552;
  assign N287 = N542 & N553;
  assign N286 = N542 & N554;
  assign N285 = N542 & N555;
  assign N284 = N542 & N556;
  assign N283 = N542 & N557;
  assign N282 = N542 & N558;
  assign N281 = N542 & N559;
  assign N280 = N542 & N560;
  assign N279 = N542 & N561;
  assign N278 = N542 & N562;
  assign N277 = N542 & N563;
  assign N276 = N542 & N564;
  assign N275 = N542 & N565;
  assign N274 = N542 & N566;
  assign { N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402 } = (N12)? { N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_v_i;
  assign N13 = N273;
  assign N14 = ~r_addr_i[0];
  assign N15 = ~r_addr_i[1];
  assign N16 = N14 & N15;
  assign N17 = N14 & r_addr_i[1];
  assign N18 = r_addr_i[0] & N15;
  assign N19 = r_addr_i[0] & r_addr_i[1];
  assign N20 = ~r_addr_i[2];
  assign N21 = N16 & N20;
  assign N22 = N16 & r_addr_i[2];
  assign N23 = N18 & N20;
  assign N24 = N18 & r_addr_i[2];
  assign N25 = N17 & N20;
  assign N26 = N17 & r_addr_i[2];
  assign N27 = N19 & N20;
  assign N28 = N19 & r_addr_i[2];
  assign N29 = ~r_addr_i[3];
  assign N30 = N21 & N29;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N29;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N25 & N29;
  assign N35 = N25 & r_addr_i[3];
  assign N36 = N27 & N29;
  assign N37 = N27 & r_addr_i[3];
  assign N38 = N22 & N29;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N29;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = N26 & N29;
  assign N43 = N26 & r_addr_i[3];
  assign N44 = N28 & N29;
  assign N45 = N28 & r_addr_i[3];
  assign N46 = ~r_addr_i[4];
  assign N47 = N30 & N46;
  assign N48 = N30 & r_addr_i[4];
  assign N49 = N32 & N46;
  assign N50 = N32 & r_addr_i[4];
  assign N51 = N34 & N46;
  assign N52 = N34 & r_addr_i[4];
  assign N53 = N36 & N46;
  assign N54 = N36 & r_addr_i[4];
  assign N55 = N38 & N46;
  assign N56 = N38 & r_addr_i[4];
  assign N57 = N40 & N46;
  assign N58 = N40 & r_addr_i[4];
  assign N59 = N42 & N46;
  assign N60 = N42 & r_addr_i[4];
  assign N61 = N44 & N46;
  assign N62 = N44 & r_addr_i[4];
  assign N63 = N31 & N46;
  assign N64 = N31 & r_addr_i[4];
  assign N65 = N33 & N46;
  assign N66 = N33 & r_addr_i[4];
  assign N67 = N35 & N46;
  assign N68 = N35 & r_addr_i[4];
  assign N69 = N37 & N46;
  assign N70 = N37 & r_addr_i[4];
  assign N71 = N39 & N46;
  assign N72 = N39 & r_addr_i[4];
  assign N73 = N41 & N46;
  assign N74 = N41 & r_addr_i[4];
  assign N75 = N43 & N46;
  assign N76 = N43 & r_addr_i[4];
  assign N77 = N45 & N46;
  assign N78 = N45 & r_addr_i[4];
  assign N79 = ~r_addr_i[5];
  assign N80 = N47 & N79;
  assign N81 = N47 & r_addr_i[5];
  assign N82 = N49 & N79;
  assign N83 = N49 & r_addr_i[5];
  assign N84 = N51 & N79;
  assign N85 = N51 & r_addr_i[5];
  assign N86 = N53 & N79;
  assign N87 = N53 & r_addr_i[5];
  assign N88 = N55 & N79;
  assign N89 = N55 & r_addr_i[5];
  assign N90 = N57 & N79;
  assign N91 = N57 & r_addr_i[5];
  assign N92 = N59 & N79;
  assign N93 = N59 & r_addr_i[5];
  assign N94 = N61 & N79;
  assign N95 = N61 & r_addr_i[5];
  assign N96 = N63 & N79;
  assign N97 = N63 & r_addr_i[5];
  assign N98 = N65 & N79;
  assign N99 = N65 & r_addr_i[5];
  assign N100 = N67 & N79;
  assign N101 = N67 & r_addr_i[5];
  assign N102 = N69 & N79;
  assign N103 = N69 & r_addr_i[5];
  assign N104 = N71 & N79;
  assign N105 = N71 & r_addr_i[5];
  assign N106 = N73 & N79;
  assign N107 = N73 & r_addr_i[5];
  assign N108 = N75 & N79;
  assign N109 = N75 & r_addr_i[5];
  assign N110 = N77 & N79;
  assign N111 = N77 & r_addr_i[5];
  assign N112 = N48 & N79;
  assign N113 = N48 & r_addr_i[5];
  assign N114 = N50 & N79;
  assign N115 = N50 & r_addr_i[5];
  assign N116 = N52 & N79;
  assign N117 = N52 & r_addr_i[5];
  assign N118 = N54 & N79;
  assign N119 = N54 & r_addr_i[5];
  assign N120 = N56 & N79;
  assign N121 = N56 & r_addr_i[5];
  assign N122 = N58 & N79;
  assign N123 = N58 & r_addr_i[5];
  assign N124 = N60 & N79;
  assign N125 = N60 & r_addr_i[5];
  assign N126 = N62 & N79;
  assign N127 = N62 & r_addr_i[5];
  assign N128 = N64 & N79;
  assign N129 = N64 & r_addr_i[5];
  assign N130 = N66 & N79;
  assign N131 = N66 & r_addr_i[5];
  assign N132 = N68 & N79;
  assign N133 = N68 & r_addr_i[5];
  assign N134 = N70 & N79;
  assign N135 = N70 & r_addr_i[5];
  assign N136 = N72 & N79;
  assign N137 = N72 & r_addr_i[5];
  assign N138 = N74 & N79;
  assign N139 = N74 & r_addr_i[5];
  assign N140 = N76 & N79;
  assign N141 = N76 & r_addr_i[5];
  assign N142 = N78 & N79;
  assign N143 = N78 & r_addr_i[5];
  assign N144 = ~r_addr_i[6];
  assign N145 = N80 & N144;
  assign N146 = N80 & r_addr_i[6];
  assign N147 = N82 & N144;
  assign N148 = N82 & r_addr_i[6];
  assign N149 = N84 & N144;
  assign N150 = N84 & r_addr_i[6];
  assign N151 = N86 & N144;
  assign N152 = N86 & r_addr_i[6];
  assign N153 = N88 & N144;
  assign N154 = N88 & r_addr_i[6];
  assign N155 = N90 & N144;
  assign N156 = N90 & r_addr_i[6];
  assign N157 = N92 & N144;
  assign N158 = N92 & r_addr_i[6];
  assign N159 = N94 & N144;
  assign N160 = N94 & r_addr_i[6];
  assign N161 = N96 & N144;
  assign N162 = N96 & r_addr_i[6];
  assign N163 = N98 & N144;
  assign N164 = N98 & r_addr_i[6];
  assign N165 = N100 & N144;
  assign N166 = N100 & r_addr_i[6];
  assign N167 = N102 & N144;
  assign N168 = N102 & r_addr_i[6];
  assign N169 = N104 & N144;
  assign N170 = N104 & r_addr_i[6];
  assign N171 = N106 & N144;
  assign N172 = N106 & r_addr_i[6];
  assign N173 = N108 & N144;
  assign N174 = N108 & r_addr_i[6];
  assign N175 = N110 & N144;
  assign N176 = N110 & r_addr_i[6];
  assign N177 = N112 & N144;
  assign N178 = N112 & r_addr_i[6];
  assign N179 = N114 & N144;
  assign N180 = N114 & r_addr_i[6];
  assign N181 = N116 & N144;
  assign N182 = N116 & r_addr_i[6];
  assign N183 = N118 & N144;
  assign N184 = N118 & r_addr_i[6];
  assign N185 = N120 & N144;
  assign N186 = N120 & r_addr_i[6];
  assign N187 = N122 & N144;
  assign N188 = N122 & r_addr_i[6];
  assign N189 = N124 & N144;
  assign N190 = N124 & r_addr_i[6];
  assign N191 = N126 & N144;
  assign N192 = N126 & r_addr_i[6];
  assign N193 = N128 & N144;
  assign N194 = N128 & r_addr_i[6];
  assign N195 = N130 & N144;
  assign N196 = N130 & r_addr_i[6];
  assign N197 = N132 & N144;
  assign N198 = N132 & r_addr_i[6];
  assign N199 = N134 & N144;
  assign N200 = N134 & r_addr_i[6];
  assign N201 = N136 & N144;
  assign N202 = N136 & r_addr_i[6];
  assign N203 = N138 & N144;
  assign N204 = N138 & r_addr_i[6];
  assign N205 = N140 & N144;
  assign N206 = N140 & r_addr_i[6];
  assign N207 = N142 & N144;
  assign N208 = N142 & r_addr_i[6];
  assign N209 = N81 & N144;
  assign N210 = N81 & r_addr_i[6];
  assign N211 = N83 & N144;
  assign N212 = N83 & r_addr_i[6];
  assign N213 = N85 & N144;
  assign N214 = N85 & r_addr_i[6];
  assign N215 = N87 & N144;
  assign N216 = N87 & r_addr_i[6];
  assign N217 = N89 & N144;
  assign N218 = N89 & r_addr_i[6];
  assign N219 = N91 & N144;
  assign N220 = N91 & r_addr_i[6];
  assign N221 = N93 & N144;
  assign N222 = N93 & r_addr_i[6];
  assign N223 = N95 & N144;
  assign N224 = N95 & r_addr_i[6];
  assign N225 = N97 & N144;
  assign N226 = N97 & r_addr_i[6];
  assign N227 = N99 & N144;
  assign N228 = N99 & r_addr_i[6];
  assign N229 = N101 & N144;
  assign N230 = N101 & r_addr_i[6];
  assign N231 = N103 & N144;
  assign N232 = N103 & r_addr_i[6];
  assign N233 = N105 & N144;
  assign N234 = N105 & r_addr_i[6];
  assign N235 = N107 & N144;
  assign N236 = N107 & r_addr_i[6];
  assign N237 = N109 & N144;
  assign N238 = N109 & r_addr_i[6];
  assign N239 = N111 & N144;
  assign N240 = N111 & r_addr_i[6];
  assign N241 = N113 & N144;
  assign N242 = N113 & r_addr_i[6];
  assign N243 = N115 & N144;
  assign N244 = N115 & r_addr_i[6];
  assign N245 = N117 & N144;
  assign N246 = N117 & r_addr_i[6];
  assign N247 = N119 & N144;
  assign N248 = N119 & r_addr_i[6];
  assign N249 = N121 & N144;
  assign N250 = N121 & r_addr_i[6];
  assign N251 = N123 & N144;
  assign N252 = N123 & r_addr_i[6];
  assign N253 = N125 & N144;
  assign N254 = N125 & r_addr_i[6];
  assign N255 = N127 & N144;
  assign N256 = N127 & r_addr_i[6];
  assign N257 = N129 & N144;
  assign N258 = N129 & r_addr_i[6];
  assign N259 = N131 & N144;
  assign N260 = N131 & r_addr_i[6];
  assign N261 = N133 & N144;
  assign N262 = N133 & r_addr_i[6];
  assign N263 = N135 & N144;
  assign N264 = N135 & r_addr_i[6];
  assign N265 = N137 & N144;
  assign N266 = N137 & r_addr_i[6];
  assign N267 = N139 & N144;
  assign N268 = N139 & r_addr_i[6];
  assign N269 = N141 & N144;
  assign N270 = N141 & r_addr_i[6];
  assign N271 = N143 & N144;
  assign N272 = N143 & r_addr_i[6];
  assign N273 = ~w_v_i;

endmodule