module RocketCAM
(
  clk,
  reset,
  io_clear,
  io_clear_mask,
  io_tag,
  io_hit,
  io_hits,
  io_valid_bits,
  io_write,
  io_write_tag,
  io_write_addr
);

  input [7:0] io_clear_mask;
  input [33:0] io_tag;
  output [7:0] io_hits;
  output [7:0] io_valid_bits;
  input [33:0] io_write_tag;
  input [2:0] io_write_addr;
  input clk;
  input reset;
  input io_clear;
  input io_write;
  output io_hit;
  wire [7:0] io_hits,T8,T2,T6,T3,T4,T7,T9;
  wire io_hit,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,T14,T18,T22,T25,T30,T33,T37,T40,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N52,
  N53,N54,N55;
  wire [7:7] T45;
  reg [7:0] io_valid_bits;
  reg [33:0] T41,T38,T34,T31,T26,T23,T19,T15;
  assign T4 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << io_write_addr;
  assign T14 = T15 == io_tag;
  assign T18 = T19 == io_tag;
  assign T22 = T23 == io_tag;
  assign T25 = T26 == io_tag;
  assign T30 = T31 == io_tag;
  assign T33 = T34 == io_tag;
  assign T37 = T38 == io_tag;
  assign T40 = T41 == io_tag;

  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[7] <= N22;
    end 
  end


  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[6] <= N21;
    end 
  end


  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[5] <= N20;
    end 
  end


  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[4] <= N19;
    end 
  end


  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[3] <= N18;
    end 
  end


  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[2] <= N17;
    end 
  end


  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[1] <= N16;
    end 
  end


  always @(posedge clk) begin
    if(N14) begin
      io_valid_bits[0] <= N15;
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N39) begin
      T41[0] <= io_write_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N38) begin
      T38[0] <= io_write_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N37) begin
      T34[0] <= io_write_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N36) begin
      T31[0] <= io_write_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N35) begin
      T26[0] <= io_write_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N34) begin
      T23[0] <= io_write_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N33) begin
      T19[0] <= io_write_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[33] <= io_write_tag[33];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[32] <= io_write_tag[32];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[31] <= io_write_tag[31];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[30] <= io_write_tag[30];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[29] <= io_write_tag[29];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[28] <= io_write_tag[28];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[27] <= io_write_tag[27];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[26] <= io_write_tag[26];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[25] <= io_write_tag[25];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[24] <= io_write_tag[24];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[23] <= io_write_tag[23];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[22] <= io_write_tag[22];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[21] <= io_write_tag[21];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[20] <= io_write_tag[20];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[19] <= io_write_tag[19];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[18] <= io_write_tag[18];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[17] <= io_write_tag[17];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[16] <= io_write_tag[16];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[15] <= io_write_tag[15];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[14] <= io_write_tag[14];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[13] <= io_write_tag[13];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[12] <= io_write_tag[12];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[11] <= io_write_tag[11];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[10] <= io_write_tag[10];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[9] <= io_write_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[8] <= io_write_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[7] <= io_write_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[6] <= io_write_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[5] <= io_write_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[4] <= io_write_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[3] <= io_write_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[2] <= io_write_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[1] <= io_write_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N32) begin
      T15[0] <= io_write_tag[0];
    end 
  end

  assign N45 = io_hits[6] | io_hits[7];
  assign N46 = io_hits[5] | N45;
  assign N47 = io_hits[4] | N46;
  assign N48 = io_hits[3] | N47;
  assign N49 = io_hits[2] | N48;
  assign N50 = io_hits[1] | N49;
  assign io_hit = io_hits[0] | N50;
  assign N52 = io_write_addr[0] & io_write_addr[1];
  assign N31 = N52 & io_write_addr[2];
  assign N53 = N0 & io_write_addr[1];
  assign N0 = ~io_write_addr[0];
  assign N30 = N53 & io_write_addr[2];
  assign N54 = io_write_addr[0] & N1;
  assign N1 = ~io_write_addr[1];
  assign N29 = N54 & io_write_addr[2];
  assign N55 = N2 & N3;
  assign N2 = ~io_write_addr[0];
  assign N3 = ~io_write_addr[1];
  assign N28 = N55 & io_write_addr[2];
  assign N27 = N52 & N4;
  assign N4 = ~io_write_addr[2];
  assign N26 = N53 & N5;
  assign N5 = ~io_write_addr[2];
  assign N25 = N54 & N6;
  assign N6 = ~io_write_addr[2];
  assign N24 = N55 & N7;
  assign N7 = ~io_write_addr[2];
  assign N14 = (N8)? 1'b1 : 
               (N41)? 1'b1 : 
               (N44)? 1'b1 : 
               (N13)? 1'b0 : 1'b0;
  assign N8 = reset;
  assign { N22, N21, N20, N19, N18, N17, N16, N15 } = (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                      (N41)? T8 : 
                                                      (N44)? T2 : 1'b0;
  assign { N39, N38, N37, N36, N35, N34, N33, N32 } = (N9)? { N31, N30, N29, N28, N27, N26, N25, N24 } : 
                                                      (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = io_write;
  assign N10 = N23;
  assign T2[7] = T6[7] | T3[7];
  assign T2[6] = T6[6] | T3[6];
  assign T2[5] = T6[5] | T3[5];
  assign T2[4] = T6[4] | T3[4];
  assign T2[3] = T6[3] | T3[3];
  assign T2[2] = T6[2] | T3[2];
  assign T2[1] = T6[1] | T3[1];
  assign T2[0] = T6[0] | T3[0];
  assign T3[7] = T45[7] & T4[7];
  assign T3[6] = T45[7] & T4[6];
  assign T3[5] = T45[7] & T4[5];
  assign T3[4] = T45[7] & T4[4];
  assign T3[3] = T45[7] & T4[3];
  assign T3[2] = T45[7] & T4[2];
  assign T3[1] = T45[7] & T4[1];
  assign T3[0] = T45[7] & T4[0];
  assign T45[7] = 1'b1;
  assign T6[7] = io_valid_bits[7] & T7[7];
  assign T6[6] = io_valid_bits[6] & T7[6];
  assign T6[5] = io_valid_bits[5] & T7[5];
  assign T6[4] = io_valid_bits[4] & T7[4];
  assign T6[3] = io_valid_bits[3] & T7[3];
  assign T6[2] = io_valid_bits[2] & T7[2];
  assign T6[1] = io_valid_bits[1] & T7[1];
  assign T6[0] = io_valid_bits[0] & T7[0];
  assign T7[7] = ~T4[7];
  assign T7[6] = ~T4[6];
  assign T7[5] = ~T4[5];
  assign T7[4] = ~T4[4];
  assign T7[3] = ~T4[3];
  assign T7[2] = ~T4[2];
  assign T7[1] = ~T4[1];
  assign T7[0] = ~T4[0];
  assign T8[7] = io_valid_bits[7] & T9[7];
  assign T8[6] = io_valid_bits[6] & T9[6];
  assign T8[5] = io_valid_bits[5] & T9[5];
  assign T8[4] = io_valid_bits[4] & T9[4];
  assign T8[3] = io_valid_bits[3] & T9[3];
  assign T8[2] = io_valid_bits[2] & T9[2];
  assign T8[1] = io_valid_bits[1] & T9[1];
  assign T8[0] = io_valid_bits[0] & T9[0];
  assign T9[7] = ~io_clear_mask[7];
  assign T9[6] = ~io_clear_mask[6];
  assign T9[5] = ~io_clear_mask[5];
  assign T9[4] = ~io_clear_mask[4];
  assign T9[3] = ~io_clear_mask[3];
  assign T9[2] = ~io_clear_mask[2];
  assign T9[1] = ~io_clear_mask[1];
  assign T9[0] = ~io_clear_mask[0];
  assign io_hits[0] = io_valid_bits[0] & T14;
  assign io_hits[1] = io_valid_bits[1] & T18;
  assign io_hits[2] = io_valid_bits[2] & T22;
  assign io_hits[3] = io_valid_bits[3] & T25;
  assign io_hits[4] = io_valid_bits[4] & T30;
  assign io_hits[5] = io_valid_bits[5] & T33;
  assign io_hits[6] = io_valid_bits[6] & T37;
  assign io_hits[7] = io_valid_bits[7] & T40;
  assign N11 = io_clear | reset;
  assign N12 = io_write | N11;
  assign N13 = ~N12;
  assign N23 = ~io_write;
  assign N40 = ~reset;
  assign N41 = io_clear & N40;
  assign N42 = ~io_clear;
  assign N43 = N40 & N42;
  assign N44 = io_write & N43;

endmodule