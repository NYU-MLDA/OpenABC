module bp_fe_bht_bht_indx_width_p5
(
  clk_i,
  en_i,
  reset_i,
  idx_r_i,
  idx_w_i,
  r_v_i,
  w_v_i,
  correct_i,
  predict_o
);

  input [4:0] idx_r_i;
  input [4:0] idx_w_i;
  input clk_i;
  input en_i;
  input reset_i;
  input r_v_i;
  input w_v_i;
  input correct_i;
  output predict_o;
  wire predict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413;
  reg [63:0] mem;
  assign predict_o = (N52)? mem[1] : 
                     (N54)? mem[3] : 
                     (N56)? mem[5] : 
                     (N58)? mem[7] : 
                     (N60)? mem[9] : 
                     (N62)? mem[11] : 
                     (N64)? mem[13] : 
                     (N66)? mem[15] : 
                     (N68)? mem[17] : 
                     (N70)? mem[19] : 
                     (N72)? mem[21] : 
                     (N74)? mem[23] : 
                     (N76)? mem[25] : 
                     (N78)? mem[27] : 
                     (N80)? mem[29] : 
                     (N82)? mem[31] : 
                     (N53)? mem[33] : 
                     (N55)? mem[35] : 
                     (N57)? mem[37] : 
                     (N59)? mem[39] : 
                     (N61)? mem[41] : 
                     (N63)? mem[43] : 
                     (N65)? mem[45] : 
                     (N67)? mem[47] : 
                     (N69)? mem[49] : 
                     (N71)? mem[51] : 
                     (N73)? mem[53] : 
                     (N75)? mem[55] : 
                     (N77)? mem[57] : 
                     (N79)? mem[59] : 
                     (N81)? mem[61] : 
                     (N83)? mem[63] : 1'b0;
  assign N87 = (N147)? mem[1] : 
               (N148)? mem[3] : 
               (N149)? mem[5] : 
               (N150)? mem[7] : 
               (N151)? mem[9] : 
               (N152)? mem[11] : 
               (N153)? mem[13] : 
               (N154)? mem[15] : 
               (N155)? mem[17] : 
               (N156)? mem[19] : 
               (N157)? mem[21] : 
               (N158)? mem[23] : 
               (N159)? mem[25] : 
               (N160)? mem[27] : 
               (N161)? mem[29] : 
               (N162)? mem[31] : 
               (N123)? mem[33] : 
               (N125)? mem[35] : 
               (N127)? mem[37] : 
               (N129)? mem[39] : 
               (N131)? mem[41] : 
               (N133)? mem[43] : 
               (N135)? mem[45] : 
               (N137)? mem[47] : 
               (N272)? mem[49] : 
               (N274)? mem[51] : 
               (N276)? mem[53] : 
               (N278)? mem[55] : 
               (N280)? mem[57] : 
               (N282)? mem[59] : 
               (N284)? mem[61] : 
               (N286)? mem[63] : 1'b0;
  assign N88 = (N147)? mem[0] : 
               (N148)? mem[2] : 
               (N149)? mem[4] : 
               (N150)? mem[6] : 
               (N151)? mem[8] : 
               (N152)? mem[10] : 
               (N153)? mem[12] : 
               (N154)? mem[14] : 
               (N155)? mem[16] : 
               (N156)? mem[18] : 
               (N157)? mem[20] : 
               (N158)? mem[22] : 
               (N159)? mem[24] : 
               (N160)? mem[26] : 
               (N161)? mem[28] : 
               (N162)? mem[30] : 
               (N123)? mem[32] : 
               (N125)? mem[34] : 
               (N127)? mem[36] : 
               (N129)? mem[38] : 
               (N131)? mem[40] : 
               (N133)? mem[42] : 
               (N135)? mem[44] : 
               (N137)? mem[46] : 
               (N272)? mem[48] : 
               (N274)? mem[50] : 
               (N276)? mem[52] : 
               (N278)? mem[54] : 
               (N280)? mem[56] : 
               (N282)? mem[58] : 
               (N284)? mem[60] : 
               (N286)? mem[62] : 1'b0;
  assign N92 = N89 & N90;
  assign N93 = N92 & N91;
  assign N94 = correct_i | N87;
  assign N95 = N94 | N91;
  assign N97 = correct_i | N90;
  assign N98 = N97 | N88;
  assign N100 = N97 | N91;
  assign N102 = N89 | N87;
  assign N103 = N102 | N88;
  assign N105 = N102 | N91;
  assign N107 = N89 | N90;
  assign N108 = N107 | N88;
  assign N110 = correct_i & N87;
  assign N111 = N110 & N88;
  assign N146 = (N122)? mem[1] : 
                (N124)? mem[3] : 
                (N126)? mem[5] : 
                (N128)? mem[7] : 
                (N130)? mem[9] : 
                (N132)? mem[11] : 
                (N134)? mem[13] : 
                (N136)? mem[15] : 
                (N138)? mem[17] : 
                (N139)? mem[19] : 
                (N140)? mem[21] : 
                (N141)? mem[23] : 
                (N142)? mem[25] : 
                (N143)? mem[27] : 
                (N144)? mem[29] : 
                (N145)? mem[31] : 
                (N123)? mem[33] : 
                (N125)? mem[35] : 
                (N127)? mem[37] : 
                (N129)? mem[39] : 
                (N131)? mem[41] : 
                (N133)? mem[43] : 
                (N135)? mem[45] : 
                (N137)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N163 = (N147)? mem[0] : 
                (N148)? mem[2] : 
                (N149)? mem[4] : 
                (N150)? mem[6] : 
                (N151)? mem[8] : 
                (N152)? mem[10] : 
                (N153)? mem[12] : 
                (N154)? mem[14] : 
                (N155)? mem[16] : 
                (N156)? mem[18] : 
                (N157)? mem[20] : 
                (N158)? mem[22] : 
                (N159)? mem[24] : 
                (N160)? mem[26] : 
                (N161)? mem[28] : 
                (N162)? mem[30] : 
                (N123)? mem[32] : 
                (N125)? mem[34] : 
                (N127)? mem[36] : 
                (N129)? mem[38] : 
                (N131)? mem[40] : 
                (N133)? mem[42] : 
                (N135)? mem[44] : 
                (N137)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N205 = (N197)? mem[1] : 
                (N198)? mem[3] : 
                (N199)? mem[5] : 
                (N200)? mem[7] : 
                (N201)? mem[9] : 
                (N202)? mem[11] : 
                (N203)? mem[13] : 
                (N204)? mem[15] : 
                (N155)? mem[17] : 
                (N156)? mem[19] : 
                (N157)? mem[21] : 
                (N158)? mem[23] : 
                (N159)? mem[25] : 
                (N160)? mem[27] : 
                (N161)? mem[29] : 
                (N162)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N214 = (N206)? mem[0] : 
                (N207)? mem[2] : 
                (N208)? mem[4] : 
                (N209)? mem[6] : 
                (N210)? mem[8] : 
                (N211)? mem[10] : 
                (N212)? mem[12] : 
                (N213)? mem[14] : 
                (N138)? mem[16] : 
                (N139)? mem[18] : 
                (N140)? mem[20] : 
                (N141)? mem[22] : 
                (N142)? mem[24] : 
                (N143)? mem[26] : 
                (N144)? mem[28] : 
                (N145)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N216 = (N206)? mem[1] : 
                (N207)? mem[3] : 
                (N208)? mem[5] : 
                (N209)? mem[7] : 
                (N210)? mem[9] : 
                (N211)? mem[11] : 
                (N212)? mem[13] : 
                (N213)? mem[15] : 
                (N138)? mem[17] : 
                (N139)? mem[19] : 
                (N140)? mem[21] : 
                (N141)? mem[23] : 
                (N142)? mem[25] : 
                (N143)? mem[27] : 
                (N144)? mem[29] : 
                (N145)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N217 = (N206)? mem[0] : 
                (N207)? mem[2] : 
                (N208)? mem[4] : 
                (N209)? mem[6] : 
                (N210)? mem[8] : 
                (N211)? mem[10] : 
                (N212)? mem[12] : 
                (N213)? mem[14] : 
                (N138)? mem[16] : 
                (N139)? mem[18] : 
                (N140)? mem[20] : 
                (N141)? mem[22] : 
                (N142)? mem[24] : 
                (N143)? mem[26] : 
                (N144)? mem[28] : 
                (N145)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N219 = (N206)? mem[1] : 
                (N207)? mem[3] : 
                (N208)? mem[5] : 
                (N209)? mem[7] : 
                (N210)? mem[9] : 
                (N211)? mem[11] : 
                (N212)? mem[13] : 
                (N213)? mem[15] : 
                (N138)? mem[17] : 
                (N139)? mem[19] : 
                (N140)? mem[21] : 
                (N141)? mem[23] : 
                (N142)? mem[25] : 
                (N143)? mem[27] : 
                (N144)? mem[29] : 
                (N145)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N220 = (N206)? mem[0] : 
                (N207)? mem[2] : 
                (N208)? mem[4] : 
                (N209)? mem[6] : 
                (N210)? mem[8] : 
                (N211)? mem[10] : 
                (N212)? mem[12] : 
                (N213)? mem[14] : 
                (N138)? mem[16] : 
                (N139)? mem[18] : 
                (N140)? mem[20] : 
                (N141)? mem[22] : 
                (N142)? mem[24] : 
                (N143)? mem[26] : 
                (N144)? mem[28] : 
                (N145)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N222 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N223 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N287 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N288 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N290 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N291 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N292 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N293 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N397 = idx_w_i[3] & idx_w_i[4];
  assign N398 = N0 & idx_w_i[4];
  assign N0 = ~idx_w_i[3];
  assign N399 = idx_w_i[3] & N1;
  assign N1 = ~idx_w_i[4];
  assign N400 = N2 & N3;
  assign N2 = ~idx_w_i[3];
  assign N3 = ~idx_w_i[4];
  assign N401 = ~idx_w_i[2];
  assign N402 = idx_w_i[0] & idx_w_i[1];
  assign N403 = N4 & idx_w_i[1];
  assign N4 = ~idx_w_i[0];
  assign N404 = idx_w_i[0] & N5;
  assign N5 = ~idx_w_i[1];
  assign N405 = N6 & N7;
  assign N6 = ~idx_w_i[0];
  assign N7 = ~idx_w_i[1];
  assign N406 = idx_w_i[2] & N402;
  assign N407 = idx_w_i[2] & N403;
  assign N408 = idx_w_i[2] & N404;
  assign N409 = idx_w_i[2] & N405;
  assign N410 = N401 & N402;
  assign N411 = N401 & N403;
  assign N412 = N401 & N404;
  assign N413 = N401 & N405;
  assign N195 = N397 & N406;
  assign N194 = N397 & N407;
  assign N193 = N397 & N408;
  assign N192 = N397 & N409;
  assign N191 = N397 & N410;
  assign N190 = N397 & N411;
  assign N189 = N397 & N412;
  assign N188 = N397 & N413;
  assign N187 = N398 & N406;
  assign N186 = N398 & N407;
  assign N185 = N398 & N408;
  assign N184 = N398 & N409;
  assign N183 = N398 & N410;
  assign N182 = N398 & N411;
  assign N181 = N398 & N412;
  assign N180 = N398 & N413;
  assign N179 = N399 & N406;
  assign N178 = N399 & N407;
  assign N177 = N399 & N408;
  assign N176 = N399 & N409;
  assign N175 = N399 & N410;
  assign N174 = N399 & N411;
  assign N173 = N399 & N412;
  assign N172 = N399 & N413;
  assign N171 = N400 & N406;
  assign N170 = N400 & N407;
  assign N169 = N400 & N408;
  assign N168 = N400 & N409;
  assign N167 = N400 & N410;
  assign N166 = N400 & N411;
  assign N165 = N400 & N412;
  assign N164 = N400 & N413;
  assign { N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N295 } = (N8)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N9)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N10)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N11)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N12)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N13)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N14)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N15)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 1'b0;
  assign N8 = N93;
  assign N9 = N96;
  assign N10 = N99;
  assign N11 = N101;
  assign N12 = N104;
  assign N13 = N106;
  assign N14 = N109;
  assign N15 = N111;
  assign { N297, N296 } = (N8)? { N196, 1'b1 } : 
                          (N9)? { N215, 1'b1 } : 
                          (N10)? { N218, 1'b1 } : 
                          (N11)? { N221, 1'b1 } : 
                          (N12)? { N222, N223 } : 
                          (N13)? { N287, N289 } : 
                          (N14)? { N290, N291 } : 
                          (N15)? { N292, N294 } : 1'b0;
  assign { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N329 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N396)? { N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N295 } : 
                                                                                                                                                                                                              (N86)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = reset_i;
  assign { N331, N330 } = (N16)? { 1'b0, 1'b1 } : 
                          (N396)? { N297, N296 } : 1'b0;
  assign { N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363 } = (N17)? { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N329 } : 
                                                                                                                                                                                                              (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = en_i;
  assign N18 = N84;
  assign N19 = ~idx_r_i[0];
  assign N20 = ~idx_r_i[1];
  assign N21 = N19 & N20;
  assign N22 = N19 & idx_r_i[1];
  assign N23 = idx_r_i[0] & N20;
  assign N24 = idx_r_i[0] & idx_r_i[1];
  assign N25 = ~idx_r_i[2];
  assign N26 = N21 & N25;
  assign N27 = N21 & idx_r_i[2];
  assign N28 = N23 & N25;
  assign N29 = N23 & idx_r_i[2];
  assign N30 = N22 & N25;
  assign N31 = N22 & idx_r_i[2];
  assign N32 = N24 & N25;
  assign N33 = N24 & idx_r_i[2];
  assign N34 = ~idx_r_i[3];
  assign N35 = N26 & N34;
  assign N36 = N26 & idx_r_i[3];
  assign N37 = N28 & N34;
  assign N38 = N28 & idx_r_i[3];
  assign N39 = N30 & N34;
  assign N40 = N30 & idx_r_i[3];
  assign N41 = N32 & N34;
  assign N42 = N32 & idx_r_i[3];
  assign N43 = N27 & N34;
  assign N44 = N27 & idx_r_i[3];
  assign N45 = N29 & N34;
  assign N46 = N29 & idx_r_i[3];
  assign N47 = N31 & N34;
  assign N48 = N31 & idx_r_i[3];
  assign N49 = N33 & N34;
  assign N50 = N33 & idx_r_i[3];
  assign N51 = ~idx_r_i[4];
  assign N52 = N35 & N51;
  assign N53 = N35 & idx_r_i[4];
  assign N54 = N37 & N51;
  assign N55 = N37 & idx_r_i[4];
  assign N56 = N39 & N51;
  assign N57 = N39 & idx_r_i[4];
  assign N58 = N41 & N51;
  assign N59 = N41 & idx_r_i[4];
  assign N60 = N43 & N51;
  assign N61 = N43 & idx_r_i[4];
  assign N62 = N45 & N51;
  assign N63 = N45 & idx_r_i[4];
  assign N64 = N47 & N51;
  assign N65 = N47 & idx_r_i[4];
  assign N66 = N49 & N51;
  assign N67 = N49 & idx_r_i[4];
  assign N68 = N36 & N51;
  assign N69 = N36 & idx_r_i[4];
  assign N70 = N38 & N51;
  assign N71 = N38 & idx_r_i[4];
  assign N72 = N40 & N51;
  assign N73 = N40 & idx_r_i[4];
  assign N74 = N42 & N51;
  assign N75 = N42 & idx_r_i[4];
  assign N76 = N44 & N51;
  assign N77 = N44 & idx_r_i[4];
  assign N78 = N46 & N51;
  assign N79 = N46 & idx_r_i[4];
  assign N80 = N48 & N51;
  assign N81 = N48 & idx_r_i[4];
  assign N82 = N50 & N51;
  assign N83 = N50 & idx_r_i[4];
  assign N84 = ~en_i;
  assign N85 = w_v_i | reset_i;
  assign N86 = ~N85;
  assign N89 = ~correct_i;
  assign N90 = ~N87;
  assign N91 = ~N88;
  assign N96 = ~N95;
  assign N99 = ~N98;
  assign N101 = ~N100;
  assign N104 = ~N103;
  assign N106 = ~N105;
  assign N109 = ~N108;
  assign N112 = ~idx_w_i[3];
  assign N113 = N231 & N112;
  assign N114 = N233 & N112;
  assign N115 = N235 & N112;
  assign N116 = N237 & N112;
  assign N117 = N232 & N112;
  assign N118 = N234 & N112;
  assign N119 = N236 & N112;
  assign N120 = N238 & N112;
  assign N121 = ~idx_w_i[4];
  assign N122 = N113 & N121;
  assign N123 = N113 & idx_w_i[4];
  assign N124 = N114 & N121;
  assign N125 = N114 & idx_w_i[4];
  assign N126 = N115 & N121;
  assign N127 = N115 & idx_w_i[4];
  assign N128 = N116 & N121;
  assign N129 = N116 & idx_w_i[4];
  assign N130 = N117 & N121;
  assign N131 = N117 & idx_w_i[4];
  assign N132 = N118 & N121;
  assign N133 = N118 & idx_w_i[4];
  assign N134 = N119 & N121;
  assign N135 = N119 & idx_w_i[4];
  assign N136 = N120 & N121;
  assign N137 = N120 & idx_w_i[4];
  assign N138 = N240 & N121;
  assign N139 = N242 & N121;
  assign N140 = N244 & N121;
  assign N141 = N246 & N121;
  assign N142 = N248 & N121;
  assign N143 = N250 & N121;
  assign N144 = N252 & N121;
  assign N145 = N254 & N121;
  assign N147 = N113 & N121;
  assign N148 = N114 & N121;
  assign N149 = N115 & N121;
  assign N150 = N116 & N121;
  assign N151 = N117 & N121;
  assign N152 = N118 & N121;
  assign N153 = N119 & N121;
  assign N154 = N120 & N121;
  assign N155 = N240 & N121;
  assign N156 = N242 & N121;
  assign N157 = N244 & N121;
  assign N158 = N246 & N121;
  assign N159 = N248 & N121;
  assign N160 = N250 & N121;
  assign N161 = N252 & N121;
  assign N162 = N254 & N121;
  assign N196 = N146 ^ N163;
  assign N197 = N239 & N121;
  assign N198 = N241 & N121;
  assign N199 = N243 & N121;
  assign N200 = N245 & N121;
  assign N201 = N247 & N121;
  assign N202 = N249 & N121;
  assign N203 = N251 & N121;
  assign N204 = N253 & N121;
  assign N206 = N239 & N121;
  assign N207 = N241 & N121;
  assign N208 = N243 & N121;
  assign N209 = N245 & N121;
  assign N210 = N247 & N121;
  assign N211 = N249 & N121;
  assign N212 = N251 & N121;
  assign N213 = N253 & N121;
  assign N215 = N205 ^ N214;
  assign N218 = N216 ^ N217;
  assign N221 = N219 ^ N220;
  assign N224 = ~idx_w_i[0];
  assign N225 = ~idx_w_i[1];
  assign N226 = N224 & N225;
  assign N227 = N224 & idx_w_i[1];
  assign N228 = idx_w_i[0] & N225;
  assign N229 = idx_w_i[0] & idx_w_i[1];
  assign N230 = ~idx_w_i[2];
  assign N231 = N226 & N230;
  assign N232 = N226 & idx_w_i[2];
  assign N233 = N228 & N230;
  assign N234 = N228 & idx_w_i[2];
  assign N235 = N227 & N230;
  assign N236 = N227 & idx_w_i[2];
  assign N237 = N229 & N230;
  assign N238 = N229 & idx_w_i[2];
  assign N239 = N231 & N112;
  assign N240 = N231 & idx_w_i[3];
  assign N241 = N233 & N112;
  assign N242 = N233 & idx_w_i[3];
  assign N243 = N235 & N112;
  assign N244 = N235 & idx_w_i[3];
  assign N245 = N237 & N112;
  assign N246 = N237 & idx_w_i[3];
  assign N247 = N232 & N112;
  assign N248 = N232 & idx_w_i[3];
  assign N249 = N234 & N112;
  assign N250 = N234 & idx_w_i[3];
  assign N251 = N236 & N112;
  assign N252 = N236 & idx_w_i[3];
  assign N253 = N238 & N112;
  assign N254 = N238 & idx_w_i[3];
  assign N255 = N239 & N121;
  assign N256 = N239 & idx_w_i[4];
  assign N257 = N241 & N121;
  assign N258 = N241 & idx_w_i[4];
  assign N259 = N243 & N121;
  assign N260 = N243 & idx_w_i[4];
  assign N261 = N245 & N121;
  assign N262 = N245 & idx_w_i[4];
  assign N263 = N247 & N121;
  assign N264 = N247 & idx_w_i[4];
  assign N265 = N249 & N121;
  assign N266 = N249 & idx_w_i[4];
  assign N267 = N251 & N121;
  assign N268 = N251 & idx_w_i[4];
  assign N269 = N253 & N121;
  assign N270 = N253 & idx_w_i[4];
  assign N271 = N240 & N121;
  assign N272 = N240 & idx_w_i[4];
  assign N273 = N242 & N121;
  assign N274 = N242 & idx_w_i[4];
  assign N275 = N244 & N121;
  assign N276 = N244 & idx_w_i[4];
  assign N277 = N246 & N121;
  assign N278 = N246 & idx_w_i[4];
  assign N279 = N248 & N121;
  assign N280 = N248 & idx_w_i[4];
  assign N281 = N250 & N121;
  assign N282 = N250 & idx_w_i[4];
  assign N283 = N252 & N121;
  assign N284 = N252 & idx_w_i[4];
  assign N285 = N254 & N121;
  assign N286 = N254 & idx_w_i[4];
  assign N289 = ~N288;
  assign N294 = ~N293;
  assign N395 = ~reset_i;
  assign N396 = w_v_i & N395;

  always @(posedge clk_i) begin
    if(N394) begin
      { mem[63:62] } <= { N331, N330 };
    end 
    if(N393) begin
      { mem[61:60] } <= { N331, N330 };
    end 
    if(N392) begin
      { mem[59:58] } <= { N331, N330 };
    end 
    if(N391) begin
      { mem[57:56] } <= { N331, N330 };
    end 
    if(N390) begin
      { mem[55:54] } <= { N331, N330 };
    end 
    if(N389) begin
      { mem[53:52] } <= { N331, N330 };
    end 
    if(N388) begin
      { mem[51:50] } <= { N331, N330 };
    end 
    if(N387) begin
      { mem[49:48] } <= { N331, N330 };
    end 
    if(N386) begin
      { mem[47:46] } <= { N331, N330 };
    end 
    if(N385) begin
      { mem[45:44] } <= { N331, N330 };
    end 
    if(N384) begin
      { mem[43:42] } <= { N331, N330 };
    end 
    if(N383) begin
      { mem[41:40] } <= { N331, N330 };
    end 
    if(N382) begin
      { mem[39:38] } <= { N331, N330 };
    end 
    if(N381) begin
      { mem[37:36] } <= { N331, N330 };
    end 
    if(N380) begin
      { mem[35:34] } <= { N331, N330 };
    end 
    if(N379) begin
      { mem[33:32] } <= { N331, N330 };
    end 
    if(N378) begin
      { mem[31:30] } <= { N331, N330 };
    end 
    if(N377) begin
      { mem[29:28] } <= { N331, N330 };
    end 
    if(N376) begin
      { mem[27:26] } <= { N331, N330 };
    end 
    if(N375) begin
      { mem[25:24] } <= { N331, N330 };
    end 
    if(N374) begin
      { mem[23:22] } <= { N331, N330 };
    end 
    if(N373) begin
      { mem[21:20] } <= { N331, N330 };
    end 
    if(N372) begin
      { mem[19:18] } <= { N331, N330 };
    end 
    if(N371) begin
      { mem[17:16] } <= { N331, N330 };
    end 
    if(N370) begin
      { mem[15:14] } <= { N331, N330 };
    end 
    if(N369) begin
      { mem[13:12] } <= { N331, N330 };
    end 
    if(N368) begin
      { mem[11:10] } <= { N331, N330 };
    end 
    if(N367) begin
      { mem[9:8] } <= { N331, N330 };
    end 
    if(N366) begin
      { mem[7:6] } <= { N331, N330 };
    end 
    if(N365) begin
      { mem[5:4] } <= { N331, N330 };
    end 
    if(N364) begin
      { mem[3:2] } <= { N331, N330 };
    end 
    if(N363) begin
      { mem[1:0] } <= { N331, N330 };
    end 
  end


endmodule