module tag_cmp_4_0000000c_00000008
(
  clk_i,
  rst_ni,
  req_i,
  gnt_o,
  addr_i,
  wdata_i,
  we_i,
  be_i,
  rdata_o,
  tag_i,
  hit_way_o,
  req_o,
  addr_o,
  wdata_o,
  we_o,
  be_o,
  rdata_i
);

  input [31:0] req_i;
  output [3:0] gnt_o;
  input [47:0] addr_i;
  input [695:0] wdata_i;
  input [3:0] we_i;
  input [119:0] be_i;
  output [1391:0] rdata_o;
  input [175:0] tag_i;
  output [7:0] hit_way_o;
  output [7:0] req_o;
  output [11:0] addr_o;
  output [173:0] wdata_o;
  output [29:0] be_o;
  input [1391:0] rdata_i;
  input clk_i;
  input rst_ni;
  output we_o;
  wire [3:0] gnt_o,id_d;
  wire [1391:0] rdata_o;
  wire [7:0] hit_way_o,req_o;
  wire [11:0] addr_o;
  wire [173:0] wdata_o;
  wire [29:0] be_o;
  wire we_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,
  N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,
  N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,
  N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,
  N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
  N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,
  N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,
  N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,
  N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,
  N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,
  N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,
  N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,
  N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,
  N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,
  N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,
  N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,
  N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,
  N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,
  N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,
  N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,
  N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,
  N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,
  N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,
  N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,
  N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,
  N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,
  N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,
  N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,
  N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,
  N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,
  N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,
  N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,
  N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,
  N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,
  N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,
  N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,
  N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,
  N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,
  N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,
  N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,
  N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,
  N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,
  N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,
  N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,
  N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,
  N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,
  N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,
  N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,
  N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,
  N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,
  N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343;
  wire [43:0] sel_tag;
  reg [3:0] id_q;
  assign gnt_o[0] = 1'b1;
  assign rdata_o[1391] = rdata_i[1391];
  assign rdata_o[1390] = rdata_i[1390];
  assign rdata_o[1389] = rdata_i[1389];
  assign rdata_o[1388] = rdata_i[1388];
  assign rdata_o[1387] = rdata_i[1387];
  assign rdata_o[1386] = rdata_i[1386];
  assign rdata_o[1385] = rdata_i[1385];
  assign rdata_o[1384] = rdata_i[1384];
  assign rdata_o[1383] = rdata_i[1383];
  assign rdata_o[1382] = rdata_i[1382];
  assign rdata_o[1381] = rdata_i[1381];
  assign rdata_o[1380] = rdata_i[1380];
  assign rdata_o[1379] = rdata_i[1379];
  assign rdata_o[1378] = rdata_i[1378];
  assign rdata_o[1377] = rdata_i[1377];
  assign rdata_o[1376] = rdata_i[1376];
  assign rdata_o[1375] = rdata_i[1375];
  assign rdata_o[1374] = rdata_i[1374];
  assign rdata_o[1373] = rdata_i[1373];
  assign rdata_o[1372] = rdata_i[1372];
  assign rdata_o[1371] = rdata_i[1371];
  assign rdata_o[1370] = rdata_i[1370];
  assign rdata_o[1369] = rdata_i[1369];
  assign rdata_o[1368] = rdata_i[1368];
  assign rdata_o[1367] = rdata_i[1367];
  assign rdata_o[1366] = rdata_i[1366];
  assign rdata_o[1365] = rdata_i[1365];
  assign rdata_o[1364] = rdata_i[1364];
  assign rdata_o[1363] = rdata_i[1363];
  assign rdata_o[1362] = rdata_i[1362];
  assign rdata_o[1361] = rdata_i[1361];
  assign rdata_o[1360] = rdata_i[1360];
  assign rdata_o[1359] = rdata_i[1359];
  assign rdata_o[1358] = rdata_i[1358];
  assign rdata_o[1357] = rdata_i[1357];
  assign rdata_o[1356] = rdata_i[1356];
  assign rdata_o[1355] = rdata_i[1355];
  assign rdata_o[1354] = rdata_i[1354];
  assign rdata_o[1353] = rdata_i[1353];
  assign rdata_o[1352] = rdata_i[1352];
  assign rdata_o[1351] = rdata_i[1351];
  assign rdata_o[1350] = rdata_i[1350];
  assign rdata_o[1349] = rdata_i[1349];
  assign rdata_o[1348] = rdata_i[1348];
  assign rdata_o[1347] = rdata_i[1347];
  assign rdata_o[1346] = rdata_i[1346];
  assign rdata_o[1345] = rdata_i[1345];
  assign rdata_o[1344] = rdata_i[1344];
  assign rdata_o[1343] = rdata_i[1343];
  assign rdata_o[1342] = rdata_i[1342];
  assign rdata_o[1341] = rdata_i[1341];
  assign rdata_o[1340] = rdata_i[1340];
  assign rdata_o[1339] = rdata_i[1339];
  assign rdata_o[1338] = rdata_i[1338];
  assign rdata_o[1337] = rdata_i[1337];
  assign rdata_o[1336] = rdata_i[1336];
  assign rdata_o[1335] = rdata_i[1335];
  assign rdata_o[1334] = rdata_i[1334];
  assign rdata_o[1333] = rdata_i[1333];
  assign rdata_o[1332] = rdata_i[1332];
  assign rdata_o[1331] = rdata_i[1331];
  assign rdata_o[1330] = rdata_i[1330];
  assign rdata_o[1329] = rdata_i[1329];
  assign rdata_o[1328] = rdata_i[1328];
  assign rdata_o[1327] = rdata_i[1327];
  assign rdata_o[1326] = rdata_i[1326];
  assign rdata_o[1325] = rdata_i[1325];
  assign rdata_o[1324] = rdata_i[1324];
  assign rdata_o[1323] = rdata_i[1323];
  assign rdata_o[1322] = rdata_i[1322];
  assign rdata_o[1321] = rdata_i[1321];
  assign rdata_o[1320] = rdata_i[1320];
  assign rdata_o[1319] = rdata_i[1319];
  assign rdata_o[1318] = rdata_i[1318];
  assign rdata_o[1317] = rdata_i[1317];
  assign rdata_o[1316] = rdata_i[1316];
  assign rdata_o[1315] = rdata_i[1315];
  assign rdata_o[1314] = rdata_i[1314];
  assign rdata_o[1313] = rdata_i[1313];
  assign rdata_o[1312] = rdata_i[1312];
  assign rdata_o[1311] = rdata_i[1311];
  assign rdata_o[1310] = rdata_i[1310];
  assign rdata_o[1309] = rdata_i[1309];
  assign rdata_o[1308] = rdata_i[1308];
  assign rdata_o[1307] = rdata_i[1307];
  assign rdata_o[1306] = rdata_i[1306];
  assign rdata_o[1305] = rdata_i[1305];
  assign rdata_o[1304] = rdata_i[1304];
  assign rdata_o[1303] = rdata_i[1303];
  assign rdata_o[1302] = rdata_i[1302];
  assign rdata_o[1301] = rdata_i[1301];
  assign rdata_o[1300] = rdata_i[1300];
  assign rdata_o[1299] = rdata_i[1299];
  assign rdata_o[1298] = rdata_i[1298];
  assign rdata_o[1297] = rdata_i[1297];
  assign rdata_o[1296] = rdata_i[1296];
  assign rdata_o[1295] = rdata_i[1295];
  assign rdata_o[1294] = rdata_i[1294];
  assign rdata_o[1293] = rdata_i[1293];
  assign rdata_o[1292] = rdata_i[1292];
  assign rdata_o[1291] = rdata_i[1291];
  assign rdata_o[1290] = rdata_i[1290];
  assign rdata_o[1289] = rdata_i[1289];
  assign rdata_o[1288] = rdata_i[1288];
  assign rdata_o[1287] = rdata_i[1287];
  assign rdata_o[1286] = rdata_i[1286];
  assign rdata_o[1285] = rdata_i[1285];
  assign rdata_o[1284] = rdata_i[1284];
  assign rdata_o[1283] = rdata_i[1283];
  assign rdata_o[1282] = rdata_i[1282];
  assign rdata_o[1281] = rdata_i[1281];
  assign rdata_o[1280] = rdata_i[1280];
  assign rdata_o[1279] = rdata_i[1279];
  assign rdata_o[1278] = rdata_i[1278];
  assign rdata_o[1277] = rdata_i[1277];
  assign rdata_o[1276] = rdata_i[1276];
  assign rdata_o[1275] = rdata_i[1275];
  assign rdata_o[1274] = rdata_i[1274];
  assign rdata_o[1273] = rdata_i[1273];
  assign rdata_o[1272] = rdata_i[1272];
  assign rdata_o[1271] = rdata_i[1271];
  assign rdata_o[1270] = rdata_i[1270];
  assign rdata_o[1269] = rdata_i[1269];
  assign rdata_o[1268] = rdata_i[1268];
  assign rdata_o[1267] = rdata_i[1267];
  assign rdata_o[1266] = rdata_i[1266];
  assign rdata_o[1265] = rdata_i[1265];
  assign rdata_o[1264] = rdata_i[1264];
  assign rdata_o[1263] = rdata_i[1263];
  assign rdata_o[1262] = rdata_i[1262];
  assign rdata_o[1261] = rdata_i[1261];
  assign rdata_o[1260] = rdata_i[1260];
  assign rdata_o[1259] = rdata_i[1259];
  assign rdata_o[1258] = rdata_i[1258];
  assign rdata_o[1257] = rdata_i[1257];
  assign rdata_o[1256] = rdata_i[1256];
  assign rdata_o[1255] = rdata_i[1255];
  assign rdata_o[1254] = rdata_i[1254];
  assign rdata_o[1253] = rdata_i[1253];
  assign rdata_o[1252] = rdata_i[1252];
  assign rdata_o[1251] = rdata_i[1251];
  assign rdata_o[1250] = rdata_i[1250];
  assign rdata_o[1249] = rdata_i[1249];
  assign rdata_o[1248] = rdata_i[1248];
  assign rdata_o[1247] = rdata_i[1247];
  assign rdata_o[1246] = rdata_i[1246];
  assign rdata_o[1245] = rdata_i[1245];
  assign rdata_o[1244] = rdata_i[1244];
  assign rdata_o[1243] = rdata_i[1243];
  assign rdata_o[1242] = rdata_i[1242];
  assign rdata_o[1241] = rdata_i[1241];
  assign rdata_o[1240] = rdata_i[1240];
  assign rdata_o[1239] = rdata_i[1239];
  assign rdata_o[1238] = rdata_i[1238];
  assign rdata_o[1237] = rdata_i[1237];
  assign rdata_o[1236] = rdata_i[1236];
  assign rdata_o[1235] = rdata_i[1235];
  assign rdata_o[1234] = rdata_i[1234];
  assign rdata_o[1233] = rdata_i[1233];
  assign rdata_o[1232] = rdata_i[1232];
  assign rdata_o[1231] = rdata_i[1231];
  assign rdata_o[1230] = rdata_i[1230];
  assign rdata_o[1229] = rdata_i[1229];
  assign rdata_o[1228] = rdata_i[1228];
  assign rdata_o[1227] = rdata_i[1227];
  assign rdata_o[1226] = rdata_i[1226];
  assign rdata_o[1225] = rdata_i[1225];
  assign rdata_o[1224] = rdata_i[1224];
  assign rdata_o[1223] = rdata_i[1223];
  assign rdata_o[1222] = rdata_i[1222];
  assign rdata_o[1221] = rdata_i[1221];
  assign rdata_o[1220] = rdata_i[1220];
  assign rdata_o[1219] = rdata_i[1219];
  assign rdata_o[1218] = rdata_i[1218];
  assign rdata_o[1217] = rdata_i[1217];
  assign rdata_o[1216] = rdata_i[1216];
  assign rdata_o[1215] = rdata_i[1215];
  assign rdata_o[1214] = rdata_i[1214];
  assign rdata_o[1213] = rdata_i[1213];
  assign rdata_o[1212] = rdata_i[1212];
  assign rdata_o[1211] = rdata_i[1211];
  assign rdata_o[1210] = rdata_i[1210];
  assign rdata_o[1209] = rdata_i[1209];
  assign rdata_o[1208] = rdata_i[1208];
  assign rdata_o[1207] = rdata_i[1207];
  assign rdata_o[1206] = rdata_i[1206];
  assign rdata_o[1205] = rdata_i[1205];
  assign rdata_o[1204] = rdata_i[1204];
  assign rdata_o[1203] = rdata_i[1203];
  assign rdata_o[1202] = rdata_i[1202];
  assign rdata_o[1201] = rdata_i[1201];
  assign rdata_o[1200] = rdata_i[1200];
  assign rdata_o[1199] = rdata_i[1199];
  assign rdata_o[1198] = rdata_i[1198];
  assign rdata_o[1197] = rdata_i[1197];
  assign rdata_o[1196] = rdata_i[1196];
  assign rdata_o[1195] = rdata_i[1195];
  assign rdata_o[1194] = rdata_i[1194];
  assign rdata_o[1193] = rdata_i[1193];
  assign rdata_o[1192] = rdata_i[1192];
  assign rdata_o[1191] = rdata_i[1191];
  assign rdata_o[1190] = rdata_i[1190];
  assign rdata_o[1189] = rdata_i[1189];
  assign rdata_o[1188] = rdata_i[1188];
  assign rdata_o[1187] = rdata_i[1187];
  assign rdata_o[1186] = rdata_i[1186];
  assign rdata_o[1185] = rdata_i[1185];
  assign rdata_o[1184] = rdata_i[1184];
  assign rdata_o[1183] = rdata_i[1183];
  assign rdata_o[1182] = rdata_i[1182];
  assign rdata_o[1181] = rdata_i[1181];
  assign rdata_o[1180] = rdata_i[1180];
  assign rdata_o[1179] = rdata_i[1179];
  assign rdata_o[1178] = rdata_i[1178];
  assign rdata_o[1177] = rdata_i[1177];
  assign rdata_o[1176] = rdata_i[1176];
  assign rdata_o[1175] = rdata_i[1175];
  assign rdata_o[1174] = rdata_i[1174];
  assign rdata_o[1173] = rdata_i[1173];
  assign rdata_o[1172] = rdata_i[1172];
  assign rdata_o[1171] = rdata_i[1171];
  assign rdata_o[1170] = rdata_i[1170];
  assign rdata_o[1169] = rdata_i[1169];
  assign rdata_o[1168] = rdata_i[1168];
  assign rdata_o[1167] = rdata_i[1167];
  assign rdata_o[1166] = rdata_i[1166];
  assign rdata_o[1165] = rdata_i[1165];
  assign rdata_o[1164] = rdata_i[1164];
  assign rdata_o[1163] = rdata_i[1163];
  assign rdata_o[1162] = rdata_i[1162];
  assign rdata_o[1161] = rdata_i[1161];
  assign rdata_o[1160] = rdata_i[1160];
  assign rdata_o[1159] = rdata_i[1159];
  assign rdata_o[1158] = rdata_i[1158];
  assign rdata_o[1157] = rdata_i[1157];
  assign rdata_o[1156] = rdata_i[1156];
  assign rdata_o[1155] = rdata_i[1155];
  assign rdata_o[1154] = rdata_i[1154];
  assign rdata_o[1153] = rdata_i[1153];
  assign rdata_o[1152] = rdata_i[1152];
  assign rdata_o[1151] = rdata_i[1151];
  assign rdata_o[1150] = rdata_i[1150];
  assign rdata_o[1149] = rdata_i[1149];
  assign rdata_o[1148] = rdata_i[1148];
  assign rdata_o[1147] = rdata_i[1147];
  assign rdata_o[1146] = rdata_i[1146];
  assign rdata_o[1145] = rdata_i[1145];
  assign rdata_o[1144] = rdata_i[1144];
  assign rdata_o[1143] = rdata_i[1143];
  assign rdata_o[1142] = rdata_i[1142];
  assign rdata_o[1141] = rdata_i[1141];
  assign rdata_o[1140] = rdata_i[1140];
  assign rdata_o[1139] = rdata_i[1139];
  assign rdata_o[1138] = rdata_i[1138];
  assign rdata_o[1137] = rdata_i[1137];
  assign rdata_o[1136] = rdata_i[1136];
  assign rdata_o[1135] = rdata_i[1135];
  assign rdata_o[1134] = rdata_i[1134];
  assign rdata_o[1133] = rdata_i[1133];
  assign rdata_o[1132] = rdata_i[1132];
  assign rdata_o[1131] = rdata_i[1131];
  assign rdata_o[1130] = rdata_i[1130];
  assign rdata_o[1129] = rdata_i[1129];
  assign rdata_o[1128] = rdata_i[1128];
  assign rdata_o[1127] = rdata_i[1127];
  assign rdata_o[1126] = rdata_i[1126];
  assign rdata_o[1125] = rdata_i[1125];
  assign rdata_o[1124] = rdata_i[1124];
  assign rdata_o[1123] = rdata_i[1123];
  assign rdata_o[1122] = rdata_i[1122];
  assign rdata_o[1121] = rdata_i[1121];
  assign rdata_o[1120] = rdata_i[1120];
  assign rdata_o[1119] = rdata_i[1119];
  assign rdata_o[1118] = rdata_i[1118];
  assign rdata_o[1117] = rdata_i[1117];
  assign rdata_o[1116] = rdata_i[1116];
  assign rdata_o[1115] = rdata_i[1115];
  assign rdata_o[1114] = rdata_i[1114];
  assign rdata_o[1113] = rdata_i[1113];
  assign rdata_o[1112] = rdata_i[1112];
  assign rdata_o[1111] = rdata_i[1111];
  assign rdata_o[1110] = rdata_i[1110];
  assign rdata_o[1109] = rdata_i[1109];
  assign rdata_o[1108] = rdata_i[1108];
  assign rdata_o[1107] = rdata_i[1107];
  assign rdata_o[1106] = rdata_i[1106];
  assign rdata_o[1105] = rdata_i[1105];
  assign rdata_o[1104] = rdata_i[1104];
  assign rdata_o[1103] = rdata_i[1103];
  assign rdata_o[1102] = rdata_i[1102];
  assign rdata_o[1101] = rdata_i[1101];
  assign rdata_o[1100] = rdata_i[1100];
  assign rdata_o[1099] = rdata_i[1099];
  assign rdata_o[1098] = rdata_i[1098];
  assign rdata_o[1097] = rdata_i[1097];
  assign rdata_o[1096] = rdata_i[1096];
  assign rdata_o[1095] = rdata_i[1095];
  assign rdata_o[1094] = rdata_i[1094];
  assign rdata_o[1093] = rdata_i[1093];
  assign rdata_o[1092] = rdata_i[1092];
  assign rdata_o[1091] = rdata_i[1091];
  assign rdata_o[1090] = rdata_i[1090];
  assign rdata_o[1089] = rdata_i[1089];
  assign rdata_o[1088] = rdata_i[1088];
  assign rdata_o[1087] = rdata_i[1087];
  assign rdata_o[1086] = rdata_i[1086];
  assign rdata_o[1085] = rdata_i[1085];
  assign rdata_o[1084] = rdata_i[1084];
  assign rdata_o[1083] = rdata_i[1083];
  assign rdata_o[1082] = rdata_i[1082];
  assign rdata_o[1081] = rdata_i[1081];
  assign rdata_o[1080] = rdata_i[1080];
  assign rdata_o[1079] = rdata_i[1079];
  assign rdata_o[1078] = rdata_i[1078];
  assign rdata_o[1077] = rdata_i[1077];
  assign rdata_o[1076] = rdata_i[1076];
  assign rdata_o[1075] = rdata_i[1075];
  assign rdata_o[1074] = rdata_i[1074];
  assign rdata_o[1073] = rdata_i[1073];
  assign rdata_o[1072] = rdata_i[1072];
  assign rdata_o[1071] = rdata_i[1071];
  assign rdata_o[1070] = rdata_i[1070];
  assign rdata_o[1069] = rdata_i[1069];
  assign rdata_o[1068] = rdata_i[1068];
  assign rdata_o[1067] = rdata_i[1067];
  assign rdata_o[1066] = rdata_i[1066];
  assign rdata_o[1065] = rdata_i[1065];
  assign rdata_o[1064] = rdata_i[1064];
  assign rdata_o[1063] = rdata_i[1063];
  assign rdata_o[1062] = rdata_i[1062];
  assign rdata_o[1061] = rdata_i[1061];
  assign rdata_o[1060] = rdata_i[1060];
  assign rdata_o[1059] = rdata_i[1059];
  assign rdata_o[1058] = rdata_i[1058];
  assign rdata_o[1057] = rdata_i[1057];
  assign rdata_o[1056] = rdata_i[1056];
  assign rdata_o[1055] = rdata_i[1055];
  assign rdata_o[1054] = rdata_i[1054];
  assign rdata_o[1053] = rdata_i[1053];
  assign rdata_o[1052] = rdata_i[1052];
  assign rdata_o[1051] = rdata_i[1051];
  assign rdata_o[1050] = rdata_i[1050];
  assign rdata_o[1049] = rdata_i[1049];
  assign rdata_o[1048] = rdata_i[1048];
  assign rdata_o[1047] = rdata_i[1047];
  assign rdata_o[1046] = rdata_i[1046];
  assign rdata_o[1045] = rdata_i[1045];
  assign rdata_o[1044] = rdata_i[1044];
  assign rdata_o[1043] = rdata_i[1043];
  assign rdata_o[1042] = rdata_i[1042];
  assign rdata_o[1041] = rdata_i[1041];
  assign rdata_o[1040] = rdata_i[1040];
  assign rdata_o[1039] = rdata_i[1039];
  assign rdata_o[1038] = rdata_i[1038];
  assign rdata_o[1037] = rdata_i[1037];
  assign rdata_o[1036] = rdata_i[1036];
  assign rdata_o[1035] = rdata_i[1035];
  assign rdata_o[1034] = rdata_i[1034];
  assign rdata_o[1033] = rdata_i[1033];
  assign rdata_o[1032] = rdata_i[1032];
  assign rdata_o[1031] = rdata_i[1031];
  assign rdata_o[1030] = rdata_i[1030];
  assign rdata_o[1029] = rdata_i[1029];
  assign rdata_o[1028] = rdata_i[1028];
  assign rdata_o[1027] = rdata_i[1027];
  assign rdata_o[1026] = rdata_i[1026];
  assign rdata_o[1025] = rdata_i[1025];
  assign rdata_o[1024] = rdata_i[1024];
  assign rdata_o[1023] = rdata_i[1023];
  assign rdata_o[1022] = rdata_i[1022];
  assign rdata_o[1021] = rdata_i[1021];
  assign rdata_o[1020] = rdata_i[1020];
  assign rdata_o[1019] = rdata_i[1019];
  assign rdata_o[1018] = rdata_i[1018];
  assign rdata_o[1017] = rdata_i[1017];
  assign rdata_o[1016] = rdata_i[1016];
  assign rdata_o[1015] = rdata_i[1015];
  assign rdata_o[1014] = rdata_i[1014];
  assign rdata_o[1013] = rdata_i[1013];
  assign rdata_o[1012] = rdata_i[1012];
  assign rdata_o[1011] = rdata_i[1011];
  assign rdata_o[1010] = rdata_i[1010];
  assign rdata_o[1009] = rdata_i[1009];
  assign rdata_o[1008] = rdata_i[1008];
  assign rdata_o[1007] = rdata_i[1007];
  assign rdata_o[1006] = rdata_i[1006];
  assign rdata_o[1005] = rdata_i[1005];
  assign rdata_o[1004] = rdata_i[1004];
  assign rdata_o[1003] = rdata_i[1003];
  assign rdata_o[1002] = rdata_i[1002];
  assign rdata_o[1001] = rdata_i[1001];
  assign rdata_o[1000] = rdata_i[1000];
  assign rdata_o[999] = rdata_i[999];
  assign rdata_o[998] = rdata_i[998];
  assign rdata_o[997] = rdata_i[997];
  assign rdata_o[996] = rdata_i[996];
  assign rdata_o[995] = rdata_i[995];
  assign rdata_o[994] = rdata_i[994];
  assign rdata_o[993] = rdata_i[993];
  assign rdata_o[992] = rdata_i[992];
  assign rdata_o[991] = rdata_i[991];
  assign rdata_o[990] = rdata_i[990];
  assign rdata_o[989] = rdata_i[989];
  assign rdata_o[988] = rdata_i[988];
  assign rdata_o[987] = rdata_i[987];
  assign rdata_o[986] = rdata_i[986];
  assign rdata_o[985] = rdata_i[985];
  assign rdata_o[984] = rdata_i[984];
  assign rdata_o[983] = rdata_i[983];
  assign rdata_o[982] = rdata_i[982];
  assign rdata_o[981] = rdata_i[981];
  assign rdata_o[980] = rdata_i[980];
  assign rdata_o[979] = rdata_i[979];
  assign rdata_o[978] = rdata_i[978];
  assign rdata_o[977] = rdata_i[977];
  assign rdata_o[976] = rdata_i[976];
  assign rdata_o[975] = rdata_i[975];
  assign rdata_o[974] = rdata_i[974];
  assign rdata_o[973] = rdata_i[973];
  assign rdata_o[972] = rdata_i[972];
  assign rdata_o[971] = rdata_i[971];
  assign rdata_o[970] = rdata_i[970];
  assign rdata_o[969] = rdata_i[969];
  assign rdata_o[968] = rdata_i[968];
  assign rdata_o[967] = rdata_i[967];
  assign rdata_o[966] = rdata_i[966];
  assign rdata_o[965] = rdata_i[965];
  assign rdata_o[964] = rdata_i[964];
  assign rdata_o[963] = rdata_i[963];
  assign rdata_o[962] = rdata_i[962];
  assign rdata_o[961] = rdata_i[961];
  assign rdata_o[960] = rdata_i[960];
  assign rdata_o[959] = rdata_i[959];
  assign rdata_o[958] = rdata_i[958];
  assign rdata_o[957] = rdata_i[957];
  assign rdata_o[956] = rdata_i[956];
  assign rdata_o[955] = rdata_i[955];
  assign rdata_o[954] = rdata_i[954];
  assign rdata_o[953] = rdata_i[953];
  assign rdata_o[952] = rdata_i[952];
  assign rdata_o[951] = rdata_i[951];
  assign rdata_o[950] = rdata_i[950];
  assign rdata_o[949] = rdata_i[949];
  assign rdata_o[948] = rdata_i[948];
  assign rdata_o[947] = rdata_i[947];
  assign rdata_o[946] = rdata_i[946];
  assign rdata_o[945] = rdata_i[945];
  assign rdata_o[944] = rdata_i[944];
  assign rdata_o[943] = rdata_i[943];
  assign rdata_o[942] = rdata_i[942];
  assign rdata_o[941] = rdata_i[941];
  assign rdata_o[940] = rdata_i[940];
  assign rdata_o[939] = rdata_i[939];
  assign rdata_o[938] = rdata_i[938];
  assign rdata_o[937] = rdata_i[937];
  assign rdata_o[936] = rdata_i[936];
  assign rdata_o[935] = rdata_i[935];
  assign rdata_o[934] = rdata_i[934];
  assign rdata_o[933] = rdata_i[933];
  assign rdata_o[932] = rdata_i[932];
  assign rdata_o[931] = rdata_i[931];
  assign rdata_o[930] = rdata_i[930];
  assign rdata_o[929] = rdata_i[929];
  assign rdata_o[928] = rdata_i[928];
  assign rdata_o[927] = rdata_i[927];
  assign rdata_o[926] = rdata_i[926];
  assign rdata_o[925] = rdata_i[925];
  assign rdata_o[924] = rdata_i[924];
  assign rdata_o[923] = rdata_i[923];
  assign rdata_o[922] = rdata_i[922];
  assign rdata_o[921] = rdata_i[921];
  assign rdata_o[920] = rdata_i[920];
  assign rdata_o[919] = rdata_i[919];
  assign rdata_o[918] = rdata_i[918];
  assign rdata_o[917] = rdata_i[917];
  assign rdata_o[916] = rdata_i[916];
  assign rdata_o[915] = rdata_i[915];
  assign rdata_o[914] = rdata_i[914];
  assign rdata_o[913] = rdata_i[913];
  assign rdata_o[912] = rdata_i[912];
  assign rdata_o[911] = rdata_i[911];
  assign rdata_o[910] = rdata_i[910];
  assign rdata_o[909] = rdata_i[909];
  assign rdata_o[908] = rdata_i[908];
  assign rdata_o[907] = rdata_i[907];
  assign rdata_o[906] = rdata_i[906];
  assign rdata_o[905] = rdata_i[905];
  assign rdata_o[904] = rdata_i[904];
  assign rdata_o[903] = rdata_i[903];
  assign rdata_o[902] = rdata_i[902];
  assign rdata_o[901] = rdata_i[901];
  assign rdata_o[900] = rdata_i[900];
  assign rdata_o[899] = rdata_i[899];
  assign rdata_o[898] = rdata_i[898];
  assign rdata_o[897] = rdata_i[897];
  assign rdata_o[896] = rdata_i[896];
  assign rdata_o[895] = rdata_i[895];
  assign rdata_o[894] = rdata_i[894];
  assign rdata_o[893] = rdata_i[893];
  assign rdata_o[892] = rdata_i[892];
  assign rdata_o[891] = rdata_i[891];
  assign rdata_o[890] = rdata_i[890];
  assign rdata_o[889] = rdata_i[889];
  assign rdata_o[888] = rdata_i[888];
  assign rdata_o[887] = rdata_i[887];
  assign rdata_o[886] = rdata_i[886];
  assign rdata_o[885] = rdata_i[885];
  assign rdata_o[884] = rdata_i[884];
  assign rdata_o[883] = rdata_i[883];
  assign rdata_o[882] = rdata_i[882];
  assign rdata_o[881] = rdata_i[881];
  assign rdata_o[880] = rdata_i[880];
  assign rdata_o[879] = rdata_i[879];
  assign rdata_o[878] = rdata_i[878];
  assign rdata_o[877] = rdata_i[877];
  assign rdata_o[876] = rdata_i[876];
  assign rdata_o[875] = rdata_i[875];
  assign rdata_o[874] = rdata_i[874];
  assign rdata_o[873] = rdata_i[873];
  assign rdata_o[872] = rdata_i[872];
  assign rdata_o[871] = rdata_i[871];
  assign rdata_o[870] = rdata_i[870];
  assign rdata_o[869] = rdata_i[869];
  assign rdata_o[868] = rdata_i[868];
  assign rdata_o[867] = rdata_i[867];
  assign rdata_o[866] = rdata_i[866];
  assign rdata_o[865] = rdata_i[865];
  assign rdata_o[864] = rdata_i[864];
  assign rdata_o[863] = rdata_i[863];
  assign rdata_o[862] = rdata_i[862];
  assign rdata_o[861] = rdata_i[861];
  assign rdata_o[860] = rdata_i[860];
  assign rdata_o[859] = rdata_i[859];
  assign rdata_o[858] = rdata_i[858];
  assign rdata_o[857] = rdata_i[857];
  assign rdata_o[856] = rdata_i[856];
  assign rdata_o[855] = rdata_i[855];
  assign rdata_o[854] = rdata_i[854];
  assign rdata_o[853] = rdata_i[853];
  assign rdata_o[852] = rdata_i[852];
  assign rdata_o[851] = rdata_i[851];
  assign rdata_o[850] = rdata_i[850];
  assign rdata_o[849] = rdata_i[849];
  assign rdata_o[848] = rdata_i[848];
  assign rdata_o[847] = rdata_i[847];
  assign rdata_o[846] = rdata_i[846];
  assign rdata_o[845] = rdata_i[845];
  assign rdata_o[844] = rdata_i[844];
  assign rdata_o[843] = rdata_i[843];
  assign rdata_o[842] = rdata_i[842];
  assign rdata_o[841] = rdata_i[841];
  assign rdata_o[840] = rdata_i[840];
  assign rdata_o[839] = rdata_i[839];
  assign rdata_o[838] = rdata_i[838];
  assign rdata_o[837] = rdata_i[837];
  assign rdata_o[836] = rdata_i[836];
  assign rdata_o[835] = rdata_i[835];
  assign rdata_o[834] = rdata_i[834];
  assign rdata_o[833] = rdata_i[833];
  assign rdata_o[832] = rdata_i[832];
  assign rdata_o[831] = rdata_i[831];
  assign rdata_o[830] = rdata_i[830];
  assign rdata_o[829] = rdata_i[829];
  assign rdata_o[828] = rdata_i[828];
  assign rdata_o[827] = rdata_i[827];
  assign rdata_o[826] = rdata_i[826];
  assign rdata_o[825] = rdata_i[825];
  assign rdata_o[824] = rdata_i[824];
  assign rdata_o[823] = rdata_i[823];
  assign rdata_o[822] = rdata_i[822];
  assign rdata_o[821] = rdata_i[821];
  assign rdata_o[820] = rdata_i[820];
  assign rdata_o[819] = rdata_i[819];
  assign rdata_o[818] = rdata_i[818];
  assign rdata_o[817] = rdata_i[817];
  assign rdata_o[816] = rdata_i[816];
  assign rdata_o[815] = rdata_i[815];
  assign rdata_o[814] = rdata_i[814];
  assign rdata_o[813] = rdata_i[813];
  assign rdata_o[812] = rdata_i[812];
  assign rdata_o[811] = rdata_i[811];
  assign rdata_o[810] = rdata_i[810];
  assign rdata_o[809] = rdata_i[809];
  assign rdata_o[808] = rdata_i[808];
  assign rdata_o[807] = rdata_i[807];
  assign rdata_o[806] = rdata_i[806];
  assign rdata_o[805] = rdata_i[805];
  assign rdata_o[804] = rdata_i[804];
  assign rdata_o[803] = rdata_i[803];
  assign rdata_o[802] = rdata_i[802];
  assign rdata_o[801] = rdata_i[801];
  assign rdata_o[800] = rdata_i[800];
  assign rdata_o[799] = rdata_i[799];
  assign rdata_o[798] = rdata_i[798];
  assign rdata_o[797] = rdata_i[797];
  assign rdata_o[796] = rdata_i[796];
  assign rdata_o[795] = rdata_i[795];
  assign rdata_o[794] = rdata_i[794];
  assign rdata_o[793] = rdata_i[793];
  assign rdata_o[792] = rdata_i[792];
  assign rdata_o[791] = rdata_i[791];
  assign rdata_o[790] = rdata_i[790];
  assign rdata_o[789] = rdata_i[789];
  assign rdata_o[788] = rdata_i[788];
  assign rdata_o[787] = rdata_i[787];
  assign rdata_o[786] = rdata_i[786];
  assign rdata_o[785] = rdata_i[785];
  assign rdata_o[784] = rdata_i[784];
  assign rdata_o[783] = rdata_i[783];
  assign rdata_o[782] = rdata_i[782];
  assign rdata_o[781] = rdata_i[781];
  assign rdata_o[780] = rdata_i[780];
  assign rdata_o[779] = rdata_i[779];
  assign rdata_o[778] = rdata_i[778];
  assign rdata_o[777] = rdata_i[777];
  assign rdata_o[776] = rdata_i[776];
  assign rdata_o[775] = rdata_i[775];
  assign rdata_o[774] = rdata_i[774];
  assign rdata_o[773] = rdata_i[773];
  assign rdata_o[772] = rdata_i[772];
  assign rdata_o[771] = rdata_i[771];
  assign rdata_o[770] = rdata_i[770];
  assign rdata_o[769] = rdata_i[769];
  assign rdata_o[768] = rdata_i[768];
  assign rdata_o[767] = rdata_i[767];
  assign rdata_o[766] = rdata_i[766];
  assign rdata_o[765] = rdata_i[765];
  assign rdata_o[764] = rdata_i[764];
  assign rdata_o[763] = rdata_i[763];
  assign rdata_o[762] = rdata_i[762];
  assign rdata_o[761] = rdata_i[761];
  assign rdata_o[760] = rdata_i[760];
  assign rdata_o[759] = rdata_i[759];
  assign rdata_o[758] = rdata_i[758];
  assign rdata_o[757] = rdata_i[757];
  assign rdata_o[756] = rdata_i[756];
  assign rdata_o[755] = rdata_i[755];
  assign rdata_o[754] = rdata_i[754];
  assign rdata_o[753] = rdata_i[753];
  assign rdata_o[752] = rdata_i[752];
  assign rdata_o[751] = rdata_i[751];
  assign rdata_o[750] = rdata_i[750];
  assign rdata_o[749] = rdata_i[749];
  assign rdata_o[748] = rdata_i[748];
  assign rdata_o[747] = rdata_i[747];
  assign rdata_o[746] = rdata_i[746];
  assign rdata_o[745] = rdata_i[745];
  assign rdata_o[744] = rdata_i[744];
  assign rdata_o[743] = rdata_i[743];
  assign rdata_o[742] = rdata_i[742];
  assign rdata_o[741] = rdata_i[741];
  assign rdata_o[740] = rdata_i[740];
  assign rdata_o[739] = rdata_i[739];
  assign rdata_o[738] = rdata_i[738];
  assign rdata_o[737] = rdata_i[737];
  assign rdata_o[736] = rdata_i[736];
  assign rdata_o[735] = rdata_i[735];
  assign rdata_o[734] = rdata_i[734];
  assign rdata_o[733] = rdata_i[733];
  assign rdata_o[732] = rdata_i[732];
  assign rdata_o[731] = rdata_i[731];
  assign rdata_o[730] = rdata_i[730];
  assign rdata_o[729] = rdata_i[729];
  assign rdata_o[728] = rdata_i[728];
  assign rdata_o[727] = rdata_i[727];
  assign rdata_o[726] = rdata_i[726];
  assign rdata_o[725] = rdata_i[725];
  assign rdata_o[724] = rdata_i[724];
  assign rdata_o[723] = rdata_i[723];
  assign rdata_o[722] = rdata_i[722];
  assign rdata_o[721] = rdata_i[721];
  assign rdata_o[720] = rdata_i[720];
  assign rdata_o[719] = rdata_i[719];
  assign rdata_o[718] = rdata_i[718];
  assign rdata_o[717] = rdata_i[717];
  assign rdata_o[716] = rdata_i[716];
  assign rdata_o[715] = rdata_i[715];
  assign rdata_o[714] = rdata_i[714];
  assign rdata_o[713] = rdata_i[713];
  assign rdata_o[712] = rdata_i[712];
  assign rdata_o[711] = rdata_i[711];
  assign rdata_o[710] = rdata_i[710];
  assign rdata_o[709] = rdata_i[709];
  assign rdata_o[708] = rdata_i[708];
  assign rdata_o[707] = rdata_i[707];
  assign rdata_o[706] = rdata_i[706];
  assign rdata_o[705] = rdata_i[705];
  assign rdata_o[704] = rdata_i[704];
  assign rdata_o[703] = rdata_i[703];
  assign rdata_o[702] = rdata_i[702];
  assign rdata_o[701] = rdata_i[701];
  assign rdata_o[700] = rdata_i[700];
  assign rdata_o[699] = rdata_i[699];
  assign rdata_o[698] = rdata_i[698];
  assign rdata_o[697] = rdata_i[697];
  assign rdata_o[696] = rdata_i[696];
  assign rdata_o[695] = rdata_i[695];
  assign rdata_o[694] = rdata_i[694];
  assign rdata_o[693] = rdata_i[693];
  assign rdata_o[692] = rdata_i[692];
  assign rdata_o[691] = rdata_i[691];
  assign rdata_o[690] = rdata_i[690];
  assign rdata_o[689] = rdata_i[689];
  assign rdata_o[688] = rdata_i[688];
  assign rdata_o[687] = rdata_i[687];
  assign rdata_o[686] = rdata_i[686];
  assign rdata_o[685] = rdata_i[685];
  assign rdata_o[684] = rdata_i[684];
  assign rdata_o[683] = rdata_i[683];
  assign rdata_o[682] = rdata_i[682];
  assign rdata_o[681] = rdata_i[681];
  assign rdata_o[680] = rdata_i[680];
  assign rdata_o[679] = rdata_i[679];
  assign rdata_o[678] = rdata_i[678];
  assign rdata_o[677] = rdata_i[677];
  assign rdata_o[676] = rdata_i[676];
  assign rdata_o[675] = rdata_i[675];
  assign rdata_o[674] = rdata_i[674];
  assign rdata_o[673] = rdata_i[673];
  assign rdata_o[672] = rdata_i[672];
  assign rdata_o[671] = rdata_i[671];
  assign rdata_o[670] = rdata_i[670];
  assign rdata_o[669] = rdata_i[669];
  assign rdata_o[668] = rdata_i[668];
  assign rdata_o[667] = rdata_i[667];
  assign rdata_o[666] = rdata_i[666];
  assign rdata_o[665] = rdata_i[665];
  assign rdata_o[664] = rdata_i[664];
  assign rdata_o[663] = rdata_i[663];
  assign rdata_o[662] = rdata_i[662];
  assign rdata_o[661] = rdata_i[661];
  assign rdata_o[660] = rdata_i[660];
  assign rdata_o[659] = rdata_i[659];
  assign rdata_o[658] = rdata_i[658];
  assign rdata_o[657] = rdata_i[657];
  assign rdata_o[656] = rdata_i[656];
  assign rdata_o[655] = rdata_i[655];
  assign rdata_o[654] = rdata_i[654];
  assign rdata_o[653] = rdata_i[653];
  assign rdata_o[652] = rdata_i[652];
  assign rdata_o[651] = rdata_i[651];
  assign rdata_o[650] = rdata_i[650];
  assign rdata_o[649] = rdata_i[649];
  assign rdata_o[648] = rdata_i[648];
  assign rdata_o[647] = rdata_i[647];
  assign rdata_o[646] = rdata_i[646];
  assign rdata_o[645] = rdata_i[645];
  assign rdata_o[644] = rdata_i[644];
  assign rdata_o[643] = rdata_i[643];
  assign rdata_o[642] = rdata_i[642];
  assign rdata_o[641] = rdata_i[641];
  assign rdata_o[640] = rdata_i[640];
  assign rdata_o[639] = rdata_i[639];
  assign rdata_o[638] = rdata_i[638];
  assign rdata_o[637] = rdata_i[637];
  assign rdata_o[636] = rdata_i[636];
  assign rdata_o[635] = rdata_i[635];
  assign rdata_o[634] = rdata_i[634];
  assign rdata_o[633] = rdata_i[633];
  assign rdata_o[632] = rdata_i[632];
  assign rdata_o[631] = rdata_i[631];
  assign rdata_o[630] = rdata_i[630];
  assign rdata_o[629] = rdata_i[629];
  assign rdata_o[628] = rdata_i[628];
  assign rdata_o[627] = rdata_i[627];
  assign rdata_o[626] = rdata_i[626];
  assign rdata_o[625] = rdata_i[625];
  assign rdata_o[624] = rdata_i[624];
  assign rdata_o[623] = rdata_i[623];
  assign rdata_o[622] = rdata_i[622];
  assign rdata_o[621] = rdata_i[621];
  assign rdata_o[620] = rdata_i[620];
  assign rdata_o[619] = rdata_i[619];
  assign rdata_o[618] = rdata_i[618];
  assign rdata_o[617] = rdata_i[617];
  assign rdata_o[616] = rdata_i[616];
  assign rdata_o[615] = rdata_i[615];
  assign rdata_o[614] = rdata_i[614];
  assign rdata_o[613] = rdata_i[613];
  assign rdata_o[612] = rdata_i[612];
  assign rdata_o[611] = rdata_i[611];
  assign rdata_o[610] = rdata_i[610];
  assign rdata_o[609] = rdata_i[609];
  assign rdata_o[608] = rdata_i[608];
  assign rdata_o[607] = rdata_i[607];
  assign rdata_o[606] = rdata_i[606];
  assign rdata_o[605] = rdata_i[605];
  assign rdata_o[604] = rdata_i[604];
  assign rdata_o[603] = rdata_i[603];
  assign rdata_o[602] = rdata_i[602];
  assign rdata_o[601] = rdata_i[601];
  assign rdata_o[600] = rdata_i[600];
  assign rdata_o[599] = rdata_i[599];
  assign rdata_o[598] = rdata_i[598];
  assign rdata_o[597] = rdata_i[597];
  assign rdata_o[596] = rdata_i[596];
  assign rdata_o[595] = rdata_i[595];
  assign rdata_o[594] = rdata_i[594];
  assign rdata_o[593] = rdata_i[593];
  assign rdata_o[592] = rdata_i[592];
  assign rdata_o[591] = rdata_i[591];
  assign rdata_o[590] = rdata_i[590];
  assign rdata_o[589] = rdata_i[589];
  assign rdata_o[588] = rdata_i[588];
  assign rdata_o[587] = rdata_i[587];
  assign rdata_o[586] = rdata_i[586];
  assign rdata_o[585] = rdata_i[585];
  assign rdata_o[584] = rdata_i[584];
  assign rdata_o[583] = rdata_i[583];
  assign rdata_o[582] = rdata_i[582];
  assign rdata_o[581] = rdata_i[581];
  assign rdata_o[580] = rdata_i[580];
  assign rdata_o[579] = rdata_i[579];
  assign rdata_o[578] = rdata_i[578];
  assign rdata_o[577] = rdata_i[577];
  assign rdata_o[576] = rdata_i[576];
  assign rdata_o[575] = rdata_i[575];
  assign rdata_o[574] = rdata_i[574];
  assign rdata_o[573] = rdata_i[573];
  assign rdata_o[572] = rdata_i[572];
  assign rdata_o[571] = rdata_i[571];
  assign rdata_o[570] = rdata_i[570];
  assign rdata_o[569] = rdata_i[569];
  assign rdata_o[568] = rdata_i[568];
  assign rdata_o[567] = rdata_i[567];
  assign rdata_o[566] = rdata_i[566];
  assign rdata_o[565] = rdata_i[565];
  assign rdata_o[564] = rdata_i[564];
  assign rdata_o[563] = rdata_i[563];
  assign rdata_o[562] = rdata_i[562];
  assign rdata_o[561] = rdata_i[561];
  assign rdata_o[560] = rdata_i[560];
  assign rdata_o[559] = rdata_i[559];
  assign rdata_o[558] = rdata_i[558];
  assign rdata_o[557] = rdata_i[557];
  assign rdata_o[556] = rdata_i[556];
  assign rdata_o[555] = rdata_i[555];
  assign rdata_o[554] = rdata_i[554];
  assign rdata_o[553] = rdata_i[553];
  assign rdata_o[552] = rdata_i[552];
  assign rdata_o[551] = rdata_i[551];
  assign rdata_o[550] = rdata_i[550];
  assign rdata_o[549] = rdata_i[549];
  assign rdata_o[548] = rdata_i[548];
  assign rdata_o[547] = rdata_i[547];
  assign rdata_o[546] = rdata_i[546];
  assign rdata_o[545] = rdata_i[545];
  assign rdata_o[544] = rdata_i[544];
  assign rdata_o[543] = rdata_i[543];
  assign rdata_o[542] = rdata_i[542];
  assign rdata_o[541] = rdata_i[541];
  assign rdata_o[540] = rdata_i[540];
  assign rdata_o[539] = rdata_i[539];
  assign rdata_o[538] = rdata_i[538];
  assign rdata_o[537] = rdata_i[537];
  assign rdata_o[536] = rdata_i[536];
  assign rdata_o[535] = rdata_i[535];
  assign rdata_o[534] = rdata_i[534];
  assign rdata_o[533] = rdata_i[533];
  assign rdata_o[532] = rdata_i[532];
  assign rdata_o[531] = rdata_i[531];
  assign rdata_o[530] = rdata_i[530];
  assign rdata_o[529] = rdata_i[529];
  assign rdata_o[528] = rdata_i[528];
  assign rdata_o[527] = rdata_i[527];
  assign rdata_o[526] = rdata_i[526];
  assign rdata_o[525] = rdata_i[525];
  assign rdata_o[524] = rdata_i[524];
  assign rdata_o[523] = rdata_i[523];
  assign rdata_o[522] = rdata_i[522];
  assign rdata_o[521] = rdata_i[521];
  assign rdata_o[520] = rdata_i[520];
  assign rdata_o[519] = rdata_i[519];
  assign rdata_o[518] = rdata_i[518];
  assign rdata_o[517] = rdata_i[517];
  assign rdata_o[516] = rdata_i[516];
  assign rdata_o[515] = rdata_i[515];
  assign rdata_o[514] = rdata_i[514];
  assign rdata_o[513] = rdata_i[513];
  assign rdata_o[512] = rdata_i[512];
  assign rdata_o[511] = rdata_i[511];
  assign rdata_o[510] = rdata_i[510];
  assign rdata_o[509] = rdata_i[509];
  assign rdata_o[508] = rdata_i[508];
  assign rdata_o[507] = rdata_i[507];
  assign rdata_o[506] = rdata_i[506];
  assign rdata_o[505] = rdata_i[505];
  assign rdata_o[504] = rdata_i[504];
  assign rdata_o[503] = rdata_i[503];
  assign rdata_o[502] = rdata_i[502];
  assign rdata_o[501] = rdata_i[501];
  assign rdata_o[500] = rdata_i[500];
  assign rdata_o[499] = rdata_i[499];
  assign rdata_o[498] = rdata_i[498];
  assign rdata_o[497] = rdata_i[497];
  assign rdata_o[496] = rdata_i[496];
  assign rdata_o[495] = rdata_i[495];
  assign rdata_o[494] = rdata_i[494];
  assign rdata_o[493] = rdata_i[493];
  assign rdata_o[492] = rdata_i[492];
  assign rdata_o[491] = rdata_i[491];
  assign rdata_o[490] = rdata_i[490];
  assign rdata_o[489] = rdata_i[489];
  assign rdata_o[488] = rdata_i[488];
  assign rdata_o[487] = rdata_i[487];
  assign rdata_o[486] = rdata_i[486];
  assign rdata_o[485] = rdata_i[485];
  assign rdata_o[484] = rdata_i[484];
  assign rdata_o[483] = rdata_i[483];
  assign rdata_o[482] = rdata_i[482];
  assign rdata_o[481] = rdata_i[481];
  assign rdata_o[480] = rdata_i[480];
  assign rdata_o[479] = rdata_i[479];
  assign rdata_o[478] = rdata_i[478];
  assign rdata_o[477] = rdata_i[477];
  assign rdata_o[476] = rdata_i[476];
  assign rdata_o[475] = rdata_i[475];
  assign rdata_o[474] = rdata_i[474];
  assign rdata_o[473] = rdata_i[473];
  assign rdata_o[472] = rdata_i[472];
  assign rdata_o[471] = rdata_i[471];
  assign rdata_o[470] = rdata_i[470];
  assign rdata_o[469] = rdata_i[469];
  assign rdata_o[468] = rdata_i[468];
  assign rdata_o[467] = rdata_i[467];
  assign rdata_o[466] = rdata_i[466];
  assign rdata_o[465] = rdata_i[465];
  assign rdata_o[464] = rdata_i[464];
  assign rdata_o[463] = rdata_i[463];
  assign rdata_o[462] = rdata_i[462];
  assign rdata_o[461] = rdata_i[461];
  assign rdata_o[460] = rdata_i[460];
  assign rdata_o[459] = rdata_i[459];
  assign rdata_o[458] = rdata_i[458];
  assign rdata_o[457] = rdata_i[457];
  assign rdata_o[456] = rdata_i[456];
  assign rdata_o[455] = rdata_i[455];
  assign rdata_o[454] = rdata_i[454];
  assign rdata_o[453] = rdata_i[453];
  assign rdata_o[452] = rdata_i[452];
  assign rdata_o[451] = rdata_i[451];
  assign rdata_o[450] = rdata_i[450];
  assign rdata_o[449] = rdata_i[449];
  assign rdata_o[448] = rdata_i[448];
  assign rdata_o[447] = rdata_i[447];
  assign rdata_o[446] = rdata_i[446];
  assign rdata_o[445] = rdata_i[445];
  assign rdata_o[444] = rdata_i[444];
  assign rdata_o[443] = rdata_i[443];
  assign rdata_o[442] = rdata_i[442];
  assign rdata_o[441] = rdata_i[441];
  assign rdata_o[440] = rdata_i[440];
  assign rdata_o[439] = rdata_i[439];
  assign rdata_o[438] = rdata_i[438];
  assign rdata_o[437] = rdata_i[437];
  assign rdata_o[436] = rdata_i[436];
  assign rdata_o[435] = rdata_i[435];
  assign rdata_o[434] = rdata_i[434];
  assign rdata_o[433] = rdata_i[433];
  assign rdata_o[432] = rdata_i[432];
  assign rdata_o[431] = rdata_i[431];
  assign rdata_o[430] = rdata_i[430];
  assign rdata_o[429] = rdata_i[429];
  assign rdata_o[428] = rdata_i[428];
  assign rdata_o[427] = rdata_i[427];
  assign rdata_o[426] = rdata_i[426];
  assign rdata_o[425] = rdata_i[425];
  assign rdata_o[424] = rdata_i[424];
  assign rdata_o[423] = rdata_i[423];
  assign rdata_o[422] = rdata_i[422];
  assign rdata_o[421] = rdata_i[421];
  assign rdata_o[420] = rdata_i[420];
  assign rdata_o[419] = rdata_i[419];
  assign rdata_o[418] = rdata_i[418];
  assign rdata_o[417] = rdata_i[417];
  assign rdata_o[416] = rdata_i[416];
  assign rdata_o[415] = rdata_i[415];
  assign rdata_o[414] = rdata_i[414];
  assign rdata_o[413] = rdata_i[413];
  assign rdata_o[412] = rdata_i[412];
  assign rdata_o[411] = rdata_i[411];
  assign rdata_o[410] = rdata_i[410];
  assign rdata_o[409] = rdata_i[409];
  assign rdata_o[408] = rdata_i[408];
  assign rdata_o[407] = rdata_i[407];
  assign rdata_o[406] = rdata_i[406];
  assign rdata_o[405] = rdata_i[405];
  assign rdata_o[404] = rdata_i[404];
  assign rdata_o[403] = rdata_i[403];
  assign rdata_o[402] = rdata_i[402];
  assign rdata_o[401] = rdata_i[401];
  assign rdata_o[400] = rdata_i[400];
  assign rdata_o[399] = rdata_i[399];
  assign rdata_o[398] = rdata_i[398];
  assign rdata_o[397] = rdata_i[397];
  assign rdata_o[396] = rdata_i[396];
  assign rdata_o[395] = rdata_i[395];
  assign rdata_o[394] = rdata_i[394];
  assign rdata_o[393] = rdata_i[393];
  assign rdata_o[392] = rdata_i[392];
  assign rdata_o[391] = rdata_i[391];
  assign rdata_o[390] = rdata_i[390];
  assign rdata_o[389] = rdata_i[389];
  assign rdata_o[388] = rdata_i[388];
  assign rdata_o[387] = rdata_i[387];
  assign rdata_o[386] = rdata_i[386];
  assign rdata_o[385] = rdata_i[385];
  assign rdata_o[384] = rdata_i[384];
  assign rdata_o[383] = rdata_i[383];
  assign rdata_o[382] = rdata_i[382];
  assign rdata_o[381] = rdata_i[381];
  assign rdata_o[380] = rdata_i[380];
  assign rdata_o[379] = rdata_i[379];
  assign rdata_o[378] = rdata_i[378];
  assign rdata_o[377] = rdata_i[377];
  assign rdata_o[376] = rdata_i[376];
  assign rdata_o[375] = rdata_i[375];
  assign rdata_o[374] = rdata_i[374];
  assign rdata_o[373] = rdata_i[373];
  assign rdata_o[372] = rdata_i[372];
  assign rdata_o[371] = rdata_i[371];
  assign rdata_o[370] = rdata_i[370];
  assign rdata_o[369] = rdata_i[369];
  assign rdata_o[368] = rdata_i[368];
  assign rdata_o[367] = rdata_i[367];
  assign rdata_o[366] = rdata_i[366];
  assign rdata_o[365] = rdata_i[365];
  assign rdata_o[364] = rdata_i[364];
  assign rdata_o[363] = rdata_i[363];
  assign rdata_o[362] = rdata_i[362];
  assign rdata_o[361] = rdata_i[361];
  assign rdata_o[360] = rdata_i[360];
  assign rdata_o[359] = rdata_i[359];
  assign rdata_o[358] = rdata_i[358];
  assign rdata_o[357] = rdata_i[357];
  assign rdata_o[356] = rdata_i[356];
  assign rdata_o[355] = rdata_i[355];
  assign rdata_o[354] = rdata_i[354];
  assign rdata_o[353] = rdata_i[353];
  assign rdata_o[352] = rdata_i[352];
  assign rdata_o[351] = rdata_i[351];
  assign rdata_o[350] = rdata_i[350];
  assign rdata_o[349] = rdata_i[349];
  assign rdata_o[348] = rdata_i[348];
  assign rdata_o[347] = rdata_i[347];
  assign rdata_o[346] = rdata_i[346];
  assign rdata_o[345] = rdata_i[345];
  assign rdata_o[344] = rdata_i[344];
  assign rdata_o[343] = rdata_i[343];
  assign rdata_o[342] = rdata_i[342];
  assign rdata_o[341] = rdata_i[341];
  assign rdata_o[340] = rdata_i[340];
  assign rdata_o[339] = rdata_i[339];
  assign rdata_o[338] = rdata_i[338];
  assign rdata_o[337] = rdata_i[337];
  assign rdata_o[336] = rdata_i[336];
  assign rdata_o[335] = rdata_i[335];
  assign rdata_o[334] = rdata_i[334];
  assign rdata_o[333] = rdata_i[333];
  assign rdata_o[332] = rdata_i[332];
  assign rdata_o[331] = rdata_i[331];
  assign rdata_o[330] = rdata_i[330];
  assign rdata_o[329] = rdata_i[329];
  assign rdata_o[328] = rdata_i[328];
  assign rdata_o[327] = rdata_i[327];
  assign rdata_o[326] = rdata_i[326];
  assign rdata_o[325] = rdata_i[325];
  assign rdata_o[324] = rdata_i[324];
  assign rdata_o[323] = rdata_i[323];
  assign rdata_o[322] = rdata_i[322];
  assign rdata_o[321] = rdata_i[321];
  assign rdata_o[320] = rdata_i[320];
  assign rdata_o[319] = rdata_i[319];
  assign rdata_o[318] = rdata_i[318];
  assign rdata_o[317] = rdata_i[317];
  assign rdata_o[316] = rdata_i[316];
  assign rdata_o[315] = rdata_i[315];
  assign rdata_o[314] = rdata_i[314];
  assign rdata_o[313] = rdata_i[313];
  assign rdata_o[312] = rdata_i[312];
  assign rdata_o[311] = rdata_i[311];
  assign rdata_o[310] = rdata_i[310];
  assign rdata_o[309] = rdata_i[309];
  assign rdata_o[308] = rdata_i[308];
  assign rdata_o[307] = rdata_i[307];
  assign rdata_o[306] = rdata_i[306];
  assign rdata_o[305] = rdata_i[305];
  assign rdata_o[304] = rdata_i[304];
  assign rdata_o[303] = rdata_i[303];
  assign rdata_o[302] = rdata_i[302];
  assign rdata_o[301] = rdata_i[301];
  assign rdata_o[300] = rdata_i[300];
  assign rdata_o[299] = rdata_i[299];
  assign rdata_o[298] = rdata_i[298];
  assign rdata_o[297] = rdata_i[297];
  assign rdata_o[296] = rdata_i[296];
  assign rdata_o[295] = rdata_i[295];
  assign rdata_o[294] = rdata_i[294];
  assign rdata_o[293] = rdata_i[293];
  assign rdata_o[292] = rdata_i[292];
  assign rdata_o[291] = rdata_i[291];
  assign rdata_o[290] = rdata_i[290];
  assign rdata_o[289] = rdata_i[289];
  assign rdata_o[288] = rdata_i[288];
  assign rdata_o[287] = rdata_i[287];
  assign rdata_o[286] = rdata_i[286];
  assign rdata_o[285] = rdata_i[285];
  assign rdata_o[284] = rdata_i[284];
  assign rdata_o[283] = rdata_i[283];
  assign rdata_o[282] = rdata_i[282];
  assign rdata_o[281] = rdata_i[281];
  assign rdata_o[280] = rdata_i[280];
  assign rdata_o[279] = rdata_i[279];
  assign rdata_o[278] = rdata_i[278];
  assign rdata_o[277] = rdata_i[277];
  assign rdata_o[276] = rdata_i[276];
  assign rdata_o[275] = rdata_i[275];
  assign rdata_o[274] = rdata_i[274];
  assign rdata_o[273] = rdata_i[273];
  assign rdata_o[272] = rdata_i[272];
  assign rdata_o[271] = rdata_i[271];
  assign rdata_o[270] = rdata_i[270];
  assign rdata_o[269] = rdata_i[269];
  assign rdata_o[268] = rdata_i[268];
  assign rdata_o[267] = rdata_i[267];
  assign rdata_o[266] = rdata_i[266];
  assign rdata_o[265] = rdata_i[265];
  assign rdata_o[264] = rdata_i[264];
  assign rdata_o[263] = rdata_i[263];
  assign rdata_o[262] = rdata_i[262];
  assign rdata_o[261] = rdata_i[261];
  assign rdata_o[260] = rdata_i[260];
  assign rdata_o[259] = rdata_i[259];
  assign rdata_o[258] = rdata_i[258];
  assign rdata_o[257] = rdata_i[257];
  assign rdata_o[256] = rdata_i[256];
  assign rdata_o[255] = rdata_i[255];
  assign rdata_o[254] = rdata_i[254];
  assign rdata_o[253] = rdata_i[253];
  assign rdata_o[252] = rdata_i[252];
  assign rdata_o[251] = rdata_i[251];
  assign rdata_o[250] = rdata_i[250];
  assign rdata_o[249] = rdata_i[249];
  assign rdata_o[248] = rdata_i[248];
  assign rdata_o[247] = rdata_i[247];
  assign rdata_o[246] = rdata_i[246];
  assign rdata_o[245] = rdata_i[245];
  assign rdata_o[244] = rdata_i[244];
  assign rdata_o[243] = rdata_i[243];
  assign rdata_o[242] = rdata_i[242];
  assign rdata_o[241] = rdata_i[241];
  assign rdata_o[240] = rdata_i[240];
  assign rdata_o[239] = rdata_i[239];
  assign rdata_o[238] = rdata_i[238];
  assign rdata_o[237] = rdata_i[237];
  assign rdata_o[236] = rdata_i[236];
  assign rdata_o[235] = rdata_i[235];
  assign rdata_o[234] = rdata_i[234];
  assign rdata_o[233] = rdata_i[233];
  assign rdata_o[232] = rdata_i[232];
  assign rdata_o[231] = rdata_i[231];
  assign rdata_o[230] = rdata_i[230];
  assign rdata_o[229] = rdata_i[229];
  assign rdata_o[228] = rdata_i[228];
  assign rdata_o[227] = rdata_i[227];
  assign rdata_o[226] = rdata_i[226];
  assign rdata_o[225] = rdata_i[225];
  assign rdata_o[224] = rdata_i[224];
  assign rdata_o[223] = rdata_i[223];
  assign rdata_o[222] = rdata_i[222];
  assign rdata_o[221] = rdata_i[221];
  assign rdata_o[220] = rdata_i[220];
  assign rdata_o[219] = rdata_i[219];
  assign rdata_o[218] = rdata_i[218];
  assign rdata_o[217] = rdata_i[217];
  assign rdata_o[216] = rdata_i[216];
  assign rdata_o[215] = rdata_i[215];
  assign rdata_o[214] = rdata_i[214];
  assign rdata_o[213] = rdata_i[213];
  assign rdata_o[212] = rdata_i[212];
  assign rdata_o[211] = rdata_i[211];
  assign rdata_o[210] = rdata_i[210];
  assign rdata_o[209] = rdata_i[209];
  assign rdata_o[208] = rdata_i[208];
  assign rdata_o[207] = rdata_i[207];
  assign rdata_o[206] = rdata_i[206];
  assign rdata_o[205] = rdata_i[205];
  assign rdata_o[204] = rdata_i[204];
  assign rdata_o[203] = rdata_i[203];
  assign rdata_o[202] = rdata_i[202];
  assign rdata_o[201] = rdata_i[201];
  assign rdata_o[200] = rdata_i[200];
  assign rdata_o[199] = rdata_i[199];
  assign rdata_o[198] = rdata_i[198];
  assign rdata_o[197] = rdata_i[197];
  assign rdata_o[196] = rdata_i[196];
  assign rdata_o[195] = rdata_i[195];
  assign rdata_o[194] = rdata_i[194];
  assign rdata_o[193] = rdata_i[193];
  assign rdata_o[192] = rdata_i[192];
  assign rdata_o[191] = rdata_i[191];
  assign rdata_o[190] = rdata_i[190];
  assign rdata_o[189] = rdata_i[189];
  assign rdata_o[188] = rdata_i[188];
  assign rdata_o[187] = rdata_i[187];
  assign rdata_o[186] = rdata_i[186];
  assign rdata_o[185] = rdata_i[185];
  assign rdata_o[184] = rdata_i[184];
  assign rdata_o[183] = rdata_i[183];
  assign rdata_o[182] = rdata_i[182];
  assign rdata_o[181] = rdata_i[181];
  assign rdata_o[180] = rdata_i[180];
  assign rdata_o[179] = rdata_i[179];
  assign rdata_o[178] = rdata_i[178];
  assign rdata_o[177] = rdata_i[177];
  assign rdata_o[176] = rdata_i[176];
  assign rdata_o[175] = rdata_i[175];
  assign rdata_o[174] = rdata_i[174];
  assign rdata_o[173] = rdata_i[173];
  assign rdata_o[172] = rdata_i[172];
  assign rdata_o[171] = rdata_i[171];
  assign rdata_o[170] = rdata_i[170];
  assign rdata_o[169] = rdata_i[169];
  assign rdata_o[168] = rdata_i[168];
  assign rdata_o[167] = rdata_i[167];
  assign rdata_o[166] = rdata_i[166];
  assign rdata_o[165] = rdata_i[165];
  assign rdata_o[164] = rdata_i[164];
  assign rdata_o[163] = rdata_i[163];
  assign rdata_o[162] = rdata_i[162];
  assign rdata_o[161] = rdata_i[161];
  assign rdata_o[160] = rdata_i[160];
  assign rdata_o[159] = rdata_i[159];
  assign rdata_o[158] = rdata_i[158];
  assign rdata_o[157] = rdata_i[157];
  assign rdata_o[156] = rdata_i[156];
  assign rdata_o[155] = rdata_i[155];
  assign rdata_o[154] = rdata_i[154];
  assign rdata_o[153] = rdata_i[153];
  assign rdata_o[152] = rdata_i[152];
  assign rdata_o[151] = rdata_i[151];
  assign rdata_o[150] = rdata_i[150];
  assign rdata_o[149] = rdata_i[149];
  assign rdata_o[148] = rdata_i[148];
  assign rdata_o[147] = rdata_i[147];
  assign rdata_o[146] = rdata_i[146];
  assign rdata_o[145] = rdata_i[145];
  assign rdata_o[144] = rdata_i[144];
  assign rdata_o[143] = rdata_i[143];
  assign rdata_o[142] = rdata_i[142];
  assign rdata_o[141] = rdata_i[141];
  assign rdata_o[140] = rdata_i[140];
  assign rdata_o[139] = rdata_i[139];
  assign rdata_o[138] = rdata_i[138];
  assign rdata_o[137] = rdata_i[137];
  assign rdata_o[136] = rdata_i[136];
  assign rdata_o[135] = rdata_i[135];
  assign rdata_o[134] = rdata_i[134];
  assign rdata_o[133] = rdata_i[133];
  assign rdata_o[132] = rdata_i[132];
  assign rdata_o[131] = rdata_i[131];
  assign rdata_o[130] = rdata_i[130];
  assign rdata_o[129] = rdata_i[129];
  assign rdata_o[128] = rdata_i[128];
  assign rdata_o[127] = rdata_i[127];
  assign rdata_o[126] = rdata_i[126];
  assign rdata_o[125] = rdata_i[125];
  assign rdata_o[124] = rdata_i[124];
  assign rdata_o[123] = rdata_i[123];
  assign rdata_o[122] = rdata_i[122];
  assign rdata_o[121] = rdata_i[121];
  assign rdata_o[120] = rdata_i[120];
  assign rdata_o[119] = rdata_i[119];
  assign rdata_o[118] = rdata_i[118];
  assign rdata_o[117] = rdata_i[117];
  assign rdata_o[116] = rdata_i[116];
  assign rdata_o[115] = rdata_i[115];
  assign rdata_o[114] = rdata_i[114];
  assign rdata_o[113] = rdata_i[113];
  assign rdata_o[112] = rdata_i[112];
  assign rdata_o[111] = rdata_i[111];
  assign rdata_o[110] = rdata_i[110];
  assign rdata_o[109] = rdata_i[109];
  assign rdata_o[108] = rdata_i[108];
  assign rdata_o[107] = rdata_i[107];
  assign rdata_o[106] = rdata_i[106];
  assign rdata_o[105] = rdata_i[105];
  assign rdata_o[104] = rdata_i[104];
  assign rdata_o[103] = rdata_i[103];
  assign rdata_o[102] = rdata_i[102];
  assign rdata_o[101] = rdata_i[101];
  assign rdata_o[100] = rdata_i[100];
  assign rdata_o[99] = rdata_i[99];
  assign rdata_o[98] = rdata_i[98];
  assign rdata_o[97] = rdata_i[97];
  assign rdata_o[96] = rdata_i[96];
  assign rdata_o[95] = rdata_i[95];
  assign rdata_o[94] = rdata_i[94];
  assign rdata_o[93] = rdata_i[93];
  assign rdata_o[92] = rdata_i[92];
  assign rdata_o[91] = rdata_i[91];
  assign rdata_o[90] = rdata_i[90];
  assign rdata_o[89] = rdata_i[89];
  assign rdata_o[88] = rdata_i[88];
  assign rdata_o[87] = rdata_i[87];
  assign rdata_o[86] = rdata_i[86];
  assign rdata_o[85] = rdata_i[85];
  assign rdata_o[84] = rdata_i[84];
  assign rdata_o[83] = rdata_i[83];
  assign rdata_o[82] = rdata_i[82];
  assign rdata_o[81] = rdata_i[81];
  assign rdata_o[80] = rdata_i[80];
  assign rdata_o[79] = rdata_i[79];
  assign rdata_o[78] = rdata_i[78];
  assign rdata_o[77] = rdata_i[77];
  assign rdata_o[76] = rdata_i[76];
  assign rdata_o[75] = rdata_i[75];
  assign rdata_o[74] = rdata_i[74];
  assign rdata_o[73] = rdata_i[73];
  assign rdata_o[72] = rdata_i[72];
  assign rdata_o[71] = rdata_i[71];
  assign rdata_o[70] = rdata_i[70];
  assign rdata_o[69] = rdata_i[69];
  assign rdata_o[68] = rdata_i[68];
  assign rdata_o[67] = rdata_i[67];
  assign rdata_o[66] = rdata_i[66];
  assign rdata_o[65] = rdata_i[65];
  assign rdata_o[64] = rdata_i[64];
  assign rdata_o[63] = rdata_i[63];
  assign rdata_o[62] = rdata_i[62];
  assign rdata_o[61] = rdata_i[61];
  assign rdata_o[60] = rdata_i[60];
  assign rdata_o[59] = rdata_i[59];
  assign rdata_o[58] = rdata_i[58];
  assign rdata_o[57] = rdata_i[57];
  assign rdata_o[56] = rdata_i[56];
  assign rdata_o[55] = rdata_i[55];
  assign rdata_o[54] = rdata_i[54];
  assign rdata_o[53] = rdata_i[53];
  assign rdata_o[52] = rdata_i[52];
  assign rdata_o[51] = rdata_i[51];
  assign rdata_o[50] = rdata_i[50];
  assign rdata_o[49] = rdata_i[49];
  assign rdata_o[48] = rdata_i[48];
  assign rdata_o[47] = rdata_i[47];
  assign rdata_o[46] = rdata_i[46];
  assign rdata_o[45] = rdata_i[45];
  assign rdata_o[44] = rdata_i[44];
  assign rdata_o[43] = rdata_i[43];
  assign rdata_o[42] = rdata_i[42];
  assign rdata_o[41] = rdata_i[41];
  assign rdata_o[40] = rdata_i[40];
  assign rdata_o[39] = rdata_i[39];
  assign rdata_o[38] = rdata_i[38];
  assign rdata_o[37] = rdata_i[37];
  assign rdata_o[36] = rdata_i[36];
  assign rdata_o[35] = rdata_i[35];
  assign rdata_o[34] = rdata_i[34];
  assign rdata_o[33] = rdata_i[33];
  assign rdata_o[32] = rdata_i[32];
  assign rdata_o[31] = rdata_i[31];
  assign rdata_o[30] = rdata_i[30];
  assign rdata_o[29] = rdata_i[29];
  assign rdata_o[28] = rdata_i[28];
  assign rdata_o[27] = rdata_i[27];
  assign rdata_o[26] = rdata_i[26];
  assign rdata_o[25] = rdata_i[25];
  assign rdata_o[24] = rdata_i[24];
  assign rdata_o[23] = rdata_i[23];
  assign rdata_o[22] = rdata_i[22];
  assign rdata_o[21] = rdata_i[21];
  assign rdata_o[20] = rdata_i[20];
  assign rdata_o[19] = rdata_i[19];
  assign rdata_o[18] = rdata_i[18];
  assign rdata_o[17] = rdata_i[17];
  assign rdata_o[16] = rdata_i[16];
  assign rdata_o[15] = rdata_i[15];
  assign rdata_o[14] = rdata_i[14];
  assign rdata_o[13] = rdata_i[13];
  assign rdata_o[12] = rdata_i[12];
  assign rdata_o[11] = rdata_i[11];
  assign rdata_o[10] = rdata_i[10];
  assign rdata_o[9] = rdata_i[9];
  assign rdata_o[8] = rdata_i[8];
  assign rdata_o[7] = rdata_i[7];
  assign rdata_o[6] = rdata_i[6];
  assign rdata_o[5] = rdata_i[5];
  assign rdata_o[4] = rdata_i[4];
  assign rdata_o[3] = rdata_i[3];
  assign rdata_o[2] = rdata_i[2];
  assign rdata_o[1] = rdata_i[1];
  assign rdata_o[0] = rdata_i[0];
  assign N157 = sel_tag == rdata_i[173:130];
  assign N159 = sel_tag == rdata_i[347:304];
  assign N161 = sel_tag == rdata_i[521:478];
  assign N163 = sel_tag == rdata_i[695:652];
  assign N165 = sel_tag == rdata_i[869:826];
  assign N167 = sel_tag == rdata_i[1043:1000];
  assign N169 = sel_tag == rdata_i[1217:1174];
  assign N171 = sel_tag == rdata_i[1391:1348];

  always @(posedge clk_i or posedge N1325) begin
    if(N1325) begin
      id_q[3] <= 1'b0;
    end else if(1'b1) begin
      id_q[3] <= id_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1325) begin
    if(N1325) begin
      id_q[2] <= 1'b0;
    end else if(1'b1) begin
      id_q[2] <= id_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1325) begin
    if(N1325) begin
      id_q[1] <= 1'b0;
    end else if(1'b1) begin
      id_q[1] <= id_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1325) begin
    if(N1325) begin
      id_q[0] <= 1'b0;
    end else if(1'b1) begin
      id_q[0] <= id_d[0];
    end 
  end

  assign { N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22 } = (N0)? tag_i[43:0] : 
                                                                                                                                                                                                                                          (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = id_q[0];
  assign { N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67 } = (N1)? tag_i[87:44] : 
                                                                                                                                                                                                                                                     (N66)? { N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22 } : 1'b0;
  assign N1 = id_q[1];
  assign { N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112 } = (N2)? tag_i[131:88] : 
                                                                                                                                                                                                                                                                                      (N111)? { N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67 } : 1'b0;
  assign N2 = id_q[2];
  assign sel_tag = (N3)? tag_i[175:132] : 
                   (N156)? { N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112 } : 1'b0;
  assign N3 = id_q[3];
  assign hit_way_o[0] = (N4)? rdata_i[1] : 
                        (N158)? 1'b0 : 1'b0;
  assign N4 = N157;
  assign hit_way_o[1] = (N5)? rdata_i[175] : 
                        (N160)? 1'b0 : 1'b0;
  assign N5 = N159;
  assign hit_way_o[2] = (N6)? rdata_i[349] : 
                        (N162)? 1'b0 : 1'b0;
  assign N6 = N161;
  assign hit_way_o[3] = (N7)? rdata_i[523] : 
                        (N164)? 1'b0 : 1'b0;
  assign N7 = N163;
  assign hit_way_o[4] = (N8)? rdata_i[697] : 
                        (N166)? 1'b0 : 1'b0;
  assign N8 = N165;
  assign hit_way_o[5] = (N9)? rdata_i[871] : 
                        (N168)? 1'b0 : 1'b0;
  assign N9 = N167;
  assign hit_way_o[6] = (N10)? rdata_i[1045] : 
                        (N170)? 1'b0 : 1'b0;
  assign N10 = N169;
  assign hit_way_o[7] = (N11)? rdata_i[1219] : 
                        (N172)? 1'b0 : 1'b0;
  assign N11 = N171;
  assign N174 = ~N173;
  assign N178 = (N12)? 1'b0 : 
                (N177)? N174 : 1'b0;
  assign N12 = N176;
  assign N182 = (N13)? 1'b0 : 
                (N181)? N178 : 1'b0;
  assign N13 = N180;
  assign { N192, N191, N190, N189, N188, N187, N186, N185 } = (N14)? req_i[31:24] : 
                                                              (N184)? req_i[23:16] : 1'b0;
  assign N14 = N182;
  assign N193 = ~N182;
  assign { N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194 } = (N14)? addr_i[47:36] : 
                                                                                      (N184)? addr_i[35:24] : 1'b0;
  assign { N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206 } = (N14)? be_i[119:90] : 
                                                                                                                                                                                                  (N184)? be_i[89:60] : 1'b0;
  assign N236 = (N14)? we_i[3] : 
                (N184)? we_i[2] : 1'b0;
  assign { N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237 } = (N14)? wdata_i[695:522] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N184)? wdata_i[521:348] : 1'b0;
  assign { N418, N417, N416, N415, N414, N413, N412, N411 } = (N14)? { N192, N191, N190, N189, N188, N187, N186, N185 } : 
                                                              (N15)? req_i[23:16] : 1'b0;
  assign N15 = N183;
  assign { N420, N419 } = (N14)? { N182, N193 } : 
                          (N15)? { 1'b0, 1'b1 } : 1'b0;
  assign { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421 } = (N14)? { N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194 } : 
                                                                                      (N15)? addr_i[35:24] : 1'b0;
  assign { N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433 } = (N14)? { N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206 } : 
                                                                                                                                                                                                  (N15)? be_i[89:60] : 1'b0;
  assign N463 = (N14)? N236 : 
                (N15)? we_i[2] : 1'b0;
  assign { N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } = (N14)? { N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N15)? wdata_i[521:348] : 1'b0;
  assign { N646, N645, N644, N643, N642, N641, N640, N639 } = (N16)? { N418, N417, N416, N415, N414, N413, N412, N411 } : 
                                                              (N638)? req_i[15:8] : 1'b0;
  assign N16 = N178;
  assign N647 = ~N178;
  assign { N649, N648 } = (N16)? { N420, N419 } : 
                          (N638)? { 1'b0, 1'b0 } : 1'b0;
  assign { N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650 } = (N16)? { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421 } : 
                                                                                      (N638)? addr_i[23:12] : 1'b0;
  assign { N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662 } = (N16)? { N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433 } : 
                                                                                                                                                                                                  (N638)? be_i[59:30] : 1'b0;
  assign N692 = (N16)? N463 : 
                (N638)? we_i[1] : 1'b0;
  assign { N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693 } = (N16)? { N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N638)? wdata_i[347:174] : 1'b0;
  assign { N874, N873, N872, N871, N870, N869, N868, N867 } = (N16)? { N646, N645, N644, N643, N642, N641, N640, N639 } : 
                                                              (N17)? req_i[15:8] : 1'b0;
  assign N17 = N179;
  assign { N877, N876, N875 } = (N16)? { N649, N648, N647 } : 
                                (N17)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign N878 = (N16)? N178 : 
                (N17)? 1'b0 : 1'b0;
  assign { N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879 } = (N16)? { N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650 } : 
                                                                                      (N17)? addr_i[23:12] : 1'b0;
  assign { N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891 } = (N16)? { N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662 } : 
                                                                                                                                                                                                  (N17)? be_i[59:30] : 1'b0;
  assign N921 = (N16)? N692 : 
                (N17)? we_i[1] : 1'b0;
  assign { N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922 } = (N16)? { N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N17)? wdata_i[347:174] : 1'b0;
  assign { N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096 } = (N18)? { N874, N873, N872, N871, N870, N869, N868, N867 } : 
                                                                      (N19)? req_i[7:0] : 1'b0;
  assign N18 = N175;
  assign N19 = N173;
  assign { N1106, N1105, N1104 } = (N18)? { N877, N876, N875 } : 
                                   (N19)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1107 = (N18)? N878 : 
                 (N19)? 1'b0 : 1'b0;
  assign { N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108 } = (N18)? { N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879 } : 
                                                                                                  (N19)? addr_i[11:0] : 1'b0;
  assign { N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120 } = (N18)? { N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891 } : 
                                                                                                                                                                                                                                (N19)? be_i[29:0] : 1'b0;
  assign N1150 = (N18)? N921 : 
                 (N19)? we_i[0] : 1'b0;
  assign { N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151 } = (N18)? { N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N19)? wdata_i[173:0] : 1'b0;
  assign req_o = (N20)? { N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096 } : 
                 (N19)? req_i[7:0] : 1'b0;
  assign N20 = N174;
  assign id_d = (N20)? { N1106, N1105, N1104, N173 } : 
                (N19)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign gnt_o[3:1] = (N20)? { N1106, N1107, N175 } : 
                      (N19)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign addr_o = (N20)? { N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108 } : 
                  (N19)? addr_i[11:0] : 1'b0;
  assign be_o = (N20)? { N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120 } : 
                (N19)? be_i[29:0] : 1'b0;
  assign we_o = (N20)? N1150 : 
                (N19)? we_i[0] : 1'b0;
  assign wdata_o = (N20)? { N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151 } : 
                   (N19)? wdata_i[173:0] : 1'b0;
  assign N21 = ~id_q[0];
  assign N66 = ~id_q[1];
  assign N111 = ~id_q[2];
  assign N156 = ~id_q[3];
  assign N158 = ~N157;
  assign N160 = ~N159;
  assign N162 = ~N161;
  assign N164 = ~N163;
  assign N166 = ~N165;
  assign N168 = ~N167;
  assign N170 = ~N169;
  assign N172 = ~N171;
  assign N173 = N1331 | req_i[0];
  assign N1331 = N1330 | req_i[1];
  assign N1330 = N1329 | req_i[2];
  assign N1329 = N1328 | req_i[3];
  assign N1328 = N1327 | req_i[4];
  assign N1327 = N1326 | req_i[5];
  assign N1326 = req_i[7] | req_i[6];
  assign N175 = ~N173;
  assign N176 = N1337 | req_i[8];
  assign N1337 = N1336 | req_i[9];
  assign N1336 = N1335 | req_i[10];
  assign N1335 = N1334 | req_i[11];
  assign N1334 = N1333 | req_i[12];
  assign N1333 = N1332 | req_i[13];
  assign N1332 = req_i[15] | req_i[14];
  assign N177 = ~N176;
  assign N179 = ~N178;
  assign N180 = N1343 | req_i[16];
  assign N1343 = N1342 | req_i[17];
  assign N1342 = N1341 | req_i[18];
  assign N1341 = N1340 | req_i[19];
  assign N1340 = N1339 | req_i[20];
  assign N1339 = N1338 | req_i[21];
  assign N1338 = req_i[23] | req_i[22];
  assign N181 = ~N180;
  assign N183 = ~N182;
  assign N184 = ~N182;
  assign N638 = ~N178;
  assign N1325 = ~rst_ni;

endmodule