module bsg_mem_1r1w_synth_width_p256_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [255:0] w_data_i;
  input [0:0] r_addr_i;
  output [255:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [255:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12;
  wire [511:0] mem;
  reg mem_511_sv2v_reg,mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,
  mem_507_sv2v_reg,mem_506_sv2v_reg,mem_505_sv2v_reg,mem_504_sv2v_reg,mem_503_sv2v_reg,
  mem_502_sv2v_reg,mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,mem_498_sv2v_reg,
  mem_497_sv2v_reg,mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,
  mem_493_sv2v_reg,mem_492_sv2v_reg,mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,
  mem_488_sv2v_reg,mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,mem_484_sv2v_reg,
  mem_483_sv2v_reg,mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,
  mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,
  mem_474_sv2v_reg,mem_473_sv2v_reg,mem_472_sv2v_reg,mem_471_sv2v_reg,mem_470_sv2v_reg,
  mem_469_sv2v_reg,mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,mem_465_sv2v_reg,
  mem_464_sv2v_reg,mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,
  mem_460_sv2v_reg,mem_459_sv2v_reg,mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,
  mem_455_sv2v_reg,mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,mem_451_sv2v_reg,
  mem_450_sv2v_reg,mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,
  mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,
  mem_441_sv2v_reg,mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,
  mem_436_sv2v_reg,mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,
  mem_431_sv2v_reg,mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,
  mem_427_sv2v_reg,mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,mem_423_sv2v_reg,
  mem_422_sv2v_reg,mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,
  mem_417_sv2v_reg,mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,
  mem_413_sv2v_reg,mem_412_sv2v_reg,mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,
  mem_408_sv2v_reg,mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,
  mem_403_sv2v_reg,mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,
  mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,
  mem_394_sv2v_reg,mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,mem_390_sv2v_reg,
  mem_389_sv2v_reg,mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,
  mem_384_sv2v_reg,mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,
  mem_380_sv2v_reg,mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,
  mem_375_sv2v_reg,mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,
  mem_370_sv2v_reg,mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,
  mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,
  mem_361_sv2v_reg,mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,
  mem_356_sv2v_reg,mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,
  mem_351_sv2v_reg,mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,
  mem_347_sv2v_reg,mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,mem_343_sv2v_reg,
  mem_342_sv2v_reg,mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,
  mem_337_sv2v_reg,mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,
  mem_333_sv2v_reg,mem_332_sv2v_reg,mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,
  mem_328_sv2v_reg,mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,
  mem_323_sv2v_reg,mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,
  mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,
  mem_314_sv2v_reg,mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,mem_310_sv2v_reg,
  mem_309_sv2v_reg,mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,
  mem_304_sv2v_reg,mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,
  mem_300_sv2v_reg,mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,
  mem_295_sv2v_reg,mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,
  mem_290_sv2v_reg,mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,
  mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,
  mem_281_sv2v_reg,mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,
  mem_276_sv2v_reg,mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,
  mem_271_sv2v_reg,mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,
  mem_267_sv2v_reg,mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,mem_263_sv2v_reg,
  mem_262_sv2v_reg,mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,
  mem_257_sv2v_reg,mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,
  mem_253_sv2v_reg,mem_252_sv2v_reg,mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,
  mem_248_sv2v_reg,mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,
  mem_243_sv2v_reg,mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,
  mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,
  mem_234_sv2v_reg,mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,
  mem_229_sv2v_reg,mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,
  mem_224_sv2v_reg,mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,
  mem_220_sv2v_reg,mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,
  mem_215_sv2v_reg,mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,
  mem_210_sv2v_reg,mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,
  mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,
  mem_201_sv2v_reg,mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,
  mem_196_sv2v_reg,mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,
  mem_191_sv2v_reg,mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,
  mem_187_sv2v_reg,mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,
  mem_182_sv2v_reg,mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,
  mem_177_sv2v_reg,mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,
  mem_173_sv2v_reg,mem_172_sv2v_reg,mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,
  mem_168_sv2v_reg,mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,
  mem_163_sv2v_reg,mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,
  mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,
  mem_154_sv2v_reg,mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,
  mem_149_sv2v_reg,mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,
  mem_144_sv2v_reg,mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,
  mem_140_sv2v_reg,mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,
  mem_135_sv2v_reg,mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,
  mem_130_sv2v_reg,mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,
  mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,
  mem_121_sv2v_reg,mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,
  mem_116_sv2v_reg,mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,
  mem_111_sv2v_reg,mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,
  mem_107_sv2v_reg,mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,
  mem_102_sv2v_reg,mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,
  mem_97_sv2v_reg,mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,
  mem_92_sv2v_reg,mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,
  mem_87_sv2v_reg,mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,
  mem_82_sv2v_reg,mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,
  mem_77_sv2v_reg,mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,
  mem_72_sv2v_reg,mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,
  mem_67_sv2v_reg,mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,
  mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,
  mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,
  mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,
  mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,
  mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,
  mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,
  mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,
  mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,
  mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,
  mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,
  mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,
  mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,
  mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[255] = (N3)? mem[255] : 
                         (N0)? mem[511] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[254] = (N3)? mem[254] : 
                         (N0)? mem[510] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] : 
                         (N0)? mem[509] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] : 
                         (N0)? mem[508] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] : 
                         (N0)? mem[507] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] : 
                         (N0)? mem[506] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] : 
                         (N0)? mem[505] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] : 
                         (N0)? mem[504] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] : 
                         (N0)? mem[503] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] : 
                         (N0)? mem[502] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] : 
                         (N0)? mem[501] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] : 
                         (N0)? mem[500] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] : 
                         (N0)? mem[499] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] : 
                         (N0)? mem[498] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] : 
                         (N0)? mem[497] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] : 
                         (N0)? mem[496] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] : 
                         (N0)? mem[495] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] : 
                         (N0)? mem[494] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] : 
                         (N0)? mem[493] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] : 
                         (N0)? mem[492] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] : 
                         (N0)? mem[491] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] : 
                         (N0)? mem[490] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] : 
                         (N0)? mem[489] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] : 
                         (N0)? mem[488] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] : 
                         (N0)? mem[487] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] : 
                         (N0)? mem[486] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] : 
                         (N0)? mem[485] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] : 
                         (N0)? mem[484] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] : 
                         (N0)? mem[483] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] : 
                         (N0)? mem[482] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] : 
                         (N0)? mem[481] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] : 
                         (N0)? mem[480] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] : 
                         (N0)? mem[479] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] : 
                         (N0)? mem[478] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] : 
                         (N0)? mem[477] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] : 
                         (N0)? mem[476] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] : 
                         (N0)? mem[475] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] : 
                         (N0)? mem[474] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] : 
                         (N0)? mem[473] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] : 
                         (N0)? mem[472] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] : 
                         (N0)? mem[471] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] : 
                         (N0)? mem[470] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] : 
                         (N0)? mem[469] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] : 
                         (N0)? mem[468] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] : 
                         (N0)? mem[467] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] : 
                         (N0)? mem[466] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] : 
                         (N0)? mem[465] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] : 
                         (N0)? mem[464] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] : 
                         (N0)? mem[463] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] : 
                         (N0)? mem[462] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] : 
                         (N0)? mem[461] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] : 
                         (N0)? mem[460] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] : 
                         (N0)? mem[459] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] : 
                         (N0)? mem[458] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] : 
                         (N0)? mem[457] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] : 
                         (N0)? mem[456] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] : 
                         (N0)? mem[455] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] : 
                         (N0)? mem[454] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] : 
                         (N0)? mem[453] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] : 
                         (N0)? mem[452] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] : 
                         (N0)? mem[451] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] : 
                         (N0)? mem[450] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] : 
                         (N0)? mem[449] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] : 
                         (N0)? mem[448] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] : 
                         (N0)? mem[447] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] : 
                         (N0)? mem[446] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] : 
                         (N0)? mem[445] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] : 
                         (N0)? mem[444] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] : 
                         (N0)? mem[443] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] : 
                         (N0)? mem[442] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] : 
                         (N0)? mem[441] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] : 
                         (N0)? mem[440] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] : 
                         (N0)? mem[439] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] : 
                         (N0)? mem[438] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] : 
                         (N0)? mem[437] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] : 
                         (N0)? mem[436] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] : 
                         (N0)? mem[435] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] : 
                         (N0)? mem[434] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] : 
                         (N0)? mem[433] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] : 
                         (N0)? mem[432] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] : 
                         (N0)? mem[431] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] : 
                         (N0)? mem[430] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] : 
                         (N0)? mem[429] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] : 
                         (N0)? mem[428] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] : 
                         (N0)? mem[427] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] : 
                         (N0)? mem[426] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] : 
                         (N0)? mem[425] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] : 
                         (N0)? mem[424] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] : 
                         (N0)? mem[423] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] : 
                         (N0)? mem[422] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] : 
                         (N0)? mem[421] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] : 
                         (N0)? mem[420] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] : 
                         (N0)? mem[419] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] : 
                         (N0)? mem[418] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] : 
                         (N0)? mem[417] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] : 
                         (N0)? mem[416] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] : 
                         (N0)? mem[415] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] : 
                         (N0)? mem[414] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] : 
                         (N0)? mem[413] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] : 
                         (N0)? mem[412] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] : 
                         (N0)? mem[411] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] : 
                         (N0)? mem[410] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] : 
                         (N0)? mem[409] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] : 
                         (N0)? mem[408] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] : 
                         (N0)? mem[407] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] : 
                         (N0)? mem[406] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] : 
                         (N0)? mem[405] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] : 
                         (N0)? mem[404] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] : 
                         (N0)? mem[403] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] : 
                         (N0)? mem[402] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] : 
                         (N0)? mem[401] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] : 
                         (N0)? mem[400] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] : 
                         (N0)? mem[399] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] : 
                         (N0)? mem[398] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] : 
                         (N0)? mem[397] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] : 
                         (N0)? mem[396] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] : 
                         (N0)? mem[395] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] : 
                         (N0)? mem[394] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] : 
                         (N0)? mem[393] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] : 
                         (N0)? mem[392] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] : 
                         (N0)? mem[391] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] : 
                         (N0)? mem[390] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] : 
                         (N0)? mem[389] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] : 
                         (N0)? mem[388] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] : 
                         (N0)? mem[387] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] : 
                         (N0)? mem[386] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] : 
                         (N0)? mem[385] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] : 
                         (N0)? mem[384] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[383] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[382] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[381] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[380] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[379] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[378] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[377] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[376] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[375] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[374] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[373] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[372] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[371] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[370] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[369] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[368] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[367] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[366] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[365] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[364] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[363] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[362] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[361] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[360] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[359] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[358] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[357] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[356] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[355] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[354] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[353] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[352] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[351] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[350] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[349] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[348] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[347] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[346] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[345] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[344] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[343] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[342] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[341] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[340] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[339] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[338] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[337] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[336] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[335] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[334] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[333] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[332] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[331] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[330] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[329] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[328] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[327] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[326] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[325] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[324] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[323] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[322] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[321] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[320] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[319] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[318] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[317] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[316] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[315] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[314] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[313] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[312] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[311] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[310] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[309] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[308] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[307] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[306] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[305] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[304] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[303] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[302] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[301] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[300] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[299] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[298] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[297] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[296] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[295] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[294] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[293] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[292] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[291] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[290] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[289] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[288] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[287] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[286] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[285] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[284] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[283] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[282] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[281] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[280] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[279] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[278] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[277] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[276] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[275] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[274] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[273] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[272] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[271] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[270] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[269] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[268] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[267] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[266] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[265] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[264] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[263] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[262] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[261] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[260] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[259] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[258] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[257] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[256] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_511_sv2v_reg <= w_data_i[255];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_510_sv2v_reg <= w_data_i[254];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_509_sv2v_reg <= w_data_i[253];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_508_sv2v_reg <= w_data_i[252];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_507_sv2v_reg <= w_data_i[251];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_506_sv2v_reg <= w_data_i[250];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_505_sv2v_reg <= w_data_i[249];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_504_sv2v_reg <= w_data_i[248];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_503_sv2v_reg <= w_data_i[247];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_502_sv2v_reg <= w_data_i[246];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_501_sv2v_reg <= w_data_i[245];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_500_sv2v_reg <= w_data_i[244];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_499_sv2v_reg <= w_data_i[243];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_498_sv2v_reg <= w_data_i[242];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_497_sv2v_reg <= w_data_i[241];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_496_sv2v_reg <= w_data_i[240];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_495_sv2v_reg <= w_data_i[239];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_494_sv2v_reg <= w_data_i[238];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_493_sv2v_reg <= w_data_i[237];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_492_sv2v_reg <= w_data_i[236];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_491_sv2v_reg <= w_data_i[235];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_490_sv2v_reg <= w_data_i[234];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_489_sv2v_reg <= w_data_i[233];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_488_sv2v_reg <= w_data_i[232];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_487_sv2v_reg <= w_data_i[231];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_486_sv2v_reg <= w_data_i[230];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_485_sv2v_reg <= w_data_i[229];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_484_sv2v_reg <= w_data_i[228];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_483_sv2v_reg <= w_data_i[227];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_482_sv2v_reg <= w_data_i[226];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_481_sv2v_reg <= w_data_i[225];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_480_sv2v_reg <= w_data_i[224];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_479_sv2v_reg <= w_data_i[223];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_478_sv2v_reg <= w_data_i[222];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_477_sv2v_reg <= w_data_i[221];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_476_sv2v_reg <= w_data_i[220];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_475_sv2v_reg <= w_data_i[219];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_474_sv2v_reg <= w_data_i[218];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_473_sv2v_reg <= w_data_i[217];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_472_sv2v_reg <= w_data_i[216];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_471_sv2v_reg <= w_data_i[215];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_470_sv2v_reg <= w_data_i[214];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_469_sv2v_reg <= w_data_i[213];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_468_sv2v_reg <= w_data_i[212];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_467_sv2v_reg <= w_data_i[211];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_466_sv2v_reg <= w_data_i[210];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_465_sv2v_reg <= w_data_i[209];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_464_sv2v_reg <= w_data_i[208];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_463_sv2v_reg <= w_data_i[207];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_462_sv2v_reg <= w_data_i[206];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_461_sv2v_reg <= w_data_i[205];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_460_sv2v_reg <= w_data_i[204];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_459_sv2v_reg <= w_data_i[203];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_458_sv2v_reg <= w_data_i[202];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_457_sv2v_reg <= w_data_i[201];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_456_sv2v_reg <= w_data_i[200];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_455_sv2v_reg <= w_data_i[199];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_454_sv2v_reg <= w_data_i[198];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_453_sv2v_reg <= w_data_i[197];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_452_sv2v_reg <= w_data_i[196];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_451_sv2v_reg <= w_data_i[195];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_450_sv2v_reg <= w_data_i[194];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_449_sv2v_reg <= w_data_i[193];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_448_sv2v_reg <= w_data_i[192];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_447_sv2v_reg <= w_data_i[191];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_446_sv2v_reg <= w_data_i[190];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_445_sv2v_reg <= w_data_i[189];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_444_sv2v_reg <= w_data_i[188];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_443_sv2v_reg <= w_data_i[187];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_442_sv2v_reg <= w_data_i[186];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_441_sv2v_reg <= w_data_i[185];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_440_sv2v_reg <= w_data_i[184];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_439_sv2v_reg <= w_data_i[183];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_438_sv2v_reg <= w_data_i[182];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_437_sv2v_reg <= w_data_i[181];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_436_sv2v_reg <= w_data_i[180];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_435_sv2v_reg <= w_data_i[179];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_434_sv2v_reg <= w_data_i[178];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_433_sv2v_reg <= w_data_i[177];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_432_sv2v_reg <= w_data_i[176];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_431_sv2v_reg <= w_data_i[175];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_430_sv2v_reg <= w_data_i[174];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_429_sv2v_reg <= w_data_i[173];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_428_sv2v_reg <= w_data_i[172];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_427_sv2v_reg <= w_data_i[171];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_426_sv2v_reg <= w_data_i[170];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_425_sv2v_reg <= w_data_i[169];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_424_sv2v_reg <= w_data_i[168];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_423_sv2v_reg <= w_data_i[167];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_422_sv2v_reg <= w_data_i[166];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_421_sv2v_reg <= w_data_i[165];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_420_sv2v_reg <= w_data_i[164];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_419_sv2v_reg <= w_data_i[163];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_418_sv2v_reg <= w_data_i[162];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_417_sv2v_reg <= w_data_i[161];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_416_sv2v_reg <= w_data_i[160];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_415_sv2v_reg <= w_data_i[159];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_414_sv2v_reg <= w_data_i[158];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_413_sv2v_reg <= w_data_i[157];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_412_sv2v_reg <= w_data_i[156];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_411_sv2v_reg <= w_data_i[155];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_410_sv2v_reg <= w_data_i[154];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_409_sv2v_reg <= w_data_i[153];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_408_sv2v_reg <= w_data_i[152];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_407_sv2v_reg <= w_data_i[151];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_406_sv2v_reg <= w_data_i[150];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_405_sv2v_reg <= w_data_i[149];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_404_sv2v_reg <= w_data_i[148];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_403_sv2v_reg <= w_data_i[147];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_402_sv2v_reg <= w_data_i[146];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_401_sv2v_reg <= w_data_i[145];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_400_sv2v_reg <= w_data_i[144];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_399_sv2v_reg <= w_data_i[143];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_398_sv2v_reg <= w_data_i[142];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_397_sv2v_reg <= w_data_i[141];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_396_sv2v_reg <= w_data_i[140];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_395_sv2v_reg <= w_data_i[139];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_394_sv2v_reg <= w_data_i[138];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_393_sv2v_reg <= w_data_i[137];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_392_sv2v_reg <= w_data_i[136];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_391_sv2v_reg <= w_data_i[135];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_390_sv2v_reg <= w_data_i[134];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_389_sv2v_reg <= w_data_i[133];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_388_sv2v_reg <= w_data_i[132];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_387_sv2v_reg <= w_data_i[131];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_386_sv2v_reg <= w_data_i[130];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_385_sv2v_reg <= w_data_i[129];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_384_sv2v_reg <= w_data_i[128];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_383_sv2v_reg <= w_data_i[127];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_382_sv2v_reg <= w_data_i[126];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_381_sv2v_reg <= w_data_i[125];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_380_sv2v_reg <= w_data_i[124];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_379_sv2v_reg <= w_data_i[123];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_378_sv2v_reg <= w_data_i[122];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_377_sv2v_reg <= w_data_i[121];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_376_sv2v_reg <= w_data_i[120];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_375_sv2v_reg <= w_data_i[119];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_374_sv2v_reg <= w_data_i[118];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_373_sv2v_reg <= w_data_i[117];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_372_sv2v_reg <= w_data_i[116];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_371_sv2v_reg <= w_data_i[115];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_370_sv2v_reg <= w_data_i[114];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_369_sv2v_reg <= w_data_i[113];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_368_sv2v_reg <= w_data_i[112];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_367_sv2v_reg <= w_data_i[111];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_366_sv2v_reg <= w_data_i[110];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_365_sv2v_reg <= w_data_i[109];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_364_sv2v_reg <= w_data_i[108];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_363_sv2v_reg <= w_data_i[107];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_362_sv2v_reg <= w_data_i[106];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_361_sv2v_reg <= w_data_i[105];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_360_sv2v_reg <= w_data_i[104];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_359_sv2v_reg <= w_data_i[103];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_358_sv2v_reg <= w_data_i[102];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_357_sv2v_reg <= w_data_i[101];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_356_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_355_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_354_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_353_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_352_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_351_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_350_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_349_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_348_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_347_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_346_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_345_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_344_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_343_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_342_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_341_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_340_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_339_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_338_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_337_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_336_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_335_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_334_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_333_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_332_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_331_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_330_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_329_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_328_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_327_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_326_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_325_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_324_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_323_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_322_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_321_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_320_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_319_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_318_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_317_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_316_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_315_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_314_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_313_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_312_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_311_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_310_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_309_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_308_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_307_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_306_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_305_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_304_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_303_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_302_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_301_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_300_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_299_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_298_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_297_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_296_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_295_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_294_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_293_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_292_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_291_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_290_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_289_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_288_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_287_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_286_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_285_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_284_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_283_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_282_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_281_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_280_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_279_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_278_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_277_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_276_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_275_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_274_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_273_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_272_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_271_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_270_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_269_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_268_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_267_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_266_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_265_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_264_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_263_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_262_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_261_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_260_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_259_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N12) begin
      mem_258_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N11) begin
      mem_257_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N10) begin
      mem_256_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_255_sv2v_reg <= w_data_i[255];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_254_sv2v_reg <= w_data_i[254];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_253_sv2v_reg <= w_data_i[253];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_252_sv2v_reg <= w_data_i[252];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_251_sv2v_reg <= w_data_i[251];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_250_sv2v_reg <= w_data_i[250];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_249_sv2v_reg <= w_data_i[249];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_248_sv2v_reg <= w_data_i[248];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_247_sv2v_reg <= w_data_i[247];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_246_sv2v_reg <= w_data_i[246];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_245_sv2v_reg <= w_data_i[245];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_244_sv2v_reg <= w_data_i[244];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_243_sv2v_reg <= w_data_i[243];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_242_sv2v_reg <= w_data_i[242];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_241_sv2v_reg <= w_data_i[241];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_240_sv2v_reg <= w_data_i[240];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_239_sv2v_reg <= w_data_i[239];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_238_sv2v_reg <= w_data_i[238];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_237_sv2v_reg <= w_data_i[237];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_236_sv2v_reg <= w_data_i[236];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_235_sv2v_reg <= w_data_i[235];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_234_sv2v_reg <= w_data_i[234];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_233_sv2v_reg <= w_data_i[233];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_232_sv2v_reg <= w_data_i[232];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_231_sv2v_reg <= w_data_i[231];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_230_sv2v_reg <= w_data_i[230];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_229_sv2v_reg <= w_data_i[229];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_228_sv2v_reg <= w_data_i[228];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_227_sv2v_reg <= w_data_i[227];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_226_sv2v_reg <= w_data_i[226];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_225_sv2v_reg <= w_data_i[225];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_224_sv2v_reg <= w_data_i[224];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_223_sv2v_reg <= w_data_i[223];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_222_sv2v_reg <= w_data_i[222];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_221_sv2v_reg <= w_data_i[221];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_220_sv2v_reg <= w_data_i[220];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_219_sv2v_reg <= w_data_i[219];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_218_sv2v_reg <= w_data_i[218];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_217_sv2v_reg <= w_data_i[217];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_216_sv2v_reg <= w_data_i[216];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_215_sv2v_reg <= w_data_i[215];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_214_sv2v_reg <= w_data_i[214];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_213_sv2v_reg <= w_data_i[213];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_212_sv2v_reg <= w_data_i[212];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_211_sv2v_reg <= w_data_i[211];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_210_sv2v_reg <= w_data_i[210];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_209_sv2v_reg <= w_data_i[209];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_208_sv2v_reg <= w_data_i[208];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_207_sv2v_reg <= w_data_i[207];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_206_sv2v_reg <= w_data_i[206];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_205_sv2v_reg <= w_data_i[205];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_204_sv2v_reg <= w_data_i[204];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_203_sv2v_reg <= w_data_i[203];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_202_sv2v_reg <= w_data_i[202];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_201_sv2v_reg <= w_data_i[201];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_200_sv2v_reg <= w_data_i[200];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_199_sv2v_reg <= w_data_i[199];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_198_sv2v_reg <= w_data_i[198];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_197_sv2v_reg <= w_data_i[197];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_196_sv2v_reg <= w_data_i[196];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_195_sv2v_reg <= w_data_i[195];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_194_sv2v_reg <= w_data_i[194];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_193_sv2v_reg <= w_data_i[193];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_192_sv2v_reg <= w_data_i[192];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_191_sv2v_reg <= w_data_i[191];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_190_sv2v_reg <= w_data_i[190];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_189_sv2v_reg <= w_data_i[189];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_188_sv2v_reg <= w_data_i[188];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_187_sv2v_reg <= w_data_i[187];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_186_sv2v_reg <= w_data_i[186];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_185_sv2v_reg <= w_data_i[185];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_184_sv2v_reg <= w_data_i[184];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_183_sv2v_reg <= w_data_i[183];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_182_sv2v_reg <= w_data_i[182];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_181_sv2v_reg <= w_data_i[181];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_180_sv2v_reg <= w_data_i[180];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_179_sv2v_reg <= w_data_i[179];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_178_sv2v_reg <= w_data_i[178];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_177_sv2v_reg <= w_data_i[177];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_176_sv2v_reg <= w_data_i[176];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_175_sv2v_reg <= w_data_i[175];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_174_sv2v_reg <= w_data_i[174];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_173_sv2v_reg <= w_data_i[173];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_172_sv2v_reg <= w_data_i[172];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_171_sv2v_reg <= w_data_i[171];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_170_sv2v_reg <= w_data_i[170];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_169_sv2v_reg <= w_data_i[169];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_168_sv2v_reg <= w_data_i[168];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_167_sv2v_reg <= w_data_i[167];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_166_sv2v_reg <= w_data_i[166];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_165_sv2v_reg <= w_data_i[165];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_164_sv2v_reg <= w_data_i[164];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_163_sv2v_reg <= w_data_i[163];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_162_sv2v_reg <= w_data_i[162];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_161_sv2v_reg <= w_data_i[161];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_160_sv2v_reg <= w_data_i[160];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_159_sv2v_reg <= w_data_i[159];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_158_sv2v_reg <= w_data_i[158];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_157_sv2v_reg <= w_data_i[157];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_156_sv2v_reg <= w_data_i[156];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_155_sv2v_reg <= w_data_i[155];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_154_sv2v_reg <= w_data_i[154];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_153_sv2v_reg <= w_data_i[153];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_152_sv2v_reg <= w_data_i[152];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_151_sv2v_reg <= w_data_i[151];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_150_sv2v_reg <= w_data_i[150];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_149_sv2v_reg <= w_data_i[149];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_148_sv2v_reg <= w_data_i[148];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_147_sv2v_reg <= w_data_i[147];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_146_sv2v_reg <= w_data_i[146];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_145_sv2v_reg <= w_data_i[145];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_144_sv2v_reg <= w_data_i[144];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_143_sv2v_reg <= w_data_i[143];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_142_sv2v_reg <= w_data_i[142];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_141_sv2v_reg <= w_data_i[141];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_140_sv2v_reg <= w_data_i[140];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_139_sv2v_reg <= w_data_i[139];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_138_sv2v_reg <= w_data_i[138];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_137_sv2v_reg <= w_data_i[137];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_136_sv2v_reg <= w_data_i[136];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_135_sv2v_reg <= w_data_i[135];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_134_sv2v_reg <= w_data_i[134];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_133_sv2v_reg <= w_data_i[133];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_132_sv2v_reg <= w_data_i[132];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_131_sv2v_reg <= w_data_i[131];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_130_sv2v_reg <= w_data_i[130];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_129_sv2v_reg <= w_data_i[129];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_128_sv2v_reg <= w_data_i[128];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_127_sv2v_reg <= w_data_i[127];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_126_sv2v_reg <= w_data_i[126];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_125_sv2v_reg <= w_data_i[125];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_124_sv2v_reg <= w_data_i[124];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_123_sv2v_reg <= w_data_i[123];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_122_sv2v_reg <= w_data_i[122];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_121_sv2v_reg <= w_data_i[121];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_120_sv2v_reg <= w_data_i[120];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_119_sv2v_reg <= w_data_i[119];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_118_sv2v_reg <= w_data_i[118];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_117_sv2v_reg <= w_data_i[117];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_116_sv2v_reg <= w_data_i[116];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_115_sv2v_reg <= w_data_i[115];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_114_sv2v_reg <= w_data_i[114];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_113_sv2v_reg <= w_data_i[113];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_112_sv2v_reg <= w_data_i[112];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_111_sv2v_reg <= w_data_i[111];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_110_sv2v_reg <= w_data_i[110];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_109_sv2v_reg <= w_data_i[109];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_108_sv2v_reg <= w_data_i[108];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_107_sv2v_reg <= w_data_i[107];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_106_sv2v_reg <= w_data_i[106];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_105_sv2v_reg <= w_data_i[105];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_104_sv2v_reg <= w_data_i[104];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_103_sv2v_reg <= w_data_i[103];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_102_sv2v_reg <= w_data_i[102];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_101_sv2v_reg <= w_data_i[101];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_100_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_99_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_98_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_97_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_96_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_95_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_94_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_93_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_92_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_91_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_90_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_89_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_88_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_87_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_86_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_85_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_84_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_83_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_82_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_81_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_80_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_79_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_78_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_77_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_76_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_75_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_74_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_73_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_72_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_71_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_70_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_69_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_68_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_67_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_66_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_65_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_64_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_63_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_62_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_61_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_60_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_59_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_58_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_57_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_56_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_55_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_54_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_53_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_52_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_51_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_50_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_49_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_48_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_47_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_46_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_45_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_44_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_43_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_42_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_41_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_40_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_39_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_38_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_37_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_36_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_35_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_34_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_33_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_32_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_31_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_30_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_29_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_28_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_27_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_26_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_25_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_24_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_23_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_22_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_21_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_20_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_19_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_18_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_17_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_16_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_15_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_14_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_13_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_12_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_11_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_10_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_9_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_8_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_7_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_6_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_5_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_4_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_3_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N9) begin
      mem_2_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_1_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N7) begin
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end

  assign N5 = ~w_addr_i[0];
  assign { N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5 } : 
                                         (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

endmodule