module bsg_mesh_stitch_width_p64_x_max_p2_y_max_p2
(
  outs_i,
  ins_o,
  hor_i,
  hor_o,
  ver_i,
  ver_o
);

  input [1023:0] outs_i;
  output [1023:0] ins_o;
  input [255:0] hor_i;
  output [255:0] hor_o;
  input [255:0] ver_i;
  output [255:0] ver_o;
  wire [1023:0] ins_o;
  wire [255:0] hor_o,ver_o;
  assign ins_o[1023] = ver_i[255];
  assign ins_o[1022] = ver_i[254];
  assign ins_o[1021] = ver_i[253];
  assign ins_o[1020] = ver_i[252];
  assign ins_o[1019] = ver_i[251];
  assign ins_o[1018] = ver_i[250];
  assign ins_o[1017] = ver_i[249];
  assign ins_o[1016] = ver_i[248];
  assign ins_o[1015] = ver_i[247];
  assign ins_o[1014] = ver_i[246];
  assign ins_o[1013] = ver_i[245];
  assign ins_o[1012] = ver_i[244];
  assign ins_o[1011] = ver_i[243];
  assign ins_o[1010] = ver_i[242];
  assign ins_o[1009] = ver_i[241];
  assign ins_o[1008] = ver_i[240];
  assign ins_o[1007] = ver_i[239];
  assign ins_o[1006] = ver_i[238];
  assign ins_o[1005] = ver_i[237];
  assign ins_o[1004] = ver_i[236];
  assign ins_o[1003] = ver_i[235];
  assign ins_o[1002] = ver_i[234];
  assign ins_o[1001] = ver_i[233];
  assign ins_o[1000] = ver_i[232];
  assign ins_o[999] = ver_i[231];
  assign ins_o[998] = ver_i[230];
  assign ins_o[997] = ver_i[229];
  assign ins_o[996] = ver_i[228];
  assign ins_o[995] = ver_i[227];
  assign ins_o[994] = ver_i[226];
  assign ins_o[993] = ver_i[225];
  assign ins_o[992] = ver_i[224];
  assign ins_o[991] = ver_i[223];
  assign ins_o[990] = ver_i[222];
  assign ins_o[989] = ver_i[221];
  assign ins_o[988] = ver_i[220];
  assign ins_o[987] = ver_i[219];
  assign ins_o[986] = ver_i[218];
  assign ins_o[985] = ver_i[217];
  assign ins_o[984] = ver_i[216];
  assign ins_o[983] = ver_i[215];
  assign ins_o[982] = ver_i[214];
  assign ins_o[981] = ver_i[213];
  assign ins_o[980] = ver_i[212];
  assign ins_o[979] = ver_i[211];
  assign ins_o[978] = ver_i[210];
  assign ins_o[977] = ver_i[209];
  assign ins_o[976] = ver_i[208];
  assign ins_o[975] = ver_i[207];
  assign ins_o[974] = ver_i[206];
  assign ins_o[973] = ver_i[205];
  assign ins_o[972] = ver_i[204];
  assign ins_o[971] = ver_i[203];
  assign ins_o[970] = ver_i[202];
  assign ins_o[969] = ver_i[201];
  assign ins_o[968] = ver_i[200];
  assign ins_o[967] = ver_i[199];
  assign ins_o[966] = ver_i[198];
  assign ins_o[965] = ver_i[197];
  assign ins_o[964] = ver_i[196];
  assign ins_o[963] = ver_i[195];
  assign ins_o[962] = ver_i[194];
  assign ins_o[961] = ver_i[193];
  assign ins_o[960] = ver_i[192];
  assign ins_o[959] = outs_i[511];
  assign ins_o[958] = outs_i[510];
  assign ins_o[957] = outs_i[509];
  assign ins_o[956] = outs_i[508];
  assign ins_o[955] = outs_i[507];
  assign ins_o[954] = outs_i[506];
  assign ins_o[953] = outs_i[505];
  assign ins_o[952] = outs_i[504];
  assign ins_o[951] = outs_i[503];
  assign ins_o[950] = outs_i[502];
  assign ins_o[949] = outs_i[501];
  assign ins_o[948] = outs_i[500];
  assign ins_o[947] = outs_i[499];
  assign ins_o[946] = outs_i[498];
  assign ins_o[945] = outs_i[497];
  assign ins_o[944] = outs_i[496];
  assign ins_o[943] = outs_i[495];
  assign ins_o[942] = outs_i[494];
  assign ins_o[941] = outs_i[493];
  assign ins_o[940] = outs_i[492];
  assign ins_o[939] = outs_i[491];
  assign ins_o[938] = outs_i[490];
  assign ins_o[937] = outs_i[489];
  assign ins_o[936] = outs_i[488];
  assign ins_o[935] = outs_i[487];
  assign ins_o[934] = outs_i[486];
  assign ins_o[933] = outs_i[485];
  assign ins_o[932] = outs_i[484];
  assign ins_o[931] = outs_i[483];
  assign ins_o[930] = outs_i[482];
  assign ins_o[929] = outs_i[481];
  assign ins_o[928] = outs_i[480];
  assign ins_o[927] = outs_i[479];
  assign ins_o[926] = outs_i[478];
  assign ins_o[925] = outs_i[477];
  assign ins_o[924] = outs_i[476];
  assign ins_o[923] = outs_i[475];
  assign ins_o[922] = outs_i[474];
  assign ins_o[921] = outs_i[473];
  assign ins_o[920] = outs_i[472];
  assign ins_o[919] = outs_i[471];
  assign ins_o[918] = outs_i[470];
  assign ins_o[917] = outs_i[469];
  assign ins_o[916] = outs_i[468];
  assign ins_o[915] = outs_i[467];
  assign ins_o[914] = outs_i[466];
  assign ins_o[913] = outs_i[465];
  assign ins_o[912] = outs_i[464];
  assign ins_o[911] = outs_i[463];
  assign ins_o[910] = outs_i[462];
  assign ins_o[909] = outs_i[461];
  assign ins_o[908] = outs_i[460];
  assign ins_o[907] = outs_i[459];
  assign ins_o[906] = outs_i[458];
  assign ins_o[905] = outs_i[457];
  assign ins_o[904] = outs_i[456];
  assign ins_o[903] = outs_i[455];
  assign ins_o[902] = outs_i[454];
  assign ins_o[901] = outs_i[453];
  assign ins_o[900] = outs_i[452];
  assign ins_o[899] = outs_i[451];
  assign ins_o[898] = outs_i[450];
  assign ins_o[897] = outs_i[449];
  assign ins_o[896] = outs_i[448];
  assign ins_o[895] = hor_i[255];
  assign ins_o[894] = hor_i[254];
  assign ins_o[893] = hor_i[253];
  assign ins_o[892] = hor_i[252];
  assign ins_o[891] = hor_i[251];
  assign ins_o[890] = hor_i[250];
  assign ins_o[889] = hor_i[249];
  assign ins_o[888] = hor_i[248];
  assign ins_o[887] = hor_i[247];
  assign ins_o[886] = hor_i[246];
  assign ins_o[885] = hor_i[245];
  assign ins_o[884] = hor_i[244];
  assign ins_o[883] = hor_i[243];
  assign ins_o[882] = hor_i[242];
  assign ins_o[881] = hor_i[241];
  assign ins_o[880] = hor_i[240];
  assign ins_o[879] = hor_i[239];
  assign ins_o[878] = hor_i[238];
  assign ins_o[877] = hor_i[237];
  assign ins_o[876] = hor_i[236];
  assign ins_o[875] = hor_i[235];
  assign ins_o[874] = hor_i[234];
  assign ins_o[873] = hor_i[233];
  assign ins_o[872] = hor_i[232];
  assign ins_o[871] = hor_i[231];
  assign ins_o[870] = hor_i[230];
  assign ins_o[869] = hor_i[229];
  assign ins_o[868] = hor_i[228];
  assign ins_o[867] = hor_i[227];
  assign ins_o[866] = hor_i[226];
  assign ins_o[865] = hor_i[225];
  assign ins_o[864] = hor_i[224];
  assign ins_o[863] = hor_i[223];
  assign ins_o[862] = hor_i[222];
  assign ins_o[861] = hor_i[221];
  assign ins_o[860] = hor_i[220];
  assign ins_o[859] = hor_i[219];
  assign ins_o[858] = hor_i[218];
  assign ins_o[857] = hor_i[217];
  assign ins_o[856] = hor_i[216];
  assign ins_o[855] = hor_i[215];
  assign ins_o[854] = hor_i[214];
  assign ins_o[853] = hor_i[213];
  assign ins_o[852] = hor_i[212];
  assign ins_o[851] = hor_i[211];
  assign ins_o[850] = hor_i[210];
  assign ins_o[849] = hor_i[209];
  assign ins_o[848] = hor_i[208];
  assign ins_o[847] = hor_i[207];
  assign ins_o[846] = hor_i[206];
  assign ins_o[845] = hor_i[205];
  assign ins_o[844] = hor_i[204];
  assign ins_o[843] = hor_i[203];
  assign ins_o[842] = hor_i[202];
  assign ins_o[841] = hor_i[201];
  assign ins_o[840] = hor_i[200];
  assign ins_o[839] = hor_i[199];
  assign ins_o[838] = hor_i[198];
  assign ins_o[837] = hor_i[197];
  assign ins_o[836] = hor_i[196];
  assign ins_o[835] = hor_i[195];
  assign ins_o[834] = hor_i[194];
  assign ins_o[833] = hor_i[193];
  assign ins_o[832] = hor_i[192];
  assign ins_o[831] = outs_i[639];
  assign ins_o[830] = outs_i[638];
  assign ins_o[829] = outs_i[637];
  assign ins_o[828] = outs_i[636];
  assign ins_o[827] = outs_i[635];
  assign ins_o[826] = outs_i[634];
  assign ins_o[825] = outs_i[633];
  assign ins_o[824] = outs_i[632];
  assign ins_o[823] = outs_i[631];
  assign ins_o[822] = outs_i[630];
  assign ins_o[821] = outs_i[629];
  assign ins_o[820] = outs_i[628];
  assign ins_o[819] = outs_i[627];
  assign ins_o[818] = outs_i[626];
  assign ins_o[817] = outs_i[625];
  assign ins_o[816] = outs_i[624];
  assign ins_o[815] = outs_i[623];
  assign ins_o[814] = outs_i[622];
  assign ins_o[813] = outs_i[621];
  assign ins_o[812] = outs_i[620];
  assign ins_o[811] = outs_i[619];
  assign ins_o[810] = outs_i[618];
  assign ins_o[809] = outs_i[617];
  assign ins_o[808] = outs_i[616];
  assign ins_o[807] = outs_i[615];
  assign ins_o[806] = outs_i[614];
  assign ins_o[805] = outs_i[613];
  assign ins_o[804] = outs_i[612];
  assign ins_o[803] = outs_i[611];
  assign ins_o[802] = outs_i[610];
  assign ins_o[801] = outs_i[609];
  assign ins_o[800] = outs_i[608];
  assign ins_o[799] = outs_i[607];
  assign ins_o[798] = outs_i[606];
  assign ins_o[797] = outs_i[605];
  assign ins_o[796] = outs_i[604];
  assign ins_o[795] = outs_i[603];
  assign ins_o[794] = outs_i[602];
  assign ins_o[793] = outs_i[601];
  assign ins_o[792] = outs_i[600];
  assign ins_o[791] = outs_i[599];
  assign ins_o[790] = outs_i[598];
  assign ins_o[789] = outs_i[597];
  assign ins_o[788] = outs_i[596];
  assign ins_o[787] = outs_i[595];
  assign ins_o[786] = outs_i[594];
  assign ins_o[785] = outs_i[593];
  assign ins_o[784] = outs_i[592];
  assign ins_o[783] = outs_i[591];
  assign ins_o[782] = outs_i[590];
  assign ins_o[781] = outs_i[589];
  assign ins_o[780] = outs_i[588];
  assign ins_o[779] = outs_i[587];
  assign ins_o[778] = outs_i[586];
  assign ins_o[777] = outs_i[585];
  assign ins_o[776] = outs_i[584];
  assign ins_o[775] = outs_i[583];
  assign ins_o[774] = outs_i[582];
  assign ins_o[773] = outs_i[581];
  assign ins_o[772] = outs_i[580];
  assign ins_o[771] = outs_i[579];
  assign ins_o[770] = outs_i[578];
  assign ins_o[769] = outs_i[577];
  assign ins_o[768] = outs_i[576];
  assign ins_o[767] = ver_i[191];
  assign ins_o[766] = ver_i[190];
  assign ins_o[765] = ver_i[189];
  assign ins_o[764] = ver_i[188];
  assign ins_o[763] = ver_i[187];
  assign ins_o[762] = ver_i[186];
  assign ins_o[761] = ver_i[185];
  assign ins_o[760] = ver_i[184];
  assign ins_o[759] = ver_i[183];
  assign ins_o[758] = ver_i[182];
  assign ins_o[757] = ver_i[181];
  assign ins_o[756] = ver_i[180];
  assign ins_o[755] = ver_i[179];
  assign ins_o[754] = ver_i[178];
  assign ins_o[753] = ver_i[177];
  assign ins_o[752] = ver_i[176];
  assign ins_o[751] = ver_i[175];
  assign ins_o[750] = ver_i[174];
  assign ins_o[749] = ver_i[173];
  assign ins_o[748] = ver_i[172];
  assign ins_o[747] = ver_i[171];
  assign ins_o[746] = ver_i[170];
  assign ins_o[745] = ver_i[169];
  assign ins_o[744] = ver_i[168];
  assign ins_o[743] = ver_i[167];
  assign ins_o[742] = ver_i[166];
  assign ins_o[741] = ver_i[165];
  assign ins_o[740] = ver_i[164];
  assign ins_o[739] = ver_i[163];
  assign ins_o[738] = ver_i[162];
  assign ins_o[737] = ver_i[161];
  assign ins_o[736] = ver_i[160];
  assign ins_o[735] = ver_i[159];
  assign ins_o[734] = ver_i[158];
  assign ins_o[733] = ver_i[157];
  assign ins_o[732] = ver_i[156];
  assign ins_o[731] = ver_i[155];
  assign ins_o[730] = ver_i[154];
  assign ins_o[729] = ver_i[153];
  assign ins_o[728] = ver_i[152];
  assign ins_o[727] = ver_i[151];
  assign ins_o[726] = ver_i[150];
  assign ins_o[725] = ver_i[149];
  assign ins_o[724] = ver_i[148];
  assign ins_o[723] = ver_i[147];
  assign ins_o[722] = ver_i[146];
  assign ins_o[721] = ver_i[145];
  assign ins_o[720] = ver_i[144];
  assign ins_o[719] = ver_i[143];
  assign ins_o[718] = ver_i[142];
  assign ins_o[717] = ver_i[141];
  assign ins_o[716] = ver_i[140];
  assign ins_o[715] = ver_i[139];
  assign ins_o[714] = ver_i[138];
  assign ins_o[713] = ver_i[137];
  assign ins_o[712] = ver_i[136];
  assign ins_o[711] = ver_i[135];
  assign ins_o[710] = ver_i[134];
  assign ins_o[709] = ver_i[133];
  assign ins_o[708] = ver_i[132];
  assign ins_o[707] = ver_i[131];
  assign ins_o[706] = ver_i[130];
  assign ins_o[705] = ver_i[129];
  assign ins_o[704] = ver_i[128];
  assign ins_o[703] = outs_i[255];
  assign ins_o[702] = outs_i[254];
  assign ins_o[701] = outs_i[253];
  assign ins_o[700] = outs_i[252];
  assign ins_o[699] = outs_i[251];
  assign ins_o[698] = outs_i[250];
  assign ins_o[697] = outs_i[249];
  assign ins_o[696] = outs_i[248];
  assign ins_o[695] = outs_i[247];
  assign ins_o[694] = outs_i[246];
  assign ins_o[693] = outs_i[245];
  assign ins_o[692] = outs_i[244];
  assign ins_o[691] = outs_i[243];
  assign ins_o[690] = outs_i[242];
  assign ins_o[689] = outs_i[241];
  assign ins_o[688] = outs_i[240];
  assign ins_o[687] = outs_i[239];
  assign ins_o[686] = outs_i[238];
  assign ins_o[685] = outs_i[237];
  assign ins_o[684] = outs_i[236];
  assign ins_o[683] = outs_i[235];
  assign ins_o[682] = outs_i[234];
  assign ins_o[681] = outs_i[233];
  assign ins_o[680] = outs_i[232];
  assign ins_o[679] = outs_i[231];
  assign ins_o[678] = outs_i[230];
  assign ins_o[677] = outs_i[229];
  assign ins_o[676] = outs_i[228];
  assign ins_o[675] = outs_i[227];
  assign ins_o[674] = outs_i[226];
  assign ins_o[673] = outs_i[225];
  assign ins_o[672] = outs_i[224];
  assign ins_o[671] = outs_i[223];
  assign ins_o[670] = outs_i[222];
  assign ins_o[669] = outs_i[221];
  assign ins_o[668] = outs_i[220];
  assign ins_o[667] = outs_i[219];
  assign ins_o[666] = outs_i[218];
  assign ins_o[665] = outs_i[217];
  assign ins_o[664] = outs_i[216];
  assign ins_o[663] = outs_i[215];
  assign ins_o[662] = outs_i[214];
  assign ins_o[661] = outs_i[213];
  assign ins_o[660] = outs_i[212];
  assign ins_o[659] = outs_i[211];
  assign ins_o[658] = outs_i[210];
  assign ins_o[657] = outs_i[209];
  assign ins_o[656] = outs_i[208];
  assign ins_o[655] = outs_i[207];
  assign ins_o[654] = outs_i[206];
  assign ins_o[653] = outs_i[205];
  assign ins_o[652] = outs_i[204];
  assign ins_o[651] = outs_i[203];
  assign ins_o[650] = outs_i[202];
  assign ins_o[649] = outs_i[201];
  assign ins_o[648] = outs_i[200];
  assign ins_o[647] = outs_i[199];
  assign ins_o[646] = outs_i[198];
  assign ins_o[645] = outs_i[197];
  assign ins_o[644] = outs_i[196];
  assign ins_o[643] = outs_i[195];
  assign ins_o[642] = outs_i[194];
  assign ins_o[641] = outs_i[193];
  assign ins_o[640] = outs_i[192];
  assign ins_o[639] = outs_i[831];
  assign ins_o[638] = outs_i[830];
  assign ins_o[637] = outs_i[829];
  assign ins_o[636] = outs_i[828];
  assign ins_o[635] = outs_i[827];
  assign ins_o[634] = outs_i[826];
  assign ins_o[633] = outs_i[825];
  assign ins_o[632] = outs_i[824];
  assign ins_o[631] = outs_i[823];
  assign ins_o[630] = outs_i[822];
  assign ins_o[629] = outs_i[821];
  assign ins_o[628] = outs_i[820];
  assign ins_o[627] = outs_i[819];
  assign ins_o[626] = outs_i[818];
  assign ins_o[625] = outs_i[817];
  assign ins_o[624] = outs_i[816];
  assign ins_o[623] = outs_i[815];
  assign ins_o[622] = outs_i[814];
  assign ins_o[621] = outs_i[813];
  assign ins_o[620] = outs_i[812];
  assign ins_o[619] = outs_i[811];
  assign ins_o[618] = outs_i[810];
  assign ins_o[617] = outs_i[809];
  assign ins_o[616] = outs_i[808];
  assign ins_o[615] = outs_i[807];
  assign ins_o[614] = outs_i[806];
  assign ins_o[613] = outs_i[805];
  assign ins_o[612] = outs_i[804];
  assign ins_o[611] = outs_i[803];
  assign ins_o[610] = outs_i[802];
  assign ins_o[609] = outs_i[801];
  assign ins_o[608] = outs_i[800];
  assign ins_o[607] = outs_i[799];
  assign ins_o[606] = outs_i[798];
  assign ins_o[605] = outs_i[797];
  assign ins_o[604] = outs_i[796];
  assign ins_o[603] = outs_i[795];
  assign ins_o[602] = outs_i[794];
  assign ins_o[601] = outs_i[793];
  assign ins_o[600] = outs_i[792];
  assign ins_o[599] = outs_i[791];
  assign ins_o[598] = outs_i[790];
  assign ins_o[597] = outs_i[789];
  assign ins_o[596] = outs_i[788];
  assign ins_o[595] = outs_i[787];
  assign ins_o[594] = outs_i[786];
  assign ins_o[593] = outs_i[785];
  assign ins_o[592] = outs_i[784];
  assign ins_o[591] = outs_i[783];
  assign ins_o[590] = outs_i[782];
  assign ins_o[589] = outs_i[781];
  assign ins_o[588] = outs_i[780];
  assign ins_o[587] = outs_i[779];
  assign ins_o[586] = outs_i[778];
  assign ins_o[585] = outs_i[777];
  assign ins_o[584] = outs_i[776];
  assign ins_o[583] = outs_i[775];
  assign ins_o[582] = outs_i[774];
  assign ins_o[581] = outs_i[773];
  assign ins_o[580] = outs_i[772];
  assign ins_o[579] = outs_i[771];
  assign ins_o[578] = outs_i[770];
  assign ins_o[577] = outs_i[769];
  assign ins_o[576] = outs_i[768];
  assign ins_o[575] = hor_i[127];
  assign ins_o[574] = hor_i[126];
  assign ins_o[573] = hor_i[125];
  assign ins_o[572] = hor_i[124];
  assign ins_o[571] = hor_i[123];
  assign ins_o[570] = hor_i[122];
  assign ins_o[569] = hor_i[121];
  assign ins_o[568] = hor_i[120];
  assign ins_o[567] = hor_i[119];
  assign ins_o[566] = hor_i[118];
  assign ins_o[565] = hor_i[117];
  assign ins_o[564] = hor_i[116];
  assign ins_o[563] = hor_i[115];
  assign ins_o[562] = hor_i[114];
  assign ins_o[561] = hor_i[113];
  assign ins_o[560] = hor_i[112];
  assign ins_o[559] = hor_i[111];
  assign ins_o[558] = hor_i[110];
  assign ins_o[557] = hor_i[109];
  assign ins_o[556] = hor_i[108];
  assign ins_o[555] = hor_i[107];
  assign ins_o[554] = hor_i[106];
  assign ins_o[553] = hor_i[105];
  assign ins_o[552] = hor_i[104];
  assign ins_o[551] = hor_i[103];
  assign ins_o[550] = hor_i[102];
  assign ins_o[549] = hor_i[101];
  assign ins_o[548] = hor_i[100];
  assign ins_o[547] = hor_i[99];
  assign ins_o[546] = hor_i[98];
  assign ins_o[545] = hor_i[97];
  assign ins_o[544] = hor_i[96];
  assign ins_o[543] = hor_i[95];
  assign ins_o[542] = hor_i[94];
  assign ins_o[541] = hor_i[93];
  assign ins_o[540] = hor_i[92];
  assign ins_o[539] = hor_i[91];
  assign ins_o[538] = hor_i[90];
  assign ins_o[537] = hor_i[89];
  assign ins_o[536] = hor_i[88];
  assign ins_o[535] = hor_i[87];
  assign ins_o[534] = hor_i[86];
  assign ins_o[533] = hor_i[85];
  assign ins_o[532] = hor_i[84];
  assign ins_o[531] = hor_i[83];
  assign ins_o[530] = hor_i[82];
  assign ins_o[529] = hor_i[81];
  assign ins_o[528] = hor_i[80];
  assign ins_o[527] = hor_i[79];
  assign ins_o[526] = hor_i[78];
  assign ins_o[525] = hor_i[77];
  assign ins_o[524] = hor_i[76];
  assign ins_o[523] = hor_i[75];
  assign ins_o[522] = hor_i[74];
  assign ins_o[521] = hor_i[73];
  assign ins_o[520] = hor_i[72];
  assign ins_o[519] = hor_i[71];
  assign ins_o[518] = hor_i[70];
  assign ins_o[517] = hor_i[69];
  assign ins_o[516] = hor_i[68];
  assign ins_o[515] = hor_i[67];
  assign ins_o[514] = hor_i[66];
  assign ins_o[513] = hor_i[65];
  assign ins_o[512] = hor_i[64];
  assign ins_o[511] = outs_i[959];
  assign ins_o[510] = outs_i[958];
  assign ins_o[509] = outs_i[957];
  assign ins_o[508] = outs_i[956];
  assign ins_o[507] = outs_i[955];
  assign ins_o[506] = outs_i[954];
  assign ins_o[505] = outs_i[953];
  assign ins_o[504] = outs_i[952];
  assign ins_o[503] = outs_i[951];
  assign ins_o[502] = outs_i[950];
  assign ins_o[501] = outs_i[949];
  assign ins_o[500] = outs_i[948];
  assign ins_o[499] = outs_i[947];
  assign ins_o[498] = outs_i[946];
  assign ins_o[497] = outs_i[945];
  assign ins_o[496] = outs_i[944];
  assign ins_o[495] = outs_i[943];
  assign ins_o[494] = outs_i[942];
  assign ins_o[493] = outs_i[941];
  assign ins_o[492] = outs_i[940];
  assign ins_o[491] = outs_i[939];
  assign ins_o[490] = outs_i[938];
  assign ins_o[489] = outs_i[937];
  assign ins_o[488] = outs_i[936];
  assign ins_o[487] = outs_i[935];
  assign ins_o[486] = outs_i[934];
  assign ins_o[485] = outs_i[933];
  assign ins_o[484] = outs_i[932];
  assign ins_o[483] = outs_i[931];
  assign ins_o[482] = outs_i[930];
  assign ins_o[481] = outs_i[929];
  assign ins_o[480] = outs_i[928];
  assign ins_o[479] = outs_i[927];
  assign ins_o[478] = outs_i[926];
  assign ins_o[477] = outs_i[925];
  assign ins_o[476] = outs_i[924];
  assign ins_o[475] = outs_i[923];
  assign ins_o[474] = outs_i[922];
  assign ins_o[473] = outs_i[921];
  assign ins_o[472] = outs_i[920];
  assign ins_o[471] = outs_i[919];
  assign ins_o[470] = outs_i[918];
  assign ins_o[469] = outs_i[917];
  assign ins_o[468] = outs_i[916];
  assign ins_o[467] = outs_i[915];
  assign ins_o[466] = outs_i[914];
  assign ins_o[465] = outs_i[913];
  assign ins_o[464] = outs_i[912];
  assign ins_o[463] = outs_i[911];
  assign ins_o[462] = outs_i[910];
  assign ins_o[461] = outs_i[909];
  assign ins_o[460] = outs_i[908];
  assign ins_o[459] = outs_i[907];
  assign ins_o[458] = outs_i[906];
  assign ins_o[457] = outs_i[905];
  assign ins_o[456] = outs_i[904];
  assign ins_o[455] = outs_i[903];
  assign ins_o[454] = outs_i[902];
  assign ins_o[453] = outs_i[901];
  assign ins_o[452] = outs_i[900];
  assign ins_o[451] = outs_i[899];
  assign ins_o[450] = outs_i[898];
  assign ins_o[449] = outs_i[897];
  assign ins_o[448] = outs_i[896];
  assign ins_o[447] = ver_i[127];
  assign ins_o[446] = ver_i[126];
  assign ins_o[445] = ver_i[125];
  assign ins_o[444] = ver_i[124];
  assign ins_o[443] = ver_i[123];
  assign ins_o[442] = ver_i[122];
  assign ins_o[441] = ver_i[121];
  assign ins_o[440] = ver_i[120];
  assign ins_o[439] = ver_i[119];
  assign ins_o[438] = ver_i[118];
  assign ins_o[437] = ver_i[117];
  assign ins_o[436] = ver_i[116];
  assign ins_o[435] = ver_i[115];
  assign ins_o[434] = ver_i[114];
  assign ins_o[433] = ver_i[113];
  assign ins_o[432] = ver_i[112];
  assign ins_o[431] = ver_i[111];
  assign ins_o[430] = ver_i[110];
  assign ins_o[429] = ver_i[109];
  assign ins_o[428] = ver_i[108];
  assign ins_o[427] = ver_i[107];
  assign ins_o[426] = ver_i[106];
  assign ins_o[425] = ver_i[105];
  assign ins_o[424] = ver_i[104];
  assign ins_o[423] = ver_i[103];
  assign ins_o[422] = ver_i[102];
  assign ins_o[421] = ver_i[101];
  assign ins_o[420] = ver_i[100];
  assign ins_o[419] = ver_i[99];
  assign ins_o[418] = ver_i[98];
  assign ins_o[417] = ver_i[97];
  assign ins_o[416] = ver_i[96];
  assign ins_o[415] = ver_i[95];
  assign ins_o[414] = ver_i[94];
  assign ins_o[413] = ver_i[93];
  assign ins_o[412] = ver_i[92];
  assign ins_o[411] = ver_i[91];
  assign ins_o[410] = ver_i[90];
  assign ins_o[409] = ver_i[89];
  assign ins_o[408] = ver_i[88];
  assign ins_o[407] = ver_i[87];
  assign ins_o[406] = ver_i[86];
  assign ins_o[405] = ver_i[85];
  assign ins_o[404] = ver_i[84];
  assign ins_o[403] = ver_i[83];
  assign ins_o[402] = ver_i[82];
  assign ins_o[401] = ver_i[81];
  assign ins_o[400] = ver_i[80];
  assign ins_o[399] = ver_i[79];
  assign ins_o[398] = ver_i[78];
  assign ins_o[397] = ver_i[77];
  assign ins_o[396] = ver_i[76];
  assign ins_o[395] = ver_i[75];
  assign ins_o[394] = ver_i[74];
  assign ins_o[393] = ver_i[73];
  assign ins_o[392] = ver_i[72];
  assign ins_o[391] = ver_i[71];
  assign ins_o[390] = ver_i[70];
  assign ins_o[389] = ver_i[69];
  assign ins_o[388] = ver_i[68];
  assign ins_o[387] = ver_i[67];
  assign ins_o[386] = ver_i[66];
  assign ins_o[385] = ver_i[65];
  assign ins_o[384] = ver_i[64];
  assign ins_o[383] = hor_i[191];
  assign ins_o[382] = hor_i[190];
  assign ins_o[381] = hor_i[189];
  assign ins_o[380] = hor_i[188];
  assign ins_o[379] = hor_i[187];
  assign ins_o[378] = hor_i[186];
  assign ins_o[377] = hor_i[185];
  assign ins_o[376] = hor_i[184];
  assign ins_o[375] = hor_i[183];
  assign ins_o[374] = hor_i[182];
  assign ins_o[373] = hor_i[181];
  assign ins_o[372] = hor_i[180];
  assign ins_o[371] = hor_i[179];
  assign ins_o[370] = hor_i[178];
  assign ins_o[369] = hor_i[177];
  assign ins_o[368] = hor_i[176];
  assign ins_o[367] = hor_i[175];
  assign ins_o[366] = hor_i[174];
  assign ins_o[365] = hor_i[173];
  assign ins_o[364] = hor_i[172];
  assign ins_o[363] = hor_i[171];
  assign ins_o[362] = hor_i[170];
  assign ins_o[361] = hor_i[169];
  assign ins_o[360] = hor_i[168];
  assign ins_o[359] = hor_i[167];
  assign ins_o[358] = hor_i[166];
  assign ins_o[357] = hor_i[165];
  assign ins_o[356] = hor_i[164];
  assign ins_o[355] = hor_i[163];
  assign ins_o[354] = hor_i[162];
  assign ins_o[353] = hor_i[161];
  assign ins_o[352] = hor_i[160];
  assign ins_o[351] = hor_i[159];
  assign ins_o[350] = hor_i[158];
  assign ins_o[349] = hor_i[157];
  assign ins_o[348] = hor_i[156];
  assign ins_o[347] = hor_i[155];
  assign ins_o[346] = hor_i[154];
  assign ins_o[345] = hor_i[153];
  assign ins_o[344] = hor_i[152];
  assign ins_o[343] = hor_i[151];
  assign ins_o[342] = hor_i[150];
  assign ins_o[341] = hor_i[149];
  assign ins_o[340] = hor_i[148];
  assign ins_o[339] = hor_i[147];
  assign ins_o[338] = hor_i[146];
  assign ins_o[337] = hor_i[145];
  assign ins_o[336] = hor_i[144];
  assign ins_o[335] = hor_i[143];
  assign ins_o[334] = hor_i[142];
  assign ins_o[333] = hor_i[141];
  assign ins_o[332] = hor_i[140];
  assign ins_o[331] = hor_i[139];
  assign ins_o[330] = hor_i[138];
  assign ins_o[329] = hor_i[137];
  assign ins_o[328] = hor_i[136];
  assign ins_o[327] = hor_i[135];
  assign ins_o[326] = hor_i[134];
  assign ins_o[325] = hor_i[133];
  assign ins_o[324] = hor_i[132];
  assign ins_o[323] = hor_i[131];
  assign ins_o[322] = hor_i[130];
  assign ins_o[321] = hor_i[129];
  assign ins_o[320] = hor_i[128];
  assign ins_o[319] = outs_i[127];
  assign ins_o[318] = outs_i[126];
  assign ins_o[317] = outs_i[125];
  assign ins_o[316] = outs_i[124];
  assign ins_o[315] = outs_i[123];
  assign ins_o[314] = outs_i[122];
  assign ins_o[313] = outs_i[121];
  assign ins_o[312] = outs_i[120];
  assign ins_o[311] = outs_i[119];
  assign ins_o[310] = outs_i[118];
  assign ins_o[309] = outs_i[117];
  assign ins_o[308] = outs_i[116];
  assign ins_o[307] = outs_i[115];
  assign ins_o[306] = outs_i[114];
  assign ins_o[305] = outs_i[113];
  assign ins_o[304] = outs_i[112];
  assign ins_o[303] = outs_i[111];
  assign ins_o[302] = outs_i[110];
  assign ins_o[301] = outs_i[109];
  assign ins_o[300] = outs_i[108];
  assign ins_o[299] = outs_i[107];
  assign ins_o[298] = outs_i[106];
  assign ins_o[297] = outs_i[105];
  assign ins_o[296] = outs_i[104];
  assign ins_o[295] = outs_i[103];
  assign ins_o[294] = outs_i[102];
  assign ins_o[293] = outs_i[101];
  assign ins_o[292] = outs_i[100];
  assign ins_o[291] = outs_i[99];
  assign ins_o[290] = outs_i[98];
  assign ins_o[289] = outs_i[97];
  assign ins_o[288] = outs_i[96];
  assign ins_o[287] = outs_i[95];
  assign ins_o[286] = outs_i[94];
  assign ins_o[285] = outs_i[93];
  assign ins_o[284] = outs_i[92];
  assign ins_o[283] = outs_i[91];
  assign ins_o[282] = outs_i[90];
  assign ins_o[281] = outs_i[89];
  assign ins_o[280] = outs_i[88];
  assign ins_o[279] = outs_i[87];
  assign ins_o[278] = outs_i[86];
  assign ins_o[277] = outs_i[85];
  assign ins_o[276] = outs_i[84];
  assign ins_o[275] = outs_i[83];
  assign ins_o[274] = outs_i[82];
  assign ins_o[273] = outs_i[81];
  assign ins_o[272] = outs_i[80];
  assign ins_o[271] = outs_i[79];
  assign ins_o[270] = outs_i[78];
  assign ins_o[269] = outs_i[77];
  assign ins_o[268] = outs_i[76];
  assign ins_o[267] = outs_i[75];
  assign ins_o[266] = outs_i[74];
  assign ins_o[265] = outs_i[73];
  assign ins_o[264] = outs_i[72];
  assign ins_o[263] = outs_i[71];
  assign ins_o[262] = outs_i[70];
  assign ins_o[261] = outs_i[69];
  assign ins_o[260] = outs_i[68];
  assign ins_o[259] = outs_i[67];
  assign ins_o[258] = outs_i[66];
  assign ins_o[257] = outs_i[65];
  assign ins_o[256] = outs_i[64];
  assign ins_o[255] = outs_i[703];
  assign ins_o[254] = outs_i[702];
  assign ins_o[253] = outs_i[701];
  assign ins_o[252] = outs_i[700];
  assign ins_o[251] = outs_i[699];
  assign ins_o[250] = outs_i[698];
  assign ins_o[249] = outs_i[697];
  assign ins_o[248] = outs_i[696];
  assign ins_o[247] = outs_i[695];
  assign ins_o[246] = outs_i[694];
  assign ins_o[245] = outs_i[693];
  assign ins_o[244] = outs_i[692];
  assign ins_o[243] = outs_i[691];
  assign ins_o[242] = outs_i[690];
  assign ins_o[241] = outs_i[689];
  assign ins_o[240] = outs_i[688];
  assign ins_o[239] = outs_i[687];
  assign ins_o[238] = outs_i[686];
  assign ins_o[237] = outs_i[685];
  assign ins_o[236] = outs_i[684];
  assign ins_o[235] = outs_i[683];
  assign ins_o[234] = outs_i[682];
  assign ins_o[233] = outs_i[681];
  assign ins_o[232] = outs_i[680];
  assign ins_o[231] = outs_i[679];
  assign ins_o[230] = outs_i[678];
  assign ins_o[229] = outs_i[677];
  assign ins_o[228] = outs_i[676];
  assign ins_o[227] = outs_i[675];
  assign ins_o[226] = outs_i[674];
  assign ins_o[225] = outs_i[673];
  assign ins_o[224] = outs_i[672];
  assign ins_o[223] = outs_i[671];
  assign ins_o[222] = outs_i[670];
  assign ins_o[221] = outs_i[669];
  assign ins_o[220] = outs_i[668];
  assign ins_o[219] = outs_i[667];
  assign ins_o[218] = outs_i[666];
  assign ins_o[217] = outs_i[665];
  assign ins_o[216] = outs_i[664];
  assign ins_o[215] = outs_i[663];
  assign ins_o[214] = outs_i[662];
  assign ins_o[213] = outs_i[661];
  assign ins_o[212] = outs_i[660];
  assign ins_o[211] = outs_i[659];
  assign ins_o[210] = outs_i[658];
  assign ins_o[209] = outs_i[657];
  assign ins_o[208] = outs_i[656];
  assign ins_o[207] = outs_i[655];
  assign ins_o[206] = outs_i[654];
  assign ins_o[205] = outs_i[653];
  assign ins_o[204] = outs_i[652];
  assign ins_o[203] = outs_i[651];
  assign ins_o[202] = outs_i[650];
  assign ins_o[201] = outs_i[649];
  assign ins_o[200] = outs_i[648];
  assign ins_o[199] = outs_i[647];
  assign ins_o[198] = outs_i[646];
  assign ins_o[197] = outs_i[645];
  assign ins_o[196] = outs_i[644];
  assign ins_o[195] = outs_i[643];
  assign ins_o[194] = outs_i[642];
  assign ins_o[193] = outs_i[641];
  assign ins_o[192] = outs_i[640];
  assign ins_o[191] = ver_i[63];
  assign ins_o[190] = ver_i[62];
  assign ins_o[189] = ver_i[61];
  assign ins_o[188] = ver_i[60];
  assign ins_o[187] = ver_i[59];
  assign ins_o[186] = ver_i[58];
  assign ins_o[185] = ver_i[57];
  assign ins_o[184] = ver_i[56];
  assign ins_o[183] = ver_i[55];
  assign ins_o[182] = ver_i[54];
  assign ins_o[181] = ver_i[53];
  assign ins_o[180] = ver_i[52];
  assign ins_o[179] = ver_i[51];
  assign ins_o[178] = ver_i[50];
  assign ins_o[177] = ver_i[49];
  assign ins_o[176] = ver_i[48];
  assign ins_o[175] = ver_i[47];
  assign ins_o[174] = ver_i[46];
  assign ins_o[173] = ver_i[45];
  assign ins_o[172] = ver_i[44];
  assign ins_o[171] = ver_i[43];
  assign ins_o[170] = ver_i[42];
  assign ins_o[169] = ver_i[41];
  assign ins_o[168] = ver_i[40];
  assign ins_o[167] = ver_i[39];
  assign ins_o[166] = ver_i[38];
  assign ins_o[165] = ver_i[37];
  assign ins_o[164] = ver_i[36];
  assign ins_o[163] = ver_i[35];
  assign ins_o[162] = ver_i[34];
  assign ins_o[161] = ver_i[33];
  assign ins_o[160] = ver_i[32];
  assign ins_o[159] = ver_i[31];
  assign ins_o[158] = ver_i[30];
  assign ins_o[157] = ver_i[29];
  assign ins_o[156] = ver_i[28];
  assign ins_o[155] = ver_i[27];
  assign ins_o[154] = ver_i[26];
  assign ins_o[153] = ver_i[25];
  assign ins_o[152] = ver_i[24];
  assign ins_o[151] = ver_i[23];
  assign ins_o[150] = ver_i[22];
  assign ins_o[149] = ver_i[21];
  assign ins_o[148] = ver_i[20];
  assign ins_o[147] = ver_i[19];
  assign ins_o[146] = ver_i[18];
  assign ins_o[145] = ver_i[17];
  assign ins_o[144] = ver_i[16];
  assign ins_o[143] = ver_i[15];
  assign ins_o[142] = ver_i[14];
  assign ins_o[141] = ver_i[13];
  assign ins_o[140] = ver_i[12];
  assign ins_o[139] = ver_i[11];
  assign ins_o[138] = ver_i[10];
  assign ins_o[137] = ver_i[9];
  assign ins_o[136] = ver_i[8];
  assign ins_o[135] = ver_i[7];
  assign ins_o[134] = ver_i[6];
  assign ins_o[133] = ver_i[5];
  assign ins_o[132] = ver_i[4];
  assign ins_o[131] = ver_i[3];
  assign ins_o[130] = ver_i[2];
  assign ins_o[129] = ver_i[1];
  assign ins_o[128] = ver_i[0];
  assign ins_o[127] = outs_i[319];
  assign ins_o[126] = outs_i[318];
  assign ins_o[125] = outs_i[317];
  assign ins_o[124] = outs_i[316];
  assign ins_o[123] = outs_i[315];
  assign ins_o[122] = outs_i[314];
  assign ins_o[121] = outs_i[313];
  assign ins_o[120] = outs_i[312];
  assign ins_o[119] = outs_i[311];
  assign ins_o[118] = outs_i[310];
  assign ins_o[117] = outs_i[309];
  assign ins_o[116] = outs_i[308];
  assign ins_o[115] = outs_i[307];
  assign ins_o[114] = outs_i[306];
  assign ins_o[113] = outs_i[305];
  assign ins_o[112] = outs_i[304];
  assign ins_o[111] = outs_i[303];
  assign ins_o[110] = outs_i[302];
  assign ins_o[109] = outs_i[301];
  assign ins_o[108] = outs_i[300];
  assign ins_o[107] = outs_i[299];
  assign ins_o[106] = outs_i[298];
  assign ins_o[105] = outs_i[297];
  assign ins_o[104] = outs_i[296];
  assign ins_o[103] = outs_i[295];
  assign ins_o[102] = outs_i[294];
  assign ins_o[101] = outs_i[293];
  assign ins_o[100] = outs_i[292];
  assign ins_o[99] = outs_i[291];
  assign ins_o[98] = outs_i[290];
  assign ins_o[97] = outs_i[289];
  assign ins_o[96] = outs_i[288];
  assign ins_o[95] = outs_i[287];
  assign ins_o[94] = outs_i[286];
  assign ins_o[93] = outs_i[285];
  assign ins_o[92] = outs_i[284];
  assign ins_o[91] = outs_i[283];
  assign ins_o[90] = outs_i[282];
  assign ins_o[89] = outs_i[281];
  assign ins_o[88] = outs_i[280];
  assign ins_o[87] = outs_i[279];
  assign ins_o[86] = outs_i[278];
  assign ins_o[85] = outs_i[277];
  assign ins_o[84] = outs_i[276];
  assign ins_o[83] = outs_i[275];
  assign ins_o[82] = outs_i[274];
  assign ins_o[81] = outs_i[273];
  assign ins_o[80] = outs_i[272];
  assign ins_o[79] = outs_i[271];
  assign ins_o[78] = outs_i[270];
  assign ins_o[77] = outs_i[269];
  assign ins_o[76] = outs_i[268];
  assign ins_o[75] = outs_i[267];
  assign ins_o[74] = outs_i[266];
  assign ins_o[73] = outs_i[265];
  assign ins_o[72] = outs_i[264];
  assign ins_o[71] = outs_i[263];
  assign ins_o[70] = outs_i[262];
  assign ins_o[69] = outs_i[261];
  assign ins_o[68] = outs_i[260];
  assign ins_o[67] = outs_i[259];
  assign ins_o[66] = outs_i[258];
  assign ins_o[65] = outs_i[257];
  assign ins_o[64] = outs_i[256];
  assign ins_o[63] = hor_i[63];
  assign ins_o[62] = hor_i[62];
  assign ins_o[61] = hor_i[61];
  assign ins_o[60] = hor_i[60];
  assign ins_o[59] = hor_i[59];
  assign ins_o[58] = hor_i[58];
  assign ins_o[57] = hor_i[57];
  assign ins_o[56] = hor_i[56];
  assign ins_o[55] = hor_i[55];
  assign ins_o[54] = hor_i[54];
  assign ins_o[53] = hor_i[53];
  assign ins_o[52] = hor_i[52];
  assign ins_o[51] = hor_i[51];
  assign ins_o[50] = hor_i[50];
  assign ins_o[49] = hor_i[49];
  assign ins_o[48] = hor_i[48];
  assign ins_o[47] = hor_i[47];
  assign ins_o[46] = hor_i[46];
  assign ins_o[45] = hor_i[45];
  assign ins_o[44] = hor_i[44];
  assign ins_o[43] = hor_i[43];
  assign ins_o[42] = hor_i[42];
  assign ins_o[41] = hor_i[41];
  assign ins_o[40] = hor_i[40];
  assign ins_o[39] = hor_i[39];
  assign ins_o[38] = hor_i[38];
  assign ins_o[37] = hor_i[37];
  assign ins_o[36] = hor_i[36];
  assign ins_o[35] = hor_i[35];
  assign ins_o[34] = hor_i[34];
  assign ins_o[33] = hor_i[33];
  assign ins_o[32] = hor_i[32];
  assign ins_o[31] = hor_i[31];
  assign ins_o[30] = hor_i[30];
  assign ins_o[29] = hor_i[29];
  assign ins_o[28] = hor_i[28];
  assign ins_o[27] = hor_i[27];
  assign ins_o[26] = hor_i[26];
  assign ins_o[25] = hor_i[25];
  assign ins_o[24] = hor_i[24];
  assign ins_o[23] = hor_i[23];
  assign ins_o[22] = hor_i[22];
  assign ins_o[21] = hor_i[21];
  assign ins_o[20] = hor_i[20];
  assign ins_o[19] = hor_i[19];
  assign ins_o[18] = hor_i[18];
  assign ins_o[17] = hor_i[17];
  assign ins_o[16] = hor_i[16];
  assign ins_o[15] = hor_i[15];
  assign ins_o[14] = hor_i[14];
  assign ins_o[13] = hor_i[13];
  assign ins_o[12] = hor_i[12];
  assign ins_o[11] = hor_i[11];
  assign ins_o[10] = hor_i[10];
  assign ins_o[9] = hor_i[9];
  assign ins_o[8] = hor_i[8];
  assign ins_o[7] = hor_i[7];
  assign ins_o[6] = hor_i[6];
  assign ins_o[5] = hor_i[5];
  assign ins_o[4] = hor_i[4];
  assign ins_o[3] = hor_i[3];
  assign ins_o[2] = hor_i[2];
  assign ins_o[1] = hor_i[1];
  assign ins_o[0] = hor_i[0];
  assign hor_o[255] = outs_i[895];
  assign hor_o[254] = outs_i[894];
  assign hor_o[253] = outs_i[893];
  assign hor_o[252] = outs_i[892];
  assign hor_o[251] = outs_i[891];
  assign hor_o[250] = outs_i[890];
  assign hor_o[249] = outs_i[889];
  assign hor_o[248] = outs_i[888];
  assign hor_o[247] = outs_i[887];
  assign hor_o[246] = outs_i[886];
  assign hor_o[245] = outs_i[885];
  assign hor_o[244] = outs_i[884];
  assign hor_o[243] = outs_i[883];
  assign hor_o[242] = outs_i[882];
  assign hor_o[241] = outs_i[881];
  assign hor_o[240] = outs_i[880];
  assign hor_o[239] = outs_i[879];
  assign hor_o[238] = outs_i[878];
  assign hor_o[237] = outs_i[877];
  assign hor_o[236] = outs_i[876];
  assign hor_o[235] = outs_i[875];
  assign hor_o[234] = outs_i[874];
  assign hor_o[233] = outs_i[873];
  assign hor_o[232] = outs_i[872];
  assign hor_o[231] = outs_i[871];
  assign hor_o[230] = outs_i[870];
  assign hor_o[229] = outs_i[869];
  assign hor_o[228] = outs_i[868];
  assign hor_o[227] = outs_i[867];
  assign hor_o[226] = outs_i[866];
  assign hor_o[225] = outs_i[865];
  assign hor_o[224] = outs_i[864];
  assign hor_o[223] = outs_i[863];
  assign hor_o[222] = outs_i[862];
  assign hor_o[221] = outs_i[861];
  assign hor_o[220] = outs_i[860];
  assign hor_o[219] = outs_i[859];
  assign hor_o[218] = outs_i[858];
  assign hor_o[217] = outs_i[857];
  assign hor_o[216] = outs_i[856];
  assign hor_o[215] = outs_i[855];
  assign hor_o[214] = outs_i[854];
  assign hor_o[213] = outs_i[853];
  assign hor_o[212] = outs_i[852];
  assign hor_o[211] = outs_i[851];
  assign hor_o[210] = outs_i[850];
  assign hor_o[209] = outs_i[849];
  assign hor_o[208] = outs_i[848];
  assign hor_o[207] = outs_i[847];
  assign hor_o[206] = outs_i[846];
  assign hor_o[205] = outs_i[845];
  assign hor_o[204] = outs_i[844];
  assign hor_o[203] = outs_i[843];
  assign hor_o[202] = outs_i[842];
  assign hor_o[201] = outs_i[841];
  assign hor_o[200] = outs_i[840];
  assign hor_o[199] = outs_i[839];
  assign hor_o[198] = outs_i[838];
  assign hor_o[197] = outs_i[837];
  assign hor_o[196] = outs_i[836];
  assign hor_o[195] = outs_i[835];
  assign hor_o[194] = outs_i[834];
  assign hor_o[193] = outs_i[833];
  assign hor_o[192] = outs_i[832];
  assign hor_o[191] = outs_i[383];
  assign hor_o[190] = outs_i[382];
  assign hor_o[189] = outs_i[381];
  assign hor_o[188] = outs_i[380];
  assign hor_o[187] = outs_i[379];
  assign hor_o[186] = outs_i[378];
  assign hor_o[185] = outs_i[377];
  assign hor_o[184] = outs_i[376];
  assign hor_o[183] = outs_i[375];
  assign hor_o[182] = outs_i[374];
  assign hor_o[181] = outs_i[373];
  assign hor_o[180] = outs_i[372];
  assign hor_o[179] = outs_i[371];
  assign hor_o[178] = outs_i[370];
  assign hor_o[177] = outs_i[369];
  assign hor_o[176] = outs_i[368];
  assign hor_o[175] = outs_i[367];
  assign hor_o[174] = outs_i[366];
  assign hor_o[173] = outs_i[365];
  assign hor_o[172] = outs_i[364];
  assign hor_o[171] = outs_i[363];
  assign hor_o[170] = outs_i[362];
  assign hor_o[169] = outs_i[361];
  assign hor_o[168] = outs_i[360];
  assign hor_o[167] = outs_i[359];
  assign hor_o[166] = outs_i[358];
  assign hor_o[165] = outs_i[357];
  assign hor_o[164] = outs_i[356];
  assign hor_o[163] = outs_i[355];
  assign hor_o[162] = outs_i[354];
  assign hor_o[161] = outs_i[353];
  assign hor_o[160] = outs_i[352];
  assign hor_o[159] = outs_i[351];
  assign hor_o[158] = outs_i[350];
  assign hor_o[157] = outs_i[349];
  assign hor_o[156] = outs_i[348];
  assign hor_o[155] = outs_i[347];
  assign hor_o[154] = outs_i[346];
  assign hor_o[153] = outs_i[345];
  assign hor_o[152] = outs_i[344];
  assign hor_o[151] = outs_i[343];
  assign hor_o[150] = outs_i[342];
  assign hor_o[149] = outs_i[341];
  assign hor_o[148] = outs_i[340];
  assign hor_o[147] = outs_i[339];
  assign hor_o[146] = outs_i[338];
  assign hor_o[145] = outs_i[337];
  assign hor_o[144] = outs_i[336];
  assign hor_o[143] = outs_i[335];
  assign hor_o[142] = outs_i[334];
  assign hor_o[141] = outs_i[333];
  assign hor_o[140] = outs_i[332];
  assign hor_o[139] = outs_i[331];
  assign hor_o[138] = outs_i[330];
  assign hor_o[137] = outs_i[329];
  assign hor_o[136] = outs_i[328];
  assign hor_o[135] = outs_i[327];
  assign hor_o[134] = outs_i[326];
  assign hor_o[133] = outs_i[325];
  assign hor_o[132] = outs_i[324];
  assign hor_o[131] = outs_i[323];
  assign hor_o[130] = outs_i[322];
  assign hor_o[129] = outs_i[321];
  assign hor_o[128] = outs_i[320];
  assign hor_o[127] = outs_i[575];
  assign hor_o[126] = outs_i[574];
  assign hor_o[125] = outs_i[573];
  assign hor_o[124] = outs_i[572];
  assign hor_o[123] = outs_i[571];
  assign hor_o[122] = outs_i[570];
  assign hor_o[121] = outs_i[569];
  assign hor_o[120] = outs_i[568];
  assign hor_o[119] = outs_i[567];
  assign hor_o[118] = outs_i[566];
  assign hor_o[117] = outs_i[565];
  assign hor_o[116] = outs_i[564];
  assign hor_o[115] = outs_i[563];
  assign hor_o[114] = outs_i[562];
  assign hor_o[113] = outs_i[561];
  assign hor_o[112] = outs_i[560];
  assign hor_o[111] = outs_i[559];
  assign hor_o[110] = outs_i[558];
  assign hor_o[109] = outs_i[557];
  assign hor_o[108] = outs_i[556];
  assign hor_o[107] = outs_i[555];
  assign hor_o[106] = outs_i[554];
  assign hor_o[105] = outs_i[553];
  assign hor_o[104] = outs_i[552];
  assign hor_o[103] = outs_i[551];
  assign hor_o[102] = outs_i[550];
  assign hor_o[101] = outs_i[549];
  assign hor_o[100] = outs_i[548];
  assign hor_o[99] = outs_i[547];
  assign hor_o[98] = outs_i[546];
  assign hor_o[97] = outs_i[545];
  assign hor_o[96] = outs_i[544];
  assign hor_o[95] = outs_i[543];
  assign hor_o[94] = outs_i[542];
  assign hor_o[93] = outs_i[541];
  assign hor_o[92] = outs_i[540];
  assign hor_o[91] = outs_i[539];
  assign hor_o[90] = outs_i[538];
  assign hor_o[89] = outs_i[537];
  assign hor_o[88] = outs_i[536];
  assign hor_o[87] = outs_i[535];
  assign hor_o[86] = outs_i[534];
  assign hor_o[85] = outs_i[533];
  assign hor_o[84] = outs_i[532];
  assign hor_o[83] = outs_i[531];
  assign hor_o[82] = outs_i[530];
  assign hor_o[81] = outs_i[529];
  assign hor_o[80] = outs_i[528];
  assign hor_o[79] = outs_i[527];
  assign hor_o[78] = outs_i[526];
  assign hor_o[77] = outs_i[525];
  assign hor_o[76] = outs_i[524];
  assign hor_o[75] = outs_i[523];
  assign hor_o[74] = outs_i[522];
  assign hor_o[73] = outs_i[521];
  assign hor_o[72] = outs_i[520];
  assign hor_o[71] = outs_i[519];
  assign hor_o[70] = outs_i[518];
  assign hor_o[69] = outs_i[517];
  assign hor_o[68] = outs_i[516];
  assign hor_o[67] = outs_i[515];
  assign hor_o[66] = outs_i[514];
  assign hor_o[65] = outs_i[513];
  assign hor_o[64] = outs_i[512];
  assign hor_o[63] = outs_i[63];
  assign hor_o[62] = outs_i[62];
  assign hor_o[61] = outs_i[61];
  assign hor_o[60] = outs_i[60];
  assign hor_o[59] = outs_i[59];
  assign hor_o[58] = outs_i[58];
  assign hor_o[57] = outs_i[57];
  assign hor_o[56] = outs_i[56];
  assign hor_o[55] = outs_i[55];
  assign hor_o[54] = outs_i[54];
  assign hor_o[53] = outs_i[53];
  assign hor_o[52] = outs_i[52];
  assign hor_o[51] = outs_i[51];
  assign hor_o[50] = outs_i[50];
  assign hor_o[49] = outs_i[49];
  assign hor_o[48] = outs_i[48];
  assign hor_o[47] = outs_i[47];
  assign hor_o[46] = outs_i[46];
  assign hor_o[45] = outs_i[45];
  assign hor_o[44] = outs_i[44];
  assign hor_o[43] = outs_i[43];
  assign hor_o[42] = outs_i[42];
  assign hor_o[41] = outs_i[41];
  assign hor_o[40] = outs_i[40];
  assign hor_o[39] = outs_i[39];
  assign hor_o[38] = outs_i[38];
  assign hor_o[37] = outs_i[37];
  assign hor_o[36] = outs_i[36];
  assign hor_o[35] = outs_i[35];
  assign hor_o[34] = outs_i[34];
  assign hor_o[33] = outs_i[33];
  assign hor_o[32] = outs_i[32];
  assign hor_o[31] = outs_i[31];
  assign hor_o[30] = outs_i[30];
  assign hor_o[29] = outs_i[29];
  assign hor_o[28] = outs_i[28];
  assign hor_o[27] = outs_i[27];
  assign hor_o[26] = outs_i[26];
  assign hor_o[25] = outs_i[25];
  assign hor_o[24] = outs_i[24];
  assign hor_o[23] = outs_i[23];
  assign hor_o[22] = outs_i[22];
  assign hor_o[21] = outs_i[21];
  assign hor_o[20] = outs_i[20];
  assign hor_o[19] = outs_i[19];
  assign hor_o[18] = outs_i[18];
  assign hor_o[17] = outs_i[17];
  assign hor_o[16] = outs_i[16];
  assign hor_o[15] = outs_i[15];
  assign hor_o[14] = outs_i[14];
  assign hor_o[13] = outs_i[13];
  assign hor_o[12] = outs_i[12];
  assign hor_o[11] = outs_i[11];
  assign hor_o[10] = outs_i[10];
  assign hor_o[9] = outs_i[9];
  assign hor_o[8] = outs_i[8];
  assign hor_o[7] = outs_i[7];
  assign hor_o[6] = outs_i[6];
  assign hor_o[5] = outs_i[5];
  assign hor_o[4] = outs_i[4];
  assign hor_o[3] = outs_i[3];
  assign hor_o[2] = outs_i[2];
  assign hor_o[1] = outs_i[1];
  assign hor_o[0] = outs_i[0];
  assign ver_o[255] = outs_i[1023];
  assign ver_o[254] = outs_i[1022];
  assign ver_o[253] = outs_i[1021];
  assign ver_o[252] = outs_i[1020];
  assign ver_o[251] = outs_i[1019];
  assign ver_o[250] = outs_i[1018];
  assign ver_o[249] = outs_i[1017];
  assign ver_o[248] = outs_i[1016];
  assign ver_o[247] = outs_i[1015];
  assign ver_o[246] = outs_i[1014];
  assign ver_o[245] = outs_i[1013];
  assign ver_o[244] = outs_i[1012];
  assign ver_o[243] = outs_i[1011];
  assign ver_o[242] = outs_i[1010];
  assign ver_o[241] = outs_i[1009];
  assign ver_o[240] = outs_i[1008];
  assign ver_o[239] = outs_i[1007];
  assign ver_o[238] = outs_i[1006];
  assign ver_o[237] = outs_i[1005];
  assign ver_o[236] = outs_i[1004];
  assign ver_o[235] = outs_i[1003];
  assign ver_o[234] = outs_i[1002];
  assign ver_o[233] = outs_i[1001];
  assign ver_o[232] = outs_i[1000];
  assign ver_o[231] = outs_i[999];
  assign ver_o[230] = outs_i[998];
  assign ver_o[229] = outs_i[997];
  assign ver_o[228] = outs_i[996];
  assign ver_o[227] = outs_i[995];
  assign ver_o[226] = outs_i[994];
  assign ver_o[225] = outs_i[993];
  assign ver_o[224] = outs_i[992];
  assign ver_o[223] = outs_i[991];
  assign ver_o[222] = outs_i[990];
  assign ver_o[221] = outs_i[989];
  assign ver_o[220] = outs_i[988];
  assign ver_o[219] = outs_i[987];
  assign ver_o[218] = outs_i[986];
  assign ver_o[217] = outs_i[985];
  assign ver_o[216] = outs_i[984];
  assign ver_o[215] = outs_i[983];
  assign ver_o[214] = outs_i[982];
  assign ver_o[213] = outs_i[981];
  assign ver_o[212] = outs_i[980];
  assign ver_o[211] = outs_i[979];
  assign ver_o[210] = outs_i[978];
  assign ver_o[209] = outs_i[977];
  assign ver_o[208] = outs_i[976];
  assign ver_o[207] = outs_i[975];
  assign ver_o[206] = outs_i[974];
  assign ver_o[205] = outs_i[973];
  assign ver_o[204] = outs_i[972];
  assign ver_o[203] = outs_i[971];
  assign ver_o[202] = outs_i[970];
  assign ver_o[201] = outs_i[969];
  assign ver_o[200] = outs_i[968];
  assign ver_o[199] = outs_i[967];
  assign ver_o[198] = outs_i[966];
  assign ver_o[197] = outs_i[965];
  assign ver_o[196] = outs_i[964];
  assign ver_o[195] = outs_i[963];
  assign ver_o[194] = outs_i[962];
  assign ver_o[193] = outs_i[961];
  assign ver_o[192] = outs_i[960];
  assign ver_o[191] = outs_i[767];
  assign ver_o[190] = outs_i[766];
  assign ver_o[189] = outs_i[765];
  assign ver_o[188] = outs_i[764];
  assign ver_o[187] = outs_i[763];
  assign ver_o[186] = outs_i[762];
  assign ver_o[185] = outs_i[761];
  assign ver_o[184] = outs_i[760];
  assign ver_o[183] = outs_i[759];
  assign ver_o[182] = outs_i[758];
  assign ver_o[181] = outs_i[757];
  assign ver_o[180] = outs_i[756];
  assign ver_o[179] = outs_i[755];
  assign ver_o[178] = outs_i[754];
  assign ver_o[177] = outs_i[753];
  assign ver_o[176] = outs_i[752];
  assign ver_o[175] = outs_i[751];
  assign ver_o[174] = outs_i[750];
  assign ver_o[173] = outs_i[749];
  assign ver_o[172] = outs_i[748];
  assign ver_o[171] = outs_i[747];
  assign ver_o[170] = outs_i[746];
  assign ver_o[169] = outs_i[745];
  assign ver_o[168] = outs_i[744];
  assign ver_o[167] = outs_i[743];
  assign ver_o[166] = outs_i[742];
  assign ver_o[165] = outs_i[741];
  assign ver_o[164] = outs_i[740];
  assign ver_o[163] = outs_i[739];
  assign ver_o[162] = outs_i[738];
  assign ver_o[161] = outs_i[737];
  assign ver_o[160] = outs_i[736];
  assign ver_o[159] = outs_i[735];
  assign ver_o[158] = outs_i[734];
  assign ver_o[157] = outs_i[733];
  assign ver_o[156] = outs_i[732];
  assign ver_o[155] = outs_i[731];
  assign ver_o[154] = outs_i[730];
  assign ver_o[153] = outs_i[729];
  assign ver_o[152] = outs_i[728];
  assign ver_o[151] = outs_i[727];
  assign ver_o[150] = outs_i[726];
  assign ver_o[149] = outs_i[725];
  assign ver_o[148] = outs_i[724];
  assign ver_o[147] = outs_i[723];
  assign ver_o[146] = outs_i[722];
  assign ver_o[145] = outs_i[721];
  assign ver_o[144] = outs_i[720];
  assign ver_o[143] = outs_i[719];
  assign ver_o[142] = outs_i[718];
  assign ver_o[141] = outs_i[717];
  assign ver_o[140] = outs_i[716];
  assign ver_o[139] = outs_i[715];
  assign ver_o[138] = outs_i[714];
  assign ver_o[137] = outs_i[713];
  assign ver_o[136] = outs_i[712];
  assign ver_o[135] = outs_i[711];
  assign ver_o[134] = outs_i[710];
  assign ver_o[133] = outs_i[709];
  assign ver_o[132] = outs_i[708];
  assign ver_o[131] = outs_i[707];
  assign ver_o[130] = outs_i[706];
  assign ver_o[129] = outs_i[705];
  assign ver_o[128] = outs_i[704];
  assign ver_o[127] = outs_i[447];
  assign ver_o[126] = outs_i[446];
  assign ver_o[125] = outs_i[445];
  assign ver_o[124] = outs_i[444];
  assign ver_o[123] = outs_i[443];
  assign ver_o[122] = outs_i[442];
  assign ver_o[121] = outs_i[441];
  assign ver_o[120] = outs_i[440];
  assign ver_o[119] = outs_i[439];
  assign ver_o[118] = outs_i[438];
  assign ver_o[117] = outs_i[437];
  assign ver_o[116] = outs_i[436];
  assign ver_o[115] = outs_i[435];
  assign ver_o[114] = outs_i[434];
  assign ver_o[113] = outs_i[433];
  assign ver_o[112] = outs_i[432];
  assign ver_o[111] = outs_i[431];
  assign ver_o[110] = outs_i[430];
  assign ver_o[109] = outs_i[429];
  assign ver_o[108] = outs_i[428];
  assign ver_o[107] = outs_i[427];
  assign ver_o[106] = outs_i[426];
  assign ver_o[105] = outs_i[425];
  assign ver_o[104] = outs_i[424];
  assign ver_o[103] = outs_i[423];
  assign ver_o[102] = outs_i[422];
  assign ver_o[101] = outs_i[421];
  assign ver_o[100] = outs_i[420];
  assign ver_o[99] = outs_i[419];
  assign ver_o[98] = outs_i[418];
  assign ver_o[97] = outs_i[417];
  assign ver_o[96] = outs_i[416];
  assign ver_o[95] = outs_i[415];
  assign ver_o[94] = outs_i[414];
  assign ver_o[93] = outs_i[413];
  assign ver_o[92] = outs_i[412];
  assign ver_o[91] = outs_i[411];
  assign ver_o[90] = outs_i[410];
  assign ver_o[89] = outs_i[409];
  assign ver_o[88] = outs_i[408];
  assign ver_o[87] = outs_i[407];
  assign ver_o[86] = outs_i[406];
  assign ver_o[85] = outs_i[405];
  assign ver_o[84] = outs_i[404];
  assign ver_o[83] = outs_i[403];
  assign ver_o[82] = outs_i[402];
  assign ver_o[81] = outs_i[401];
  assign ver_o[80] = outs_i[400];
  assign ver_o[79] = outs_i[399];
  assign ver_o[78] = outs_i[398];
  assign ver_o[77] = outs_i[397];
  assign ver_o[76] = outs_i[396];
  assign ver_o[75] = outs_i[395];
  assign ver_o[74] = outs_i[394];
  assign ver_o[73] = outs_i[393];
  assign ver_o[72] = outs_i[392];
  assign ver_o[71] = outs_i[391];
  assign ver_o[70] = outs_i[390];
  assign ver_o[69] = outs_i[389];
  assign ver_o[68] = outs_i[388];
  assign ver_o[67] = outs_i[387];
  assign ver_o[66] = outs_i[386];
  assign ver_o[65] = outs_i[385];
  assign ver_o[64] = outs_i[384];
  assign ver_o[63] = outs_i[191];
  assign ver_o[62] = outs_i[190];
  assign ver_o[61] = outs_i[189];
  assign ver_o[60] = outs_i[188];
  assign ver_o[59] = outs_i[187];
  assign ver_o[58] = outs_i[186];
  assign ver_o[57] = outs_i[185];
  assign ver_o[56] = outs_i[184];
  assign ver_o[55] = outs_i[183];
  assign ver_o[54] = outs_i[182];
  assign ver_o[53] = outs_i[181];
  assign ver_o[52] = outs_i[180];
  assign ver_o[51] = outs_i[179];
  assign ver_o[50] = outs_i[178];
  assign ver_o[49] = outs_i[177];
  assign ver_o[48] = outs_i[176];
  assign ver_o[47] = outs_i[175];
  assign ver_o[46] = outs_i[174];
  assign ver_o[45] = outs_i[173];
  assign ver_o[44] = outs_i[172];
  assign ver_o[43] = outs_i[171];
  assign ver_o[42] = outs_i[170];
  assign ver_o[41] = outs_i[169];
  assign ver_o[40] = outs_i[168];
  assign ver_o[39] = outs_i[167];
  assign ver_o[38] = outs_i[166];
  assign ver_o[37] = outs_i[165];
  assign ver_o[36] = outs_i[164];
  assign ver_o[35] = outs_i[163];
  assign ver_o[34] = outs_i[162];
  assign ver_o[33] = outs_i[161];
  assign ver_o[32] = outs_i[160];
  assign ver_o[31] = outs_i[159];
  assign ver_o[30] = outs_i[158];
  assign ver_o[29] = outs_i[157];
  assign ver_o[28] = outs_i[156];
  assign ver_o[27] = outs_i[155];
  assign ver_o[26] = outs_i[154];
  assign ver_o[25] = outs_i[153];
  assign ver_o[24] = outs_i[152];
  assign ver_o[23] = outs_i[151];
  assign ver_o[22] = outs_i[150];
  assign ver_o[21] = outs_i[149];
  assign ver_o[20] = outs_i[148];
  assign ver_o[19] = outs_i[147];
  assign ver_o[18] = outs_i[146];
  assign ver_o[17] = outs_i[145];
  assign ver_o[16] = outs_i[144];
  assign ver_o[15] = outs_i[143];
  assign ver_o[14] = outs_i[142];
  assign ver_o[13] = outs_i[141];
  assign ver_o[12] = outs_i[140];
  assign ver_o[11] = outs_i[139];
  assign ver_o[10] = outs_i[138];
  assign ver_o[9] = outs_i[137];
  assign ver_o[8] = outs_i[136];
  assign ver_o[7] = outs_i[135];
  assign ver_o[6] = outs_i[134];
  assign ver_o[5] = outs_i[133];
  assign ver_o[4] = outs_i[132];
  assign ver_o[3] = outs_i[131];
  assign ver_o[2] = outs_i[130];
  assign ver_o[1] = outs_i[129];
  assign ver_o[0] = outs_i[128];

endmodule