module TLXbar_9( // @[:freechips.rocketchip.system.TinyConfig.fir@102674.2]
  output        auto_in_a_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input         auto_in_a_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [2:0]  auto_in_a_bits_opcode, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [2:0]  auto_in_a_bits_param, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [2:0]  auto_in_a_bits_size, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [4:0]  auto_in_a_bits_source, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [31:0] auto_in_a_bits_address, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [3:0]  auto_in_a_bits_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [31:0] auto_in_a_bits_data, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input         auto_in_d_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output        auto_in_d_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [2:0]  auto_in_d_bits_opcode, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [2:0]  auto_in_d_bits_size, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [4:0]  auto_in_d_bits_source, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [31:0] auto_in_d_bits_data, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input         auto_out_a_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output        auto_out_a_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [2:0]  auto_out_a_bits_opcode, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [2:0]  auto_out_a_bits_param, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [2:0]  auto_out_a_bits_size, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [4:0]  auto_out_a_bits_source, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [31:0] auto_out_a_bits_address, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [3:0]  auto_out_a_bits_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output [31:0] auto_out_a_bits_data, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  output        auto_out_d_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input         auto_out_d_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [2:0]  auto_out_d_bits_opcode, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [2:0]  auto_out_d_bits_size, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [4:0]  auto_out_d_bits_source, // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
  input  [31:0] auto_out_d_bits_data // @[:freechips.rocketchip.system.TinyConfig.fir@102677.4]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[LazyModule.scala 173:31:freechips.rocketchip.system.TinyConfig.fir@102687.4]
  assign auto_in_d_valid = auto_out_d_valid; // @[LazyModule.scala 173:31:freechips.rocketchip.system.TinyConfig.fir@102687.4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[LazyModule.scala 173:31:freechips.rocketchip.system.TinyConfig.fir@102687.4]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[LazyModule.scala 173:31:freechips.rocketchip.system.TinyConfig.fir@102687.4]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[LazyModule.scala 173:31:freechips.rocketchip.system.TinyConfig.fir@102687.4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[LazyModule.scala 173:31:freechips.rocketchip.system.TinyConfig.fir@102687.4]
  assign auto_out_a_valid = auto_in_a_valid; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
  assign auto_out_d_ready = auto_in_d_ready; // @[LazyModule.scala 173:49:freechips.rocketchip.system.TinyConfig.fir@102686.4]
endmodule