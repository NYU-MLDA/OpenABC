module ifu_compress_ctl
(
  din,
  dout,
  legal
);

  input [15:0] din;
  output [31:0] dout;
  output legal;
  wire [31:0] dout;
  wire legal,l1_30,rdrd,rdprd,rs2prd,rdeq1,rdeq2,rdrs1,rdprs1,rs1eq2,rs2rs2,rs2prs2,
  simm5_0,uimm9_2,simm9_4,ulwimm6_2,ulwspimm7_2,uimm5_0,sjaloffset11_1,sluimm17_12,
  sbroffset8_1,uswimm6_2,uswspimm7_2,l3_11,l3_10,l3_9,l3_8,l3_7,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,
  N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,
  N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,
  N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,
  N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,
  N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,
  N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,
  N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,
  N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,
  N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,
  N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,
  N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,
  N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,
  N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,
  N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,
  N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,
  N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
  N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,
  N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,
  N746,N747;
  wire [24:2] l1;
  wire [20:20] o;
  wire [31:12] l2;
  wire [31:25] l3;
  assign l1[11] = N14 | N15;
  assign N14 = N12 | N13;
  assign N12 = 1'b0 | N11;
  assign N11 = rdrd & din[11];
  assign N13 = rdprd & 1'b0;
  assign N15 = rs2prd & 1'b0;
  assign l1[10] = N19 | N20;
  assign N19 = N17 | N18;
  assign N17 = 1'b0 | N16;
  assign N16 = rdrd & din[10];
  assign N18 = rdprd & 1'b1;
  assign N20 = rs2prd & 1'b1;
  assign l1[9] = N24 | N25;
  assign N24 = N22 | N23;
  assign N22 = 1'b0 | N21;
  assign N21 = rdrd & din[9];
  assign N23 = rdprd & din[9];
  assign N25 = rs2prd & din[4];
  assign l1[8] = N31 | rdeq2;
  assign N31 = N29 | N30;
  assign N29 = N27 | N28;
  assign N27 = 1'b0 | N26;
  assign N26 = rdrd & din[8];
  assign N28 = rdprd & din[8];
  assign N30 = rs2prd & din[3];
  assign l1[7] = N37 | rdeq1;
  assign N37 = N35 | N36;
  assign N35 = N33 | N34;
  assign N33 = 1'b0 | N32;
  assign N32 = rdrd & din[7];
  assign N34 = rdprd & din[7];
  assign N36 = rs2prd & din[2];
  assign l1[19] = N39 | N40;
  assign N39 = 1'b0 | N38;
  assign N38 = rdrs1 & din[11];
  assign N40 = rdprs1 & 1'b0;
  assign l1[18] = N42 | N43;
  assign N42 = 1'b0 | N41;
  assign N41 = rdrs1 & din[10];
  assign N43 = rdprs1 & 1'b1;
  assign l1[17] = N45 | N46;
  assign N45 = 1'b0 | N44;
  assign N44 = rdrs1 & din[9];
  assign N46 = rdprs1 & din[9];
  assign l1[16] = N50 | rs1eq2;
  assign N50 = N48 | N49;
  assign N48 = 1'b0 | N47;
  assign N47 = rdrs1 & din[8];
  assign N49 = rdprs1 & din[8];
  assign l1[15] = N52 | N53;
  assign N52 = 1'b0 | N51;
  assign N51 = rdrs1 & din[7];
  assign N53 = rdprs1 & din[7];
  assign l1[24] = N55 | N56;
  assign N55 = 1'b0 | N54;
  assign N54 = rs2rs2 & din[6];
  assign N56 = rs2prs2 & 1'b0;
  assign l1[23] = N58 | N59;
  assign N58 = 1'b0 | N57;
  assign N57 = rs2rs2 & din[5];
  assign N59 = rs2prs2 & 1'b1;
  assign l1[22] = N61 | N62;
  assign N61 = 1'b0 | N60;
  assign N60 = rs2rs2 & din[4];
  assign N62 = rs2prs2 & din[4];
  assign l1[21] = N64 | N65;
  assign N64 = 1'b0 | N63;
  assign N63 = rs2rs2 & din[3];
  assign N65 = rs2prs2 & din[3];
  assign l1[20] = N67 | N68;
  assign N67 = o[20] | N66;
  assign N66 = rs2rs2 & din[2];
  assign N68 = rs2prs2 & din[2];
  assign l2[31] = N74 | N75;
  assign N74 = N72 | N73;
  assign N72 = N70 | N71;
  assign N70 = 1'b0 | N69;
  assign N69 = simm5_0 & din[12];
  assign N71 = simm9_4 & din[12];
  assign N73 = sjaloffset11_1 & din[12];
  assign N75 = sluimm17_12 & din[12];
  assign l2[30] = N81 | N82;
  assign N81 = N79 | N80;
  assign N79 = N77 | N78;
  assign N77 = l1_30 | N76;
  assign N76 = simm5_0 & din[12];
  assign N78 = simm9_4 & din[12];
  assign N80 = sjaloffset11_1 & din[8];
  assign N82 = sluimm17_12 & din[12];
  assign l2[29] = N90 | N91;
  assign N90 = N88 | N89;
  assign N88 = N86 | N87;
  assign N86 = N84 | N85;
  assign N84 = 1'b0 | N83;
  assign N83 = simm5_0 & din[12];
  assign N85 = uimm9_2 & din[10];
  assign N87 = simm9_4 & din[12];
  assign N89 = sjaloffset11_1 & din[10];
  assign N91 = sluimm17_12 & din[12];
  assign l2[28] = N99 | N100;
  assign N99 = N97 | N98;
  assign N97 = N95 | N96;
  assign N95 = N93 | N94;
  assign N93 = 1'b0 | N92;
  assign N92 = simm5_0 & din[12];
  assign N94 = uimm9_2 & din[9];
  assign N96 = simm9_4 & din[4];
  assign N98 = sjaloffset11_1 & din[9];
  assign N100 = sluimm17_12 & din[12];
  assign l2[27] = N110 | N111;
  assign N110 = N108 | N109;
  assign N108 = N106 | N107;
  assign N106 = N104 | N105;
  assign N104 = N102 | N103;
  assign N102 = 1'b0 | N101;
  assign N101 = simm5_0 & din[12];
  assign N103 = uimm9_2 & din[8];
  assign N105 = simm9_4 & din[3];
  assign N107 = ulwspimm7_2 & din[3];
  assign N109 = sjaloffset11_1 & din[6];
  assign N111 = sluimm17_12 & din[12];
  assign l2[26] = N123 | N124;
  assign N123 = N121 | N122;
  assign N121 = N119 | N120;
  assign N119 = N117 | N118;
  assign N117 = N115 | N116;
  assign N115 = N113 | N114;
  assign N113 = 1'b0 | N112;
  assign N112 = simm5_0 & din[12];
  assign N114 = uimm9_2 & din[7];
  assign N116 = simm9_4 & din[5];
  assign N118 = ulwimm6_2 & din[5];
  assign N120 = ulwspimm7_2 & din[2];
  assign N122 = sjaloffset11_1 & din[7];
  assign N124 = sluimm17_12 & din[12];
  assign l2[25] = N138 | N139;
  assign N138 = N136 | N137;
  assign N136 = N134 | N135;
  assign N134 = N132 | N133;
  assign N132 = N130 | N131;
  assign N130 = N128 | N129;
  assign N128 = N126 | N127;
  assign N126 = 1'b0 | N125;
  assign N125 = simm5_0 & din[12];
  assign N127 = uimm9_2 & din[12];
  assign N129 = simm9_4 & din[2];
  assign N131 = ulwimm6_2 & din[12];
  assign N133 = ulwspimm7_2 & din[12];
  assign N135 = uimm5_0 & din[12];
  assign N137 = sjaloffset11_1 & din[2];
  assign N139 = sluimm17_12 & din[12];
  assign l2[24] = N153 | N154;
  assign N153 = N151 | N152;
  assign N151 = N149 | N150;
  assign N149 = N147 | N148;
  assign N147 = N145 | N146;
  assign N145 = N143 | N144;
  assign N143 = N141 | N142;
  assign N141 = l1[24] | N140;
  assign N140 = simm5_0 & din[6];
  assign N142 = uimm9_2 & din[11];
  assign N144 = simm9_4 & din[6];
  assign N146 = ulwimm6_2 & din[11];
  assign N148 = ulwspimm7_2 & din[6];
  assign N150 = uimm5_0 & din[6];
  assign N152 = sjaloffset11_1 & din[11];
  assign N154 = sluimm17_12 & din[12];
  assign l2[23] = N166 | N167;
  assign N166 = N164 | N165;
  assign N164 = N162 | N163;
  assign N162 = N160 | N161;
  assign N160 = N158 | N159;
  assign N158 = N156 | N157;
  assign N156 = l1[23] | N155;
  assign N155 = simm5_0 & din[5];
  assign N157 = uimm9_2 & din[5];
  assign N159 = ulwimm6_2 & din[10];
  assign N161 = ulwspimm7_2 & din[5];
  assign N163 = uimm5_0 & din[5];
  assign N165 = sjaloffset11_1 & din[5];
  assign N167 = sluimm17_12 & din[12];
  assign l2[22] = N179 | N180;
  assign N179 = N177 | N178;
  assign N177 = N175 | N176;
  assign N175 = N173 | N174;
  assign N173 = N171 | N172;
  assign N171 = N169 | N170;
  assign N169 = l1[22] | N168;
  assign N168 = simm5_0 & din[4];
  assign N170 = uimm9_2 & din[6];
  assign N172 = ulwimm6_2 & din[6];
  assign N174 = ulwspimm7_2 & din[4];
  assign N176 = uimm5_0 & din[4];
  assign N178 = sjaloffset11_1 & din[4];
  assign N180 = sluimm17_12 & din[12];
  assign l2[21] = N186 | N187;
  assign N186 = N184 | N185;
  assign N184 = N182 | N183;
  assign N182 = l1[21] | N181;
  assign N181 = simm5_0 & din[3];
  assign N183 = uimm5_0 & din[3];
  assign N185 = sjaloffset11_1 & din[3];
  assign N187 = sluimm17_12 & din[12];
  assign l2[20] = N193 | N194;
  assign N193 = N191 | N192;
  assign N191 = N189 | N190;
  assign N189 = l1[20] | N188;
  assign N188 = simm5_0 & din[2];
  assign N190 = uimm5_0 & din[2];
  assign N192 = sjaloffset11_1 & din[12];
  assign N194 = sluimm17_12 & din[12];
  assign l2[19] = N196 | N197;
  assign N196 = l1[19] | N195;
  assign N195 = sjaloffset11_1 & din[12];
  assign N197 = sluimm17_12 & din[12];
  assign l2[18] = N199 | N200;
  assign N199 = l1[18] | N198;
  assign N198 = sjaloffset11_1 & din[12];
  assign N200 = sluimm17_12 & din[12];
  assign l2[17] = N202 | N203;
  assign N202 = l1[17] | N201;
  assign N201 = sjaloffset11_1 & din[12];
  assign N203 = sluimm17_12 & din[12];
  assign l2[16] = N205 | N206;
  assign N205 = l1[16] | N204;
  assign N204 = sjaloffset11_1 & din[12];
  assign N206 = sluimm17_12 & din[6];
  assign l2[15] = N208 | N209;
  assign N208 = l1[15] | N207;
  assign N207 = sjaloffset11_1 & din[12];
  assign N209 = sluimm17_12 & din[5];
  assign l2[14] = N211 | N212;
  assign N211 = l1[14] | N210;
  assign N210 = sjaloffset11_1 & din[12];
  assign N212 = sluimm17_12 & din[4];
  assign l2[13] = N214 | N215;
  assign N214 = l1[13] | N213;
  assign N213 = sjaloffset11_1 & din[12];
  assign N215 = sluimm17_12 & din[3];
  assign l2[12] = N217 | N218;
  assign N217 = l1[12] | N216;
  assign N216 = sjaloffset11_1 & din[12];
  assign N218 = sluimm17_12 & din[2];
  assign l3[31] = l2[31] | N219;
  assign N219 = sbroffset8_1 & din[12];
  assign l3[30] = l2[30] | N220;
  assign N220 = sbroffset8_1 & din[12];
  assign l3[29] = l2[29] | N221;
  assign N221 = sbroffset8_1 & din[12];
  assign l3[28] = l2[28] | N222;
  assign N222 = sbroffset8_1 & din[12];
  assign l3[27] = N224 | N225;
  assign N224 = l2[27] | N223;
  assign N223 = sbroffset8_1 & din[6];
  assign N225 = uswspimm7_2 & din[8];
  assign l3[26] = N229 | N230;
  assign N229 = N227 | N228;
  assign N227 = l2[26] | N226;
  assign N226 = sbroffset8_1 & din[5];
  assign N228 = uswimm6_2 & din[5];
  assign N230 = uswspimm7_2 & din[7];
  assign l3[25] = N234 | N235;
  assign N234 = N232 | N233;
  assign N232 = l2[25] | N231;
  assign N231 = sbroffset8_1 & din[2];
  assign N233 = uswimm6_2 & din[12];
  assign N235 = uswspimm7_2 & din[12];
  assign l3_11 = N239 | N240;
  assign N239 = N237 | N238;
  assign N237 = l1[11] | N236;
  assign N236 = sbroffset8_1 & din[11];
  assign N238 = uswimm6_2 & din[11];
  assign N240 = uswspimm7_2 & din[11];
  assign l3_10 = N244 | N245;
  assign N244 = N242 | N243;
  assign N242 = l1[10] | N241;
  assign N241 = sbroffset8_1 & din[10];
  assign N243 = uswimm6_2 & din[10];
  assign N245 = uswspimm7_2 & din[10];
  assign l3_9 = N249 | N250;
  assign N249 = N247 | N248;
  assign N247 = l1[9] | N246;
  assign N246 = sbroffset8_1 & din[4];
  assign N248 = uswimm6_2 & din[6];
  assign N250 = uswspimm7_2 & din[9];
  assign l3_8 = l1[8] | N251;
  assign N251 = sbroffset8_1 & din[3];
  assign l3_7 = l1[7] | N252;
  assign N252 = sbroffset8_1 & din[12];
  assign dout[31] = l3[31] & legal;
  assign dout[30] = l3[30] & legal;
  assign dout[29] = l3[29] & legal;
  assign dout[28] = l3[28] & legal;
  assign dout[27] = l3[27] & legal;
  assign dout[26] = l3[26] & legal;
  assign dout[25] = l3[25] & legal;
  assign dout[24] = l2[24] & legal;
  assign dout[23] = l2[23] & legal;
  assign dout[22] = l2[22] & legal;
  assign dout[21] = l2[21] & legal;
  assign dout[20] = l2[20] & legal;
  assign dout[19] = l2[19] & legal;
  assign dout[18] = l2[18] & legal;
  assign dout[17] = l2[17] & legal;
  assign dout[16] = l2[16] & legal;
  assign dout[15] = l2[15] & legal;
  assign dout[14] = l2[14] & legal;
  assign dout[13] = l2[13] & legal;
  assign dout[12] = l2[12] & legal;
  assign dout[11] = l3_11 & legal;
  assign dout[10] = l3_10 & legal;
  assign dout[9] = l3_9 & legal;
  assign dout[8] = l3_8 & legal;
  assign dout[7] = l3_7 & legal;
  assign dout[6] = l1[6] & legal;
  assign dout[5] = l1[5] & legal;
  assign dout[4] = l1[4] & legal;
  assign dout[3] = l1[3] & legal;
  assign dout[2] = l1[2] & legal;
  assign dout[1] = 1'b1 & legal;
  assign dout[0] = 1'b1 & legal;
  assign N0 = N288 & din[14];
  assign rdrd = N284 | N287;
  assign N284 = N282 | N283;
  assign N282 = N279 | N281;
  assign N279 = N276 | N278;
  assign N276 = N272 | N275;
  assign N272 = N269 | N271;
  assign N269 = N266 | N268;
  assign N266 = N263 | N265;
  assign N263 = N260 | N262;
  assign N260 = N257 | N259;
  assign N257 = N254 | N256;
  assign N254 = N253 & din[1];
  assign N253 = N352 & din[6];
  assign N256 = N255 & din[0];
  assign N255 = N0 & din[11];
  assign N259 = N258 & din[1];
  assign N258 = N352 & din[5];
  assign N262 = N261 & din[0];
  assign N261 = N0 & din[10];
  assign N265 = N264 & din[1];
  assign N264 = N352 & din[4];
  assign N268 = N267 & din[0];
  assign N267 = N0 & din[9];
  assign N271 = N270 & din[1];
  assign N270 = N352 & din[3];
  assign N275 = N274 & din[0];
  assign N274 = N0 & N273;
  assign N273 = ~din[8];
  assign N278 = N277 & din[1];
  assign N277 = N352 & din[2];
  assign N281 = N280 & din[0];
  assign N280 = N0 & din[7];
  assign N283 = N288 & din[1];
  assign N287 = N286 & din[0];
  assign N286 = N288 & N285;
  assign N285 = ~din[13];
  assign N1 = N288 & N352;
  assign N288 = ~din[15];
  assign rdrs1 = N334 | N335;
  assign N334 = N331 | N333;
  assign N331 = N328 | N330;
  assign N328 = N325 | N327;
  assign N325 = N322 | N324;
  assign N322 = N319 | N321;
  assign N319 = N316 | N318;
  assign N316 = N302 | N315;
  assign N302 = N299 | N301;
  assign N299 = N296 | N298;
  assign N296 = N293 | N295;
  assign N293 = N290 | N292;
  assign N290 = N289 & din[1];
  assign N289 = N6 & din[11];
  assign N292 = N291 & din[1];
  assign N291 = N6 & din[10];
  assign N295 = N294 & din[1];
  assign N294 = N6 & din[9];
  assign N298 = N297 & din[1];
  assign N297 = N6 & din[8];
  assign N301 = N300 & din[1];
  assign N300 = N6 & din[7];
  assign N315 = N314 & din[1];
  assign N314 = N312 & N313;
  assign N312 = N310 & N311;
  assign N310 = N308 & N309;
  assign N308 = N306 & N307;
  assign N306 = N304 & N305;
  assign N304 = N352 & N303;
  assign N303 = ~din[12];
  assign N305 = ~din[6];
  assign N307 = ~din[5];
  assign N309 = ~din[4];
  assign N311 = ~din[3];
  assign N313 = ~din[2];
  assign N318 = N317 & din[1];
  assign N317 = N6 & din[6];
  assign N321 = N320 & din[1];
  assign N320 = N6 & din[5];
  assign N324 = N323 & din[1];
  assign N323 = N6 & din[4];
  assign N327 = N326 & din[1];
  assign N326 = N6 & din[3];
  assign N330 = N329 & din[1];
  assign N329 = N6 & din[2];
  assign N333 = N332 & din[0];
  assign N332 = N1 & N285;
  assign N335 = N1 & din[1];
  assign rs2rs2 = N349 | N351;
  assign N349 = N346 | N348;
  assign N346 = N343 | N345;
  assign N343 = N340 | N342;
  assign N340 = N337 | N339;
  assign N337 = N336 & din[1];
  assign N336 = din[15] & din[6];
  assign N339 = N338 & din[1];
  assign N338 = din[15] & din[5];
  assign N342 = N341 & din[1];
  assign N341 = din[15] & din[4];
  assign N345 = N344 & din[1];
  assign N344 = din[15] & din[3];
  assign N348 = N347 & din[1];
  assign N347 = din[15] & din[2];
  assign N351 = N350 & din[1];
  assign N350 = din[15] & din[14];
  assign rdprd = N354 & din[0];
  assign N354 = N353 & N285;
  assign N353 = din[15] & N352;
  assign N352 = ~din[14];
  assign rdprs1 = N359 | N363;
  assign N359 = N356 | N358;
  assign N356 = N355 & din[0];
  assign N355 = din[15] & N285;
  assign N358 = N357 & din[0];
  assign N357 = din[15] & din[14];
  assign N363 = N361 & N362;
  assign N361 = din[14] & N360;
  assign N360 = ~din[1];
  assign N362 = ~din[0];
  assign rs2prs2 = N368 | N370;
  assign N368 = N367 & din[0];
  assign N367 = N366 & din[10];
  assign N366 = N365 & din[11];
  assign N365 = N364 & N285;
  assign N364 = din[15] & N352;
  assign N370 = N369 & N362;
  assign N369 = din[15] & N360;
  assign rs2prd = N371 & N362;
  assign N371 = N288 & N360;
  assign uimm9_2 = N372 & N362;
  assign N372 = N352 & N360;
  assign ulwimm6_2 = N374 & N362;
  assign N374 = N373 & N360;
  assign N373 = N288 & din[14];
  assign ulwspimm7_2 = N375 & din[1];
  assign N375 = N288 & din[14];
  assign rdeq2 = N384 & N385;
  assign N384 = N383 & din[8];
  assign N383 = N381 & N382;
  assign N381 = N379 & N380;
  assign N379 = N377 & N378;
  assign N377 = N376 & din[13];
  assign N376 = N288 & din[14];
  assign N378 = ~din[11];
  assign N380 = ~din[10];
  assign N382 = ~din[9];
  assign N385 = ~din[7];
  assign rdeq1 = N424 | N426;
  assign N424 = N416 | N423;
  assign N416 = N408 | N415;
  assign N408 = N400 | N407;
  assign N400 = N392 | N399;
  assign N392 = N391 & din[1];
  assign N391 = N390 & N313;
  assign N390 = N389 & N311;
  assign N389 = N388 & N309;
  assign N388 = N387 & N307;
  assign N387 = N386 & N305;
  assign N386 = N6 & din[11];
  assign N399 = N398 & din[1];
  assign N398 = N397 & N313;
  assign N397 = N396 & N311;
  assign N396 = N395 & N309;
  assign N395 = N394 & N307;
  assign N394 = N393 & N305;
  assign N393 = N6 & din[10];
  assign N407 = N406 & din[1];
  assign N406 = N405 & N313;
  assign N405 = N404 & N311;
  assign N404 = N403 & N309;
  assign N403 = N402 & N307;
  assign N402 = N401 & N305;
  assign N401 = N6 & din[9];
  assign N415 = N414 & din[1];
  assign N414 = N413 & N313;
  assign N413 = N412 & N311;
  assign N412 = N411 & N309;
  assign N411 = N410 & N307;
  assign N410 = N409 & N305;
  assign N409 = N6 & din[8];
  assign N423 = N422 & din[1];
  assign N422 = N421 & N313;
  assign N421 = N420 & N311;
  assign N420 = N419 & N309;
  assign N419 = N418 & N307;
  assign N418 = N417 & N305;
  assign N417 = N6 & din[7];
  assign N426 = N425 & din[13];
  assign N425 = N288 & N352;
  assign rs1eq2 = N435 | N437;
  assign N435 = N433 | N434;
  assign N433 = N432 & N385;
  assign N432 = N431 & din[8];
  assign N431 = N430 & N382;
  assign N430 = N429 & N380;
  assign N429 = N428 & N378;
  assign N428 = N427 & din[13];
  assign N427 = N288 & din[14];
  assign N434 = din[14] & din[1];
  assign N437 = N436 & N362;
  assign N436 = N352 & N360;
  assign sbroffset8_1 = N438 & din[0];
  assign N438 = din[15] & din[14];
  assign simm9_4 = N444 & N385;
  assign N444 = N443 & din[8];
  assign N443 = N442 & N382;
  assign N442 = N441 & N380;
  assign N441 = N440 & N378;
  assign N440 = N439 & din[13];
  assign N439 = N288 & din[14];
  assign simm5_0 = N448 | N450;
  assign N448 = N447 & din[0];
  assign N447 = N446 & N380;
  assign N446 = N445 & din[11];
  assign N445 = N352 & N285;
  assign N450 = N449 & din[0];
  assign N449 = N288 & N285;
  assign sjaloffset11_1 = N352 & din[13];
  assign N2 = N451 & din[13];
  assign N451 = N288 & din[14];
  assign sluimm17_12 = N458 | N459;
  assign N458 = N456 | N457;
  assign N456 = N454 | N455;
  assign N454 = N452 | N453;
  assign N452 = N2 & din[7];
  assign N453 = N2 & N273;
  assign N455 = N2 & din[9];
  assign N457 = N2 & din[10];
  assign N459 = N2 & din[11];
  assign uimm5_0 = N463 | N465;
  assign N463 = N462 & din[0];
  assign N462 = N461 & N378;
  assign N461 = N460 & N285;
  assign N460 = din[15] & N352;
  assign N465 = N464 & din[1];
  assign N464 = N288 & N352;
  assign uswimm6_2 = N466 & N362;
  assign N466 = din[15] & N360;
  assign uswspimm7_2 = N467 & din[1];
  assign N467 = din[15] & din[14];
  assign l1_30 = N471 | N474;
  assign N471 = N470 & din[0];
  assign N470 = N469 & N307;
  assign N469 = N468 & N305;
  assign N468 = N3 & din[10];
  assign N474 = N473 & din[0];
  assign N473 = N472 & din[10];
  assign N472 = N3 & N378;
  assign o[20] = N485 & din[1];
  assign N485 = N484 & N313;
  assign N484 = N483 & N311;
  assign N483 = N482 & N309;
  assign N482 = N481 & N307;
  assign N481 = N480 & N305;
  assign N480 = N479 & N385;
  assign N479 = N478 & N273;
  assign N478 = N477 & N382;
  assign N477 = N476 & N380;
  assign N476 = N475 & N378;
  assign N475 = N352 & din[12];
  assign N3 = N486 & N285;
  assign N486 = din[15] & N352;
  assign l1[14] = N494 | N496;
  assign N494 = N491 | N493;
  assign N491 = N488 | N490;
  assign N488 = N487 & din[0];
  assign N487 = N3 & N378;
  assign N490 = N489 & din[0];
  assign N489 = N3 & N380;
  assign N493 = N492 & din[0];
  assign N492 = N3 & din[6];
  assign N496 = N495 & din[0];
  assign N495 = N3 & din[5];
  assign N4 = N498 & din[11];
  assign N498 = N497 & N285;
  assign N497 = din[15] & N352;
  assign l1[13] = N503 | N504;
  assign N503 = N500 | N502;
  assign N500 = N499 & din[0];
  assign N499 = N4 & N380;
  assign N502 = N501 & din[0];
  assign N501 = N4 & din[6];
  assign N504 = din[14] & N362;
  assign N5 = N505 & N285;
  assign N505 = din[15] & N352;
  assign l1[12] = N517 | N519;
  assign N517 = N514 | N516;
  assign N514 = N511 | N513;
  assign N511 = N508 | N510;
  assign N508 = N507 & din[0];
  assign N507 = N506 & din[5];
  assign N506 = N5 & din[6];
  assign N510 = N509 & din[0];
  assign N509 = N5 & N378;
  assign N513 = N512 & din[0];
  assign N512 = N5 & N380;
  assign N516 = N515 & din[1];
  assign N515 = N288 & N352;
  assign N519 = N518 & din[13];
  assign N518 = din[15] & din[14];
  assign l1[6] = N528 | N530;
  assign N528 = N526 | N527;
  assign N526 = N525 & N362;
  assign N525 = N524 & N313;
  assign N524 = N523 & N311;
  assign N523 = N522 & N309;
  assign N522 = N521 & N307;
  assign N521 = N520 & N305;
  assign N520 = din[15] & N352;
  assign N527 = N352 & din[13];
  assign N530 = N529 & din[0];
  assign N529 = din[15] & din[14];
  assign l1[5] = N546 | N547;
  assign N546 = N544 | N545;
  assign N544 = N542 | N543;
  assign N542 = N540 | N541;
  assign N540 = N538 | N539;
  assign N538 = N536 | N537;
  assign N536 = N534 | N535;
  assign N534 = N531 | N533;
  assign N531 = din[15] & N362;
  assign N533 = N532 & din[10];
  assign N532 = din[15] & din[11];
  assign N535 = din[13] & N273;
  assign N537 = din[13] & din[7];
  assign N539 = din[13] & din[9];
  assign N541 = din[13] & din[10];
  assign N543 = din[13] & din[11];
  assign N545 = N352 & din[13];
  assign N547 = din[15] & din[14];
  assign l1[4] = N574 | N576;
  assign N574 = N571 | N573;
  assign N571 = N568 | N570;
  assign N568 = N565 | N567;
  assign N565 = N562 | N564;
  assign N562 = N559 | N561;
  assign N559 = N556 | N558;
  assign N556 = N553 | N555;
  assign N553 = N552 & N362;
  assign N552 = N551 & N385;
  assign N551 = N550 & N273;
  assign N550 = N549 & N382;
  assign N549 = N548 & N380;
  assign N548 = N352 & N378;
  assign N555 = N554 & N362;
  assign N554 = N288 & N352;
  assign N558 = N557 & N362;
  assign N557 = N352 & din[6];
  assign N561 = N560 & din[0];
  assign N560 = N288 & din[14];
  assign N564 = N563 & N362;
  assign N563 = N352 & din[5];
  assign N567 = N566 & N362;
  assign N566 = N352 & din[4];
  assign N570 = N569 & din[0];
  assign N569 = N352 & N285;
  assign N573 = N572 & N362;
  assign N572 = N352 & din[3];
  assign N576 = N575 & N362;
  assign N575 = N352 & din[2];
  assign l1[3] = N352 & din[13];
  assign N6 = N352 & din[12];
  assign N7 = N288 & din[13];
  assign l1[2] = N634 | N635;
  assign N634 = N632 | N633;
  assign N632 = N630 | N631;
  assign N630 = N628 | N629;
  assign N628 = N626 | N627;
  assign N626 = N624 | N625;
  assign N624 = N615 | N623;
  assign N615 = N607 | N614;
  assign N607 = N599 | N606;
  assign N599 = N591 | N598;
  assign N591 = N583 | N590;
  assign N583 = N582 & din[1];
  assign N582 = N581 & N313;
  assign N581 = N580 & N311;
  assign N580 = N579 & N309;
  assign N579 = N578 & N307;
  assign N578 = N577 & N305;
  assign N577 = N6 & din[11];
  assign N590 = N589 & din[1];
  assign N589 = N588 & N313;
  assign N588 = N587 & N311;
  assign N587 = N586 & N309;
  assign N586 = N585 & N307;
  assign N585 = N584 & N305;
  assign N584 = N6 & din[10];
  assign N598 = N597 & din[1];
  assign N597 = N596 & N313;
  assign N596 = N595 & N311;
  assign N595 = N594 & N309;
  assign N594 = N593 & N307;
  assign N593 = N592 & N305;
  assign N592 = N6 & din[9];
  assign N606 = N605 & din[1];
  assign N605 = N604 & N313;
  assign N604 = N603 & N311;
  assign N603 = N602 & N309;
  assign N602 = N601 & N307;
  assign N601 = N600 & N305;
  assign N600 = N6 & din[8];
  assign N614 = N613 & din[1];
  assign N613 = N612 & N313;
  assign N612 = N611 & N311;
  assign N611 = N610 & N309;
  assign N610 = N609 & N307;
  assign N609 = N608 & N305;
  assign N608 = N6 & din[7];
  assign N623 = N622 & N362;
  assign N622 = N621 & N313;
  assign N621 = N620 & N311;
  assign N620 = N619 & N309;
  assign N619 = N618 & N307;
  assign N618 = N617 & N305;
  assign N617 = N616 & N303;
  assign N616 = din[15] & N352;
  assign N625 = N7 & N273;
  assign N627 = N7 & din[7];
  assign N629 = N7 & din[9];
  assign N631 = N7 & din[10];
  assign N633 = N7 & din[11];
  assign N635 = N352 & din[13];
  assign N8 = N285 & N303;
  assign N9 = N288 & N285;
  assign N10 = din[14] & N285;
  assign legal = N746 | N747;
  assign N746 = N743 | N745;
  assign N743 = N739 | N742;
  assign N739 = N734 | N738;
  assign N734 = N730 | N733;
  assign N730 = N728 | N729;
  assign N728 = N724 | N727;
  assign N724 = N720 | N723;
  assign N720 = N717 | N719;
  assign N717 = N713 | N716;
  assign N713 = N709 | N712;
  assign N709 = N705 | N708;
  assign N705 = N702 | N704;
  assign N702 = N698 | N701;
  assign N698 = N694 | N697;
  assign N694 = N691 | N693;
  assign N691 = N686 | N690;
  assign N686 = N682 | N685;
  assign N682 = N679 | N681;
  assign N679 = N675 | N678;
  assign N675 = N671 | N674;
  assign N671 = N668 | N670;
  assign N668 = N664 | N667;
  assign N664 = N660 | N663;
  assign N660 = N656 | N659;
  assign N656 = N653 | N655;
  assign N653 = N649 | N652;
  assign N649 = N645 | N648;
  assign N645 = N642 | N644;
  assign N642 = N638 | N641;
  assign N638 = N637 & N362;
  assign N637 = N636 & din[1];
  assign N636 = N8 & din[11];
  assign N641 = N640 & N362;
  assign N640 = N639 & din[1];
  assign N639 = N8 & din[6];
  assign N644 = N643 & N360;
  assign N643 = N9 & din[11];
  assign N648 = N647 & N362;
  assign N647 = N646 & din[1];
  assign N646 = N8 & din[5];
  assign N652 = N651 & N362;
  assign N651 = N650 & din[1];
  assign N650 = N8 & din[10];
  assign N655 = N654 & N360;
  assign N654 = N9 & din[6];
  assign N659 = N658 & din[0];
  assign N658 = N657 & N360;
  assign N657 = din[15] & N303;
  assign N663 = N662 & N362;
  assign N662 = N661 & din[1];
  assign N661 = N8 & din[9];
  assign N667 = N666 & din[0];
  assign N666 = N665 & N360;
  assign N665 = N303 & din[6];
  assign N670 = N669 & N360;
  assign N669 = N9 & din[5];
  assign N674 = N673 & N362;
  assign N673 = N672 & din[1];
  assign N672 = N8 & din[8];
  assign N678 = N677 & din[0];
  assign N677 = N676 & N360;
  assign N676 = N303 & din[5];
  assign N681 = N680 & N360;
  assign N680 = N9 & din[10];
  assign N685 = N684 & N362;
  assign N684 = N683 & din[1];
  assign N683 = N8 & din[7];
  assign N690 = N689 & din[0];
  assign N689 = N688 & N360;
  assign N688 = N687 & N380;
  assign N687 = din[12] & din[11];
  assign N693 = N692 & N360;
  assign N692 = N9 & din[9];
  assign N697 = N696 & N362;
  assign N696 = N695 & din[1];
  assign N695 = N8 & din[4];
  assign N701 = N700 & din[0];
  assign N700 = N699 & N360;
  assign N699 = din[13] & din[12];
  assign N704 = N703 & N360;
  assign N703 = N9 & din[8];
  assign N708 = N707 & N362;
  assign N707 = N706 & din[1];
  assign N706 = N8 & din[3];
  assign N712 = N711 & din[0];
  assign N711 = N710 & N360;
  assign N710 = din[13] & din[4];
  assign N716 = N715 & N362;
  assign N715 = N714 & din[1];
  assign N714 = N8 & din[2];
  assign N719 = N718 & N360;
  assign N718 = N9 & din[7];
  assign N723 = N722 & din[0];
  assign N722 = N721 & N360;
  assign N721 = din[13] & din[3];
  assign N727 = N726 & din[0];
  assign N726 = N725 & N360;
  assign N725 = din[13] & din[2];
  assign N729 = N10 & N360;
  assign N733 = N732 & din[0];
  assign N732 = N731 & N360;
  assign N731 = N352 & N303;
  assign N738 = N737 & N362;
  assign N737 = N736 & din[1];
  assign N736 = N735 & din[12];
  assign N735 = din[15] & N285;
  assign N742 = N741 & N362;
  assign N741 = N740 & din[1];
  assign N740 = N9 & N303;
  assign N745 = N744 & N360;
  assign N744 = N9 & din[12];
  assign N747 = N10 & N362;

endmodule