module ALU
(
  io_dw,
  io_fn,
  io_in2,
  io_in1,
  io_out,
  io_adder_out,
  io_cmp_out
);

  input [3:0] io_fn;
  input [63:0] io_in2;
  input [63:0] io_in1;
  output [63:0] io_out;
  output [63:0] io_adder_out;
  input io_dw;
  output io_cmp_out;
  wire [63:0] io_out,io_adder_out,in1_xor_in2,in2_inv,T12,T19,shift_logic,T121,shout,T117,T21,
  shout_l,T53,lg,T127,T122,T123;
  wire io_cmp_out,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,T1,T14,N23,T2,T8,N24,T3,T140_32,out_63_,out_62_,out_61_,out_60_,
  out_59_,out_58_,out_57_,out_56_,out_55_,out_54_,out_53_,out_52_,out_51_,out_50_,
  out_49_,out_48_,out_47_,out_46_,out_45_,out_44_,out_43_,out_42_,out_41_,out_40_,
  out_39_,out_38_,out_37_,out_36_,out_35_,out_34_,out_33_,out_32_,T137,N25,T22_61,
  T22_59,T22_57,T22_55,T22_53,T22_51,T22_49,T22_47,T22_45,T22_43,T22_41,T22_39,
  T22_37,T22_35,T22_33,T22_31,T22_29,T22_27,T22_25,T22_23,T22_21,T22_19,T22_17,T22_15,
  T22_13,T22_11,T22_9,T22_7,T22_5,T22_3,T22_1,T23_60,T23_58,T23_56,T23_54,T23_52,
  T23_50,T23_48,T23_46,T23_44,T23_42,T23_40,T23_38,T23_36,T23_34,T23_32,T23_30,
  T23_28,T23_26,T23_24,T23_22,T23_20,T23_18,T23_16,T23_14,T23_12,T23_10,T23_8,T23_6,
  T23_4,T23_2,T26_59,T26_58,T26_55,T26_54,T26_51,T26_50,T26_47,T26_46,T26_43,T26_42,
  T26_39,T26_38,T26_35,T26_34,T26_31,T26_30,T26_27,T26_26,T26_23,T26_22,T26_19,
  T26_18,T26_15,T26_14,T26_11,T26_10,T26_7,T26_6,T26_3,T26_2,T27_57,T27_56,T27_53,
  T27_52,T27_49,T27_48,T27_45,T27_44,T27_41,T27_40,T27_37,T27_36,T27_33,T27_32,T27_29,
  T27_28,T27_25,T27_24,T27_21,T27_20,T27_17,T27_16,T27_13,T27_12,T27_9,T27_8,T27_5,
  T27_4,T30_55,T30_54,T30_53,T30_52,T30_47,T30_46,T30_45,T30_44,T30_39,T30_38,
  T30_37,T30_36,T30_31,T30_30,T30_29,T30_28,T30_23,T30_22,T30_21,T30_20,T30_15,T30_14,
  T30_13,T30_12,T30_7,T30_6,T30_5,T30_4,T31_51,T31_50,T31_49,T31_48,T31_43,T31_42,
  T31_41,T31_40,T31_35,T31_34,T31_33,T31_32,T31_27,T31_26,T31_25,T31_24,T31_19,
  T31_18,T31_17,T31_16,T31_11,T31_10,T31_9,T31_8,T34_47,T34_46,T34_45,T34_44,T34_43,
  T34_42,T34_41,T34_40,T34_31,T34_30,T34_29,T34_28,T34_27,T34_26,T34_25,T34_24,
  T34_15,T34_14,T34_13,T34_12,T34_11,T34_10,T34_9,T34_8,T35_39,T35_38,T35_37,T35_36,
  T35_35,T35_34,T35_33,T35_32,T35_23,T35_22,T35_21,T35_20,T35_19,T35_18,T35_17,
  T35_16,T38_31,T38_30,T38_29,T38_28,T38_27,T38_26,T38_25,T38_24,T38_23,T38_22,T38_21,
  T38_20,T38_19,T38_18,T38_17,T38_16,T98,N26,T54_61,T54_59,T54_57,T54_55,T54_53,
  T54_51,T54_49,T54_47,T54_45,T54_43,T54_41,T54_39,T54_37,T54_35,T54_33,T54_31,
  T54_29,T54_27,T54_25,T54_23,T54_21,T54_19,T54_17,T54_15,T54_13,T54_11,T54_9,T54_7,
  T54_5,T54_3,T54_1,T55_60,T55_58,T55_56,T55_54,T55_52,T55_50,T55_48,T55_46,T55_44,
  T55_42,T55_40,T55_38,T55_36,T55_34,T55_32,T55_30,T55_28,T55_26,T55_24,T55_22,
  T55_20,T55_18,T55_16,T55_14,T55_12,T55_10,T55_8,T55_6,T55_4,T55_2,T58_59,T58_58,
  T58_55,T58_54,T58_51,T58_50,T58_47,T58_46,T58_43,T58_42,T58_39,T58_38,T58_35,T58_34,
  T58_31,T58_30,T58_27,T58_26,T58_23,T58_22,T58_19,T58_18,T58_15,T58_14,T58_11,
  T58_10,T58_7,T58_6,T58_3,T58_2,T59_57,T59_56,T59_53,T59_52,T59_49,T59_48,T59_45,
  T59_44,T59_41,T59_40,T59_37,T59_36,T59_33,T59_32,T59_29,T59_28,T59_25,T59_24,T59_21,
  T59_20,T59_17,T59_16,T59_13,T59_12,T59_9,T59_8,T59_5,T59_4,T62_55,T62_54,T62_53,
  T62_52,T62_47,T62_46,T62_45,T62_44,T62_39,T62_38,T62_37,T62_36,T62_31,T62_30,
  T62_29,T62_28,T62_23,T62_22,T62_21,T62_20,T62_15,T62_14,T62_13,T62_12,T62_7,T62_6,
  T62_5,T62_4,T63_51,T63_50,T63_49,T63_48,T63_43,T63_42,T63_41,T63_40,T63_35,T63_34,
  T63_33,T63_32,T63_27,T63_26,T63_25,T63_24,T63_19,T63_18,T63_17,T63_16,T63_11,
  T63_10,T63_9,T63_8,T66_47,T66_46,T66_45,T66_44,T66_43,T66_42,T66_41,T66_40,T66_31,
  T66_30,T66_29,T66_28,T66_27,T66_26,T66_25,T66_24,T66_15,T66_14,T66_13,T66_12,
  T66_11,T66_10,T66_9,T66_8,T67_39,T67_38,T67_37,T67_36,T67_35,T67_34,T67_33,T67_32,
  T67_23,T67_22,T67_21,T67_20,T67_19,T67_18,T67_17,T67_16,T70_31,T70_30,T70_29,
  T70_28,T70_27,T70_26,T70_25,T70_24,T70_23,T70_22,T70_21,T70_20,T70_19,T70_18,T70_17,
  T70_16,T91_0,T118,N27,T124,N28,T128,N29,T132,T134,T133,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  SV2V_UNCONNECTED_1;
  wire [63:63] T140,T22,T25,T54,T57;
  wire [62:62] T23,T55;
  wire [63:62] T26,T29,T58,T61;
  wire [61:60] T27,T59;
  wire [63:60] T30,T33,T62,T65;
  wire [59:56] T31,T63;
  wire [63:56] T34,T37,T66,T69;
  wire [55:48] T35,T67;
  wire [63:48] T38,T41,T70,T73;
  wire [47:32] T39,T71;
  wire [63:32] T42,shout_r;
  wire [5:5] shamt;
  wire [64:0] T51;
  wire [31:0] T77;
  wire [31:31] T91;
  wire [0:0] T153,T160;
  assign N0 = io_in1[63] ^ io_in2[63];
  assign T8 = ~N0;
  assign { SV2V_UNCONNECTED_1, shout_r, T42 } = $signed(T51) >>> { shamt[5:5], io_in2[4:0] };
  assign T133 = { 1'b1, 1'b1, 1'b0, 1'b0 } <= io_fn;
  assign N30 = ~io_dw;
  assign N31 = io_fn[2] | io_fn[3];
  assign N32 = io_fn[1] | N31;
  assign N33 = io_fn[0] | N32;
  assign N34 = ~N33;
  assign N35 = ~io_fn[3];
  assign N36 = ~io_fn[1];
  assign N37 = io_fn[2] | N35;
  assign N38 = N36 | N37;
  assign N39 = io_fn[0] | N38;
  assign N40 = ~N39;
  assign N41 = N36 | N31;
  assign N42 = io_fn[0] | N41;
  assign N43 = ~N42;
  assign N44 = ~io_fn[0];
  assign N45 = N44 | N41;
  assign N46 = ~N45;
  assign N47 = in1_xor_in2[62] | in1_xor_in2[63];
  assign N48 = in1_xor_in2[61] | N47;
  assign N49 = in1_xor_in2[60] | N48;
  assign N50 = in1_xor_in2[59] | N49;
  assign N51 = in1_xor_in2[58] | N50;
  assign N52 = in1_xor_in2[57] | N51;
  assign N53 = in1_xor_in2[56] | N52;
  assign N54 = in1_xor_in2[55] | N53;
  assign N55 = in1_xor_in2[54] | N54;
  assign N56 = in1_xor_in2[53] | N55;
  assign N57 = in1_xor_in2[52] | N56;
  assign N58 = in1_xor_in2[51] | N57;
  assign N59 = in1_xor_in2[50] | N58;
  assign N60 = in1_xor_in2[49] | N59;
  assign N61 = in1_xor_in2[48] | N60;
  assign N62 = in1_xor_in2[47] | N61;
  assign N63 = in1_xor_in2[46] | N62;
  assign N64 = in1_xor_in2[45] | N63;
  assign N65 = in1_xor_in2[44] | N64;
  assign N66 = in1_xor_in2[43] | N65;
  assign N67 = in1_xor_in2[42] | N66;
  assign N68 = in1_xor_in2[41] | N67;
  assign N69 = in1_xor_in2[40] | N68;
  assign N70 = in1_xor_in2[39] | N69;
  assign N71 = in1_xor_in2[38] | N70;
  assign N72 = in1_xor_in2[37] | N71;
  assign N73 = in1_xor_in2[36] | N72;
  assign N74 = in1_xor_in2[35] | N73;
  assign N75 = in1_xor_in2[34] | N74;
  assign N76 = in1_xor_in2[33] | N75;
  assign N77 = in1_xor_in2[32] | N76;
  assign N78 = in1_xor_in2[31] | N77;
  assign N79 = in1_xor_in2[30] | N78;
  assign N80 = in1_xor_in2[29] | N79;
  assign N81 = in1_xor_in2[28] | N80;
  assign N82 = in1_xor_in2[27] | N81;
  assign N83 = in1_xor_in2[26] | N82;
  assign N84 = in1_xor_in2[25] | N83;
  assign N85 = in1_xor_in2[24] | N84;
  assign N86 = in1_xor_in2[23] | N85;
  assign N87 = in1_xor_in2[22] | N86;
  assign N88 = in1_xor_in2[21] | N87;
  assign N89 = in1_xor_in2[20] | N88;
  assign N90 = in1_xor_in2[19] | N89;
  assign N91 = in1_xor_in2[18] | N90;
  assign N92 = in1_xor_in2[17] | N91;
  assign N93 = in1_xor_in2[16] | N92;
  assign N94 = in1_xor_in2[15] | N93;
  assign N95 = in1_xor_in2[14] | N94;
  assign N96 = in1_xor_in2[13] | N95;
  assign N97 = in1_xor_in2[12] | N96;
  assign N98 = in1_xor_in2[11] | N97;
  assign N99 = in1_xor_in2[10] | N98;
  assign N100 = in1_xor_in2[9] | N99;
  assign N101 = in1_xor_in2[8] | N100;
  assign N102 = in1_xor_in2[7] | N101;
  assign N103 = in1_xor_in2[6] | N102;
  assign N104 = in1_xor_in2[5] | N103;
  assign N105 = in1_xor_in2[4] | N104;
  assign N106 = in1_xor_in2[3] | N105;
  assign N107 = in1_xor_in2[2] | N106;
  assign N108 = in1_xor_in2[1] | N107;
  assign N109 = in1_xor_in2[0] | N108;
  assign N110 = ~N109;
  assign N111 = N44 | N32;
  assign N112 = ~N111;
  assign N113 = ~io_fn[2];
  assign N114 = N113 | io_fn[3];
  assign N115 = io_fn[1] | N114;
  assign N116 = N44 | N115;
  assign N117 = ~N116;
  assign N118 = N44 | N38;
  assign N119 = ~N118;
  assign N120 = io_fn[0] | N115;
  assign N121 = ~N120;
  assign N122 = N36 | N114;
  assign N123 = io_fn[0] | N122;
  assign N124 = ~N123;
  assign N125 = N44 | N122;
  assign N126 = ~N125;
  assign { T91[31:31], T91_0 } = 1'b0 - T153[0];
  assign T19 = io_in1 + in2_inv;
  assign io_adder_out = T19 + io_fn[3];
  assign { T140[63:63], T140_32 } = 1'b0 - io_out[31];
  assign T1 = (N1)? N110 : 
              (N2)? T2 : 1'b0;
  assign N1 = T14;
  assign N2 = N23;
  assign T2 = (N3)? io_adder_out[63] : 
              (N4)? T3 : 1'b0;
  assign N3 = T8;
  assign N4 = N24;
  assign T3 = (N5)? io_in2[63] : 
              (N6)? io_in1[63] : 1'b0;
  assign N5 = io_fn[1];
  assign N6 = N36;
  assign in2_inv = (N7)? T12 : 
                   (N8)? io_in2 : 1'b0;
  assign N7 = io_fn[3];
  assign N8 = N35;
  assign io_out[63:32] = (N9)? { T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140[63:63], T140_32 } : 
                         (N10)? { out_63_, out_62_, out_61_, out_60_, out_59_, out_58_, out_57_, out_56_, out_55_, out_54_, out_53_, out_52_, out_51_, out_50_, out_49_, out_48_, out_47_, out_46_, out_45_, out_44_, out_43_, out_42_, out_41_, out_40_, out_39_, out_38_, out_37_, out_36_, out_35_, out_34_, out_33_, out_32_ } : 1'b0;
  assign N9 = N30;
  assign N10 = io_dw;
  assign { out_63_, out_62_, out_61_, out_60_, out_59_, out_58_, out_57_, out_56_, out_55_, out_54_, out_53_, out_52_, out_51_, out_50_, out_49_, out_48_, out_47_, out_46_, out_45_, out_44_, out_43_, out_42_, out_41_, out_40_, out_39_, out_38_, out_37_, out_36_, out_35_, out_34_, out_33_, out_32_, io_out[31:0] } = (N11)? io_adder_out : 
                                                                                                                                                                                                                                                                                                                            (N12)? shift_logic : 1'b0;
  assign N11 = T137;
  assign N12 = N25;
  assign T21 = (N13)? shout_l : 
               (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N112;
  assign N14 = N111;
  assign T51[63:0] = (N15)? { T77, io_in1[31:0] } : 
                     (N16)? T53 : 1'b0;
  assign N15 = T98;
  assign N16 = N26;
  assign T77 = (N10)? io_in1[63:32] : 
               (N9)? { T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91[31:31], T91_0 } : 1'b0;
  assign T117 = (N17)? { shout_r, T42 } : 
                (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = T118;
  assign N18 = N27;
  assign T122 = (N19)? T123 : 
                (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = T124;
  assign N20 = N28;
  assign T127 = (N21)? in1_xor_in2 : 
                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = T128;
  assign N22 = N29;
  assign io_cmp_out = io_fn[0] ^ T1;
  assign N23 = ~T14;
  assign N24 = ~T8;
  assign in1_xor_in2[63] = io_in1[63] ^ in2_inv[63];
  assign in1_xor_in2[62] = io_in1[62] ^ in2_inv[62];
  assign in1_xor_in2[61] = io_in1[61] ^ in2_inv[61];
  assign in1_xor_in2[60] = io_in1[60] ^ in2_inv[60];
  assign in1_xor_in2[59] = io_in1[59] ^ in2_inv[59];
  assign in1_xor_in2[58] = io_in1[58] ^ in2_inv[58];
  assign in1_xor_in2[57] = io_in1[57] ^ in2_inv[57];
  assign in1_xor_in2[56] = io_in1[56] ^ in2_inv[56];
  assign in1_xor_in2[55] = io_in1[55] ^ in2_inv[55];
  assign in1_xor_in2[54] = io_in1[54] ^ in2_inv[54];
  assign in1_xor_in2[53] = io_in1[53] ^ in2_inv[53];
  assign in1_xor_in2[52] = io_in1[52] ^ in2_inv[52];
  assign in1_xor_in2[51] = io_in1[51] ^ in2_inv[51];
  assign in1_xor_in2[50] = io_in1[50] ^ in2_inv[50];
  assign in1_xor_in2[49] = io_in1[49] ^ in2_inv[49];
  assign in1_xor_in2[48] = io_in1[48] ^ in2_inv[48];
  assign in1_xor_in2[47] = io_in1[47] ^ in2_inv[47];
  assign in1_xor_in2[46] = io_in1[46] ^ in2_inv[46];
  assign in1_xor_in2[45] = io_in1[45] ^ in2_inv[45];
  assign in1_xor_in2[44] = io_in1[44] ^ in2_inv[44];
  assign in1_xor_in2[43] = io_in1[43] ^ in2_inv[43];
  assign in1_xor_in2[42] = io_in1[42] ^ in2_inv[42];
  assign in1_xor_in2[41] = io_in1[41] ^ in2_inv[41];
  assign in1_xor_in2[40] = io_in1[40] ^ in2_inv[40];
  assign in1_xor_in2[39] = io_in1[39] ^ in2_inv[39];
  assign in1_xor_in2[38] = io_in1[38] ^ in2_inv[38];
  assign in1_xor_in2[37] = io_in1[37] ^ in2_inv[37];
  assign in1_xor_in2[36] = io_in1[36] ^ in2_inv[36];
  assign in1_xor_in2[35] = io_in1[35] ^ in2_inv[35];
  assign in1_xor_in2[34] = io_in1[34] ^ in2_inv[34];
  assign in1_xor_in2[33] = io_in1[33] ^ in2_inv[33];
  assign in1_xor_in2[32] = io_in1[32] ^ in2_inv[32];
  assign in1_xor_in2[31] = io_in1[31] ^ in2_inv[31];
  assign in1_xor_in2[30] = io_in1[30] ^ in2_inv[30];
  assign in1_xor_in2[29] = io_in1[29] ^ in2_inv[29];
  assign in1_xor_in2[28] = io_in1[28] ^ in2_inv[28];
  assign in1_xor_in2[27] = io_in1[27] ^ in2_inv[27];
  assign in1_xor_in2[26] = io_in1[26] ^ in2_inv[26];
  assign in1_xor_in2[25] = io_in1[25] ^ in2_inv[25];
  assign in1_xor_in2[24] = io_in1[24] ^ in2_inv[24];
  assign in1_xor_in2[23] = io_in1[23] ^ in2_inv[23];
  assign in1_xor_in2[22] = io_in1[22] ^ in2_inv[22];
  assign in1_xor_in2[21] = io_in1[21] ^ in2_inv[21];
  assign in1_xor_in2[20] = io_in1[20] ^ in2_inv[20];
  assign in1_xor_in2[19] = io_in1[19] ^ in2_inv[19];
  assign in1_xor_in2[18] = io_in1[18] ^ in2_inv[18];
  assign in1_xor_in2[17] = io_in1[17] ^ in2_inv[17];
  assign in1_xor_in2[16] = io_in1[16] ^ in2_inv[16];
  assign in1_xor_in2[15] = io_in1[15] ^ in2_inv[15];
  assign in1_xor_in2[14] = io_in1[14] ^ in2_inv[14];
  assign in1_xor_in2[13] = io_in1[13] ^ in2_inv[13];
  assign in1_xor_in2[12] = io_in1[12] ^ in2_inv[12];
  assign in1_xor_in2[11] = io_in1[11] ^ in2_inv[11];
  assign in1_xor_in2[10] = io_in1[10] ^ in2_inv[10];
  assign in1_xor_in2[9] = io_in1[9] ^ in2_inv[9];
  assign in1_xor_in2[8] = io_in1[8] ^ in2_inv[8];
  assign in1_xor_in2[7] = io_in1[7] ^ in2_inv[7];
  assign in1_xor_in2[6] = io_in1[6] ^ in2_inv[6];
  assign in1_xor_in2[5] = io_in1[5] ^ in2_inv[5];
  assign in1_xor_in2[4] = io_in1[4] ^ in2_inv[4];
  assign in1_xor_in2[3] = io_in1[3] ^ in2_inv[3];
  assign in1_xor_in2[2] = io_in1[2] ^ in2_inv[2];
  assign in1_xor_in2[1] = io_in1[1] ^ in2_inv[1];
  assign in1_xor_in2[0] = io_in1[0] ^ in2_inv[0];
  assign T12[63] = ~io_in2[63];
  assign T12[62] = ~io_in2[62];
  assign T12[61] = ~io_in2[61];
  assign T12[60] = ~io_in2[60];
  assign T12[59] = ~io_in2[59];
  assign T12[58] = ~io_in2[58];
  assign T12[57] = ~io_in2[57];
  assign T12[56] = ~io_in2[56];
  assign T12[55] = ~io_in2[55];
  assign T12[54] = ~io_in2[54];
  assign T12[53] = ~io_in2[53];
  assign T12[52] = ~io_in2[52];
  assign T12[51] = ~io_in2[51];
  assign T12[50] = ~io_in2[50];
  assign T12[49] = ~io_in2[49];
  assign T12[48] = ~io_in2[48];
  assign T12[47] = ~io_in2[47];
  assign T12[46] = ~io_in2[46];
  assign T12[45] = ~io_in2[45];
  assign T12[44] = ~io_in2[44];
  assign T12[43] = ~io_in2[43];
  assign T12[42] = ~io_in2[42];
  assign T12[41] = ~io_in2[41];
  assign T12[40] = ~io_in2[40];
  assign T12[39] = ~io_in2[39];
  assign T12[38] = ~io_in2[38];
  assign T12[37] = ~io_in2[37];
  assign T12[36] = ~io_in2[36];
  assign T12[35] = ~io_in2[35];
  assign T12[34] = ~io_in2[34];
  assign T12[33] = ~io_in2[33];
  assign T12[32] = ~io_in2[32];
  assign T12[31] = ~io_in2[31];
  assign T12[30] = ~io_in2[30];
  assign T12[29] = ~io_in2[29];
  assign T12[28] = ~io_in2[28];
  assign T12[27] = ~io_in2[27];
  assign T12[26] = ~io_in2[26];
  assign T12[25] = ~io_in2[25];
  assign T12[24] = ~io_in2[24];
  assign T12[23] = ~io_in2[23];
  assign T12[22] = ~io_in2[22];
  assign T12[21] = ~io_in2[21];
  assign T12[20] = ~io_in2[20];
  assign T12[19] = ~io_in2[19];
  assign T12[18] = ~io_in2[18];
  assign T12[17] = ~io_in2[17];
  assign T12[16] = ~io_in2[16];
  assign T12[15] = ~io_in2[15];
  assign T12[14] = ~io_in2[14];
  assign T12[13] = ~io_in2[13];
  assign T12[12] = ~io_in2[12];
  assign T12[11] = ~io_in2[11];
  assign T12[10] = ~io_in2[10];
  assign T12[9] = ~io_in2[9];
  assign T12[8] = ~io_in2[8];
  assign T12[7] = ~io_in2[7];
  assign T12[6] = ~io_in2[6];
  assign T12[5] = ~io_in2[5];
  assign T12[4] = ~io_in2[4];
  assign T12[3] = ~io_in2[3];
  assign T12[2] = ~io_in2[2];
  assign T12[1] = ~io_in2[1];
  assign T12[0] = ~io_in2[0];
  assign T14 = ~io_fn[3];
  assign N25 = ~T137;
  assign shift_logic[63] = T121[63] | shout[63];
  assign shift_logic[62] = T121[62] | shout[62];
  assign shift_logic[61] = T121[61] | shout[61];
  assign shift_logic[60] = T121[60] | shout[60];
  assign shift_logic[59] = T121[59] | shout[59];
  assign shift_logic[58] = T121[58] | shout[58];
  assign shift_logic[57] = T121[57] | shout[57];
  assign shift_logic[56] = T121[56] | shout[56];
  assign shift_logic[55] = T121[55] | shout[55];
  assign shift_logic[54] = T121[54] | shout[54];
  assign shift_logic[53] = T121[53] | shout[53];
  assign shift_logic[52] = T121[52] | shout[52];
  assign shift_logic[51] = T121[51] | shout[51];
  assign shift_logic[50] = T121[50] | shout[50];
  assign shift_logic[49] = T121[49] | shout[49];
  assign shift_logic[48] = T121[48] | shout[48];
  assign shift_logic[47] = T121[47] | shout[47];
  assign shift_logic[46] = T121[46] | shout[46];
  assign shift_logic[45] = T121[45] | shout[45];
  assign shift_logic[44] = T121[44] | shout[44];
  assign shift_logic[43] = T121[43] | shout[43];
  assign shift_logic[42] = T121[42] | shout[42];
  assign shift_logic[41] = T121[41] | shout[41];
  assign shift_logic[40] = T121[40] | shout[40];
  assign shift_logic[39] = T121[39] | shout[39];
  assign shift_logic[38] = T121[38] | shout[38];
  assign shift_logic[37] = T121[37] | shout[37];
  assign shift_logic[36] = T121[36] | shout[36];
  assign shift_logic[35] = T121[35] | shout[35];
  assign shift_logic[34] = T121[34] | shout[34];
  assign shift_logic[33] = T121[33] | shout[33];
  assign shift_logic[32] = T121[32] | shout[32];
  assign shift_logic[31] = T121[31] | shout[31];
  assign shift_logic[30] = T121[30] | shout[30];
  assign shift_logic[29] = T121[29] | shout[29];
  assign shift_logic[28] = T121[28] | shout[28];
  assign shift_logic[27] = T121[27] | shout[27];
  assign shift_logic[26] = T121[26] | shout[26];
  assign shift_logic[25] = T121[25] | shout[25];
  assign shift_logic[24] = T121[24] | shout[24];
  assign shift_logic[23] = T121[23] | shout[23];
  assign shift_logic[22] = T121[22] | shout[22];
  assign shift_logic[21] = T121[21] | shout[21];
  assign shift_logic[20] = T121[20] | shout[20];
  assign shift_logic[19] = T121[19] | shout[19];
  assign shift_logic[18] = T121[18] | shout[18];
  assign shift_logic[17] = T121[17] | shout[17];
  assign shift_logic[16] = T121[16] | shout[16];
  assign shift_logic[15] = T121[15] | shout[15];
  assign shift_logic[14] = T121[14] | shout[14];
  assign shift_logic[13] = T121[13] | shout[13];
  assign shift_logic[12] = T121[12] | shout[12];
  assign shift_logic[11] = T121[11] | shout[11];
  assign shift_logic[10] = T121[10] | shout[10];
  assign shift_logic[9] = T121[9] | shout[9];
  assign shift_logic[8] = T121[8] | shout[8];
  assign shift_logic[7] = T121[7] | shout[7];
  assign shift_logic[6] = T121[6] | shout[6];
  assign shift_logic[5] = T121[5] | shout[5];
  assign shift_logic[4] = T121[4] | shout[4];
  assign shift_logic[3] = T121[3] | shout[3];
  assign shift_logic[2] = T121[2] | shout[2];
  assign shift_logic[1] = T121[1] | shout[1];
  assign shift_logic[0] = T121[0] | shout[0];
  assign shout[63] = T117[63] | T21[63];
  assign shout[62] = T117[62] | T21[62];
  assign shout[61] = T117[61] | T21[61];
  assign shout[60] = T117[60] | T21[60];
  assign shout[59] = T117[59] | T21[59];
  assign shout[58] = T117[58] | T21[58];
  assign shout[57] = T117[57] | T21[57];
  assign shout[56] = T117[56] | T21[56];
  assign shout[55] = T117[55] | T21[55];
  assign shout[54] = T117[54] | T21[54];
  assign shout[53] = T117[53] | T21[53];
  assign shout[52] = T117[52] | T21[52];
  assign shout[51] = T117[51] | T21[51];
  assign shout[50] = T117[50] | T21[50];
  assign shout[49] = T117[49] | T21[49];
  assign shout[48] = T117[48] | T21[48];
  assign shout[47] = T117[47] | T21[47];
  assign shout[46] = T117[46] | T21[46];
  assign shout[45] = T117[45] | T21[45];
  assign shout[44] = T117[44] | T21[44];
  assign shout[43] = T117[43] | T21[43];
  assign shout[42] = T117[42] | T21[42];
  assign shout[41] = T117[41] | T21[41];
  assign shout[40] = T117[40] | T21[40];
  assign shout[39] = T117[39] | T21[39];
  assign shout[38] = T117[38] | T21[38];
  assign shout[37] = T117[37] | T21[37];
  assign shout[36] = T117[36] | T21[36];
  assign shout[35] = T117[35] | T21[35];
  assign shout[34] = T117[34] | T21[34];
  assign shout[33] = T117[33] | T21[33];
  assign shout[32] = T117[32] | T21[32];
  assign shout[31] = T117[31] | T21[31];
  assign shout[30] = T117[30] | T21[30];
  assign shout[29] = T117[29] | T21[29];
  assign shout[28] = T117[28] | T21[28];
  assign shout[27] = T117[27] | T21[27];
  assign shout[26] = T117[26] | T21[26];
  assign shout[25] = T117[25] | T21[25];
  assign shout[24] = T117[24] | T21[24];
  assign shout[23] = T117[23] | T21[23];
  assign shout[22] = T117[22] | T21[22];
  assign shout[21] = T117[21] | T21[21];
  assign shout[20] = T117[20] | T21[20];
  assign shout[19] = T117[19] | T21[19];
  assign shout[18] = T117[18] | T21[18];
  assign shout[17] = T117[17] | T21[17];
  assign shout[16] = T117[16] | T21[16];
  assign shout[15] = T117[15] | T21[15];
  assign shout[14] = T117[14] | T21[14];
  assign shout[13] = T117[13] | T21[13];
  assign shout[12] = T117[12] | T21[12];
  assign shout[11] = T117[11] | T21[11];
  assign shout[10] = T117[10] | T21[10];
  assign shout[9] = T117[9] | T21[9];
  assign shout[8] = T117[8] | T21[8];
  assign shout[7] = T117[7] | T21[7];
  assign shout[6] = T117[6] | T21[6];
  assign shout[5] = T117[5] | T21[5];
  assign shout[4] = T117[4] | T21[4];
  assign shout[3] = T117[3] | T21[3];
  assign shout[2] = T117[2] | T21[2];
  assign shout[1] = T117[1] | T21[1];
  assign shout[0] = T117[0] | T21[0];
  assign shout_l[63] = 1'b0 | T22[63];
  assign shout_l[62] = T25[63] | 1'b0;
  assign shout_l[61] = 1'b0 | T22_61;
  assign shout_l[60] = T23[62] | 1'b0;
  assign shout_l[59] = 1'b0 | T22_59;
  assign shout_l[58] = T23_60 | 1'b0;
  assign shout_l[57] = 1'b0 | T22_57;
  assign shout_l[56] = T23_58 | 1'b0;
  assign shout_l[55] = 1'b0 | T22_55;
  assign shout_l[54] = T23_56 | 1'b0;
  assign shout_l[53] = 1'b0 | T22_53;
  assign shout_l[52] = T23_54 | 1'b0;
  assign shout_l[51] = 1'b0 | T22_51;
  assign shout_l[50] = T23_52 | 1'b0;
  assign shout_l[49] = 1'b0 | T22_49;
  assign shout_l[48] = T23_50 | 1'b0;
  assign shout_l[47] = 1'b0 | T22_47;
  assign shout_l[46] = T23_48 | 1'b0;
  assign shout_l[45] = 1'b0 | T22_45;
  assign shout_l[44] = T23_46 | 1'b0;
  assign shout_l[43] = 1'b0 | T22_43;
  assign shout_l[42] = T23_44 | 1'b0;
  assign shout_l[41] = 1'b0 | T22_41;
  assign shout_l[40] = T23_42 | 1'b0;
  assign shout_l[39] = 1'b0 | T22_39;
  assign shout_l[38] = T23_40 | 1'b0;
  assign shout_l[37] = 1'b0 | T22_37;
  assign shout_l[36] = T23_38 | 1'b0;
  assign shout_l[35] = 1'b0 | T22_35;
  assign shout_l[34] = T23_36 | 1'b0;
  assign shout_l[33] = 1'b0 | T22_33;
  assign shout_l[32] = T23_34 | 1'b0;
  assign shout_l[31] = 1'b0 | T22_31;
  assign shout_l[30] = T23_32 | 1'b0;
  assign shout_l[29] = 1'b0 | T22_29;
  assign shout_l[28] = T23_30 | 1'b0;
  assign shout_l[27] = 1'b0 | T22_27;
  assign shout_l[26] = T23_28 | 1'b0;
  assign shout_l[25] = 1'b0 | T22_25;
  assign shout_l[24] = T23_26 | 1'b0;
  assign shout_l[23] = 1'b0 | T22_23;
  assign shout_l[22] = T23_24 | 1'b0;
  assign shout_l[21] = 1'b0 | T22_21;
  assign shout_l[20] = T23_22 | 1'b0;
  assign shout_l[19] = 1'b0 | T22_19;
  assign shout_l[18] = T23_20 | 1'b0;
  assign shout_l[17] = 1'b0 | T22_17;
  assign shout_l[16] = T23_18 | 1'b0;
  assign shout_l[15] = 1'b0 | T22_15;
  assign shout_l[14] = T23_16 | 1'b0;
  assign shout_l[13] = 1'b0 | T22_13;
  assign shout_l[12] = T23_14 | 1'b0;
  assign shout_l[11] = 1'b0 | T22_11;
  assign shout_l[10] = T23_12 | 1'b0;
  assign shout_l[9] = 1'b0 | T22_9;
  assign shout_l[8] = T23_10 | 1'b0;
  assign shout_l[7] = 1'b0 | T22_7;
  assign shout_l[6] = T23_8 | 1'b0;
  assign shout_l[5] = 1'b0 | T22_5;
  assign shout_l[4] = T23_6 | 1'b0;
  assign shout_l[3] = 1'b0 | T22_3;
  assign shout_l[2] = T23_4 | 1'b0;
  assign shout_l[1] = 1'b0 | T22_1;
  assign shout_l[0] = T23_2 | 1'b0;
  assign T25[63] = 1'b0 | T26[63];
  assign T22[63] = 1'b0 | T26[62];
  assign T23[62] = T29[63] | 1'b0;
  assign T22_61 = T29[62] | 1'b0;
  assign T23_60 = 1'b0 | T26_59;
  assign T22_59 = 1'b0 | T26_58;
  assign T23_58 = T27[61] | 1'b0;
  assign T22_57 = T27[60] | 1'b0;
  assign T23_56 = 1'b0 | T26_55;
  assign T22_55 = 1'b0 | T26_54;
  assign T23_54 = T27_57 | 1'b0;
  assign T22_53 = T27_56 | 1'b0;
  assign T23_52 = 1'b0 | T26_51;
  assign T22_51 = 1'b0 | T26_50;
  assign T23_50 = T27_53 | 1'b0;
  assign T22_49 = T27_52 | 1'b0;
  assign T23_48 = 1'b0 | T26_47;
  assign T22_47 = 1'b0 | T26_46;
  assign T23_46 = T27_49 | 1'b0;
  assign T22_45 = T27_48 | 1'b0;
  assign T23_44 = 1'b0 | T26_43;
  assign T22_43 = 1'b0 | T26_42;
  assign T23_42 = T27_45 | 1'b0;
  assign T22_41 = T27_44 | 1'b0;
  assign T23_40 = 1'b0 | T26_39;
  assign T22_39 = 1'b0 | T26_38;
  assign T23_38 = T27_41 | 1'b0;
  assign T22_37 = T27_40 | 1'b0;
  assign T23_36 = 1'b0 | T26_35;
  assign T22_35 = 1'b0 | T26_34;
  assign T23_34 = T27_37 | 1'b0;
  assign T22_33 = T27_36 | 1'b0;
  assign T23_32 = 1'b0 | T26_31;
  assign T22_31 = 1'b0 | T26_30;
  assign T23_30 = T27_33 | 1'b0;
  assign T22_29 = T27_32 | 1'b0;
  assign T23_28 = 1'b0 | T26_27;
  assign T22_27 = 1'b0 | T26_26;
  assign T23_26 = T27_29 | 1'b0;
  assign T22_25 = T27_28 | 1'b0;
  assign T23_24 = 1'b0 | T26_23;
  assign T22_23 = 1'b0 | T26_22;
  assign T23_22 = T27_25 | 1'b0;
  assign T22_21 = T27_24 | 1'b0;
  assign T23_20 = 1'b0 | T26_19;
  assign T22_19 = 1'b0 | T26_18;
  assign T23_18 = T27_21 | 1'b0;
  assign T22_17 = T27_20 | 1'b0;
  assign T23_16 = 1'b0 | T26_15;
  assign T22_15 = 1'b0 | T26_14;
  assign T23_14 = T27_17 | 1'b0;
  assign T22_13 = T27_16 | 1'b0;
  assign T23_12 = 1'b0 | T26_11;
  assign T22_11 = 1'b0 | T26_10;
  assign T23_10 = T27_13 | 1'b0;
  assign T22_9 = T27_12 | 1'b0;
  assign T23_8 = 1'b0 | T26_7;
  assign T22_7 = 1'b0 | T26_6;
  assign T23_6 = T27_9 | 1'b0;
  assign T22_5 = T27_8 | 1'b0;
  assign T23_4 = 1'b0 | T26_3;
  assign T22_3 = 1'b0 | T26_2;
  assign T23_2 = T27_5 | 1'b0;
  assign T22_1 = T27_4 | 1'b0;
  assign T29[63] = 1'b0 | T30[63];
  assign T29[62] = 1'b0 | T30[62];
  assign T26[63] = 1'b0 | T30[61];
  assign T26[62] = 1'b0 | T30[60];
  assign T27[61] = T33[63] | 1'b0;
  assign T27[60] = T33[62] | 1'b0;
  assign T26_59 = T33[61] | 1'b0;
  assign T26_58 = T33[60] | 1'b0;
  assign T27_57 = 1'b0 | T30_55;
  assign T27_56 = 1'b0 | T30_54;
  assign T26_55 = 1'b0 | T30_53;
  assign T26_54 = 1'b0 | T30_52;
  assign T27_53 = T31[59] | 1'b0;
  assign T27_52 = T31[58] | 1'b0;
  assign T26_51 = T31[57] | 1'b0;
  assign T26_50 = T31[56] | 1'b0;
  assign T27_49 = 1'b0 | T30_47;
  assign T27_48 = 1'b0 | T30_46;
  assign T26_47 = 1'b0 | T30_45;
  assign T26_46 = 1'b0 | T30_44;
  assign T27_45 = T31_51 | 1'b0;
  assign T27_44 = T31_50 | 1'b0;
  assign T26_43 = T31_49 | 1'b0;
  assign T26_42 = T31_48 | 1'b0;
  assign T27_41 = 1'b0 | T30_39;
  assign T27_40 = 1'b0 | T30_38;
  assign T26_39 = 1'b0 | T30_37;
  assign T26_38 = 1'b0 | T30_36;
  assign T27_37 = T31_43 | 1'b0;
  assign T27_36 = T31_42 | 1'b0;
  assign T26_35 = T31_41 | 1'b0;
  assign T26_34 = T31_40 | 1'b0;
  assign T27_33 = 1'b0 | T30_31;
  assign T27_32 = 1'b0 | T30_30;
  assign T26_31 = 1'b0 | T30_29;
  assign T26_30 = 1'b0 | T30_28;
  assign T27_29 = T31_35 | 1'b0;
  assign T27_28 = T31_34 | 1'b0;
  assign T26_27 = T31_33 | 1'b0;
  assign T26_26 = T31_32 | 1'b0;
  assign T27_25 = 1'b0 | T30_23;
  assign T27_24 = 1'b0 | T30_22;
  assign T26_23 = 1'b0 | T30_21;
  assign T26_22 = 1'b0 | T30_20;
  assign T27_21 = T31_27 | 1'b0;
  assign T27_20 = T31_26 | 1'b0;
  assign T26_19 = T31_25 | 1'b0;
  assign T26_18 = T31_24 | 1'b0;
  assign T27_17 = 1'b0 | T30_15;
  assign T27_16 = 1'b0 | T30_14;
  assign T26_15 = 1'b0 | T30_13;
  assign T26_14 = 1'b0 | T30_12;
  assign T27_13 = T31_19 | 1'b0;
  assign T27_12 = T31_18 | 1'b0;
  assign T26_11 = T31_17 | 1'b0;
  assign T26_10 = T31_16 | 1'b0;
  assign T27_9 = 1'b0 | T30_7;
  assign T27_8 = 1'b0 | T30_6;
  assign T26_7 = 1'b0 | T30_5;
  assign T26_6 = 1'b0 | T30_4;
  assign T27_5 = T31_11 | 1'b0;
  assign T27_4 = T31_10 | 1'b0;
  assign T26_3 = T31_9 | 1'b0;
  assign T26_2 = T31_8 | 1'b0;
  assign T33[63] = 1'b0 | T34[63];
  assign T33[62] = 1'b0 | T34[62];
  assign T33[61] = 1'b0 | T34[61];
  assign T33[60] = 1'b0 | T34[60];
  assign T30[63] = 1'b0 | T34[59];
  assign T30[62] = 1'b0 | T34[58];
  assign T30[61] = 1'b0 | T34[57];
  assign T30[60] = 1'b0 | T34[56];
  assign T31[59] = T37[63] | 1'b0;
  assign T31[58] = T37[62] | 1'b0;
  assign T31[57] = T37[61] | 1'b0;
  assign T31[56] = T37[60] | 1'b0;
  assign T30_55 = T37[59] | 1'b0;
  assign T30_54 = T37[58] | 1'b0;
  assign T30_53 = T37[57] | 1'b0;
  assign T30_52 = T37[56] | 1'b0;
  assign T31_51 = 1'b0 | T34_47;
  assign T31_50 = 1'b0 | T34_46;
  assign T31_49 = 1'b0 | T34_45;
  assign T31_48 = 1'b0 | T34_44;
  assign T30_47 = 1'b0 | T34_43;
  assign T30_46 = 1'b0 | T34_42;
  assign T30_45 = 1'b0 | T34_41;
  assign T30_44 = 1'b0 | T34_40;
  assign T31_43 = T35[55] | 1'b0;
  assign T31_42 = T35[54] | 1'b0;
  assign T31_41 = T35[53] | 1'b0;
  assign T31_40 = T35[52] | 1'b0;
  assign T30_39 = T35[51] | 1'b0;
  assign T30_38 = T35[50] | 1'b0;
  assign T30_37 = T35[49] | 1'b0;
  assign T30_36 = T35[48] | 1'b0;
  assign T31_35 = 1'b0 | T34_31;
  assign T31_34 = 1'b0 | T34_30;
  assign T31_33 = 1'b0 | T34_29;
  assign T31_32 = 1'b0 | T34_28;
  assign T30_31 = 1'b0 | T34_27;
  assign T30_30 = 1'b0 | T34_26;
  assign T30_29 = 1'b0 | T34_25;
  assign T30_28 = 1'b0 | T34_24;
  assign T31_27 = T35_39 | 1'b0;
  assign T31_26 = T35_38 | 1'b0;
  assign T31_25 = T35_37 | 1'b0;
  assign T31_24 = T35_36 | 1'b0;
  assign T30_23 = T35_35 | 1'b0;
  assign T30_22 = T35_34 | 1'b0;
  assign T30_21 = T35_33 | 1'b0;
  assign T30_20 = T35_32 | 1'b0;
  assign T31_19 = 1'b0 | T34_15;
  assign T31_18 = 1'b0 | T34_14;
  assign T31_17 = 1'b0 | T34_13;
  assign T31_16 = 1'b0 | T34_12;
  assign T30_15 = 1'b0 | T34_11;
  assign T30_14 = 1'b0 | T34_10;
  assign T30_13 = 1'b0 | T34_9;
  assign T30_12 = 1'b0 | T34_8;
  assign T31_11 = T35_23 | 1'b0;
  assign T31_10 = T35_22 | 1'b0;
  assign T31_9 = T35_21 | 1'b0;
  assign T31_8 = T35_20 | 1'b0;
  assign T30_7 = T35_19 | 1'b0;
  assign T30_6 = T35_18 | 1'b0;
  assign T30_5 = T35_17 | 1'b0;
  assign T30_4 = T35_16 | 1'b0;
  assign T37[63] = 1'b0 | T38[63];
  assign T37[62] = 1'b0 | T38[62];
  assign T37[61] = 1'b0 | T38[61];
  assign T37[60] = 1'b0 | T38[60];
  assign T37[59] = 1'b0 | T38[59];
  assign T37[58] = 1'b0 | T38[58];
  assign T37[57] = 1'b0 | T38[57];
  assign T37[56] = 1'b0 | T38[56];
  assign T34[63] = 1'b0 | T38[55];
  assign T34[62] = 1'b0 | T38[54];
  assign T34[61] = 1'b0 | T38[53];
  assign T34[60] = 1'b0 | T38[52];
  assign T34[59] = 1'b0 | T38[51];
  assign T34[58] = 1'b0 | T38[50];
  assign T34[57] = 1'b0 | T38[49];
  assign T34[56] = 1'b0 | T38[48];
  assign T35[55] = T41[63] | 1'b0;
  assign T35[54] = T41[62] | 1'b0;
  assign T35[53] = T41[61] | 1'b0;
  assign T35[52] = T41[60] | 1'b0;
  assign T35[51] = T41[59] | 1'b0;
  assign T35[50] = T41[58] | 1'b0;
  assign T35[49] = T41[57] | 1'b0;
  assign T35[48] = T41[56] | 1'b0;
  assign T34_47 = T41[55] | 1'b0;
  assign T34_46 = T41[54] | 1'b0;
  assign T34_45 = T41[53] | 1'b0;
  assign T34_44 = T41[52] | 1'b0;
  assign T34_43 = T41[51] | 1'b0;
  assign T34_42 = T41[50] | 1'b0;
  assign T34_41 = T41[49] | 1'b0;
  assign T34_40 = T41[48] | 1'b0;
  assign T35_39 = 1'b0 | T38_31;
  assign T35_38 = 1'b0 | T38_30;
  assign T35_37 = 1'b0 | T38_29;
  assign T35_36 = 1'b0 | T38_28;
  assign T35_35 = 1'b0 | T38_27;
  assign T35_34 = 1'b0 | T38_26;
  assign T35_33 = 1'b0 | T38_25;
  assign T35_32 = 1'b0 | T38_24;
  assign T34_31 = 1'b0 | T38_23;
  assign T34_30 = 1'b0 | T38_22;
  assign T34_29 = 1'b0 | T38_21;
  assign T34_28 = 1'b0 | T38_20;
  assign T34_27 = 1'b0 | T38_19;
  assign T34_26 = 1'b0 | T38_18;
  assign T34_25 = 1'b0 | T38_17;
  assign T34_24 = 1'b0 | T38_16;
  assign T35_23 = T39[47] | 1'b0;
  assign T35_22 = T39[46] | 1'b0;
  assign T35_21 = T39[45] | 1'b0;
  assign T35_20 = T39[44] | 1'b0;
  assign T35_19 = T39[43] | 1'b0;
  assign T35_18 = T39[42] | 1'b0;
  assign T35_17 = T39[41] | 1'b0;
  assign T35_16 = T39[40] | 1'b0;
  assign T34_15 = T39[39] | 1'b0;
  assign T34_14 = T39[38] | 1'b0;
  assign T34_13 = T39[37] | 1'b0;
  assign T34_12 = T39[36] | 1'b0;
  assign T34_11 = T39[35] | 1'b0;
  assign T34_10 = T39[34] | 1'b0;
  assign T34_9 = T39[33] | 1'b0;
  assign T34_8 = T39[32] | 1'b0;
  assign T41[63] = 1'b0 | T42[63];
  assign T41[62] = 1'b0 | T42[62];
  assign T41[61] = 1'b0 | T42[61];
  assign T41[60] = 1'b0 | T42[60];
  assign T41[59] = 1'b0 | T42[59];
  assign T41[58] = 1'b0 | T42[58];
  assign T41[57] = 1'b0 | T42[57];
  assign T41[56] = 1'b0 | T42[56];
  assign T41[55] = 1'b0 | T42[55];
  assign T41[54] = 1'b0 | T42[54];
  assign T41[53] = 1'b0 | T42[53];
  assign T41[52] = 1'b0 | T42[52];
  assign T41[51] = 1'b0 | T42[51];
  assign T41[50] = 1'b0 | T42[50];
  assign T41[49] = 1'b0 | T42[49];
  assign T41[48] = 1'b0 | T42[48];
  assign T38[63] = 1'b0 | T42[47];
  assign T38[62] = 1'b0 | T42[46];
  assign T38[61] = 1'b0 | T42[45];
  assign T38[60] = 1'b0 | T42[44];
  assign T38[59] = 1'b0 | T42[43];
  assign T38[58] = 1'b0 | T42[42];
  assign T38[57] = 1'b0 | T42[41];
  assign T38[56] = 1'b0 | T42[40];
  assign T38[55] = 1'b0 | T42[39];
  assign T38[54] = 1'b0 | T42[38];
  assign T38[53] = 1'b0 | T42[37];
  assign T38[52] = 1'b0 | T42[36];
  assign T38[51] = 1'b0 | T42[35];
  assign T38[50] = 1'b0 | T42[34];
  assign T38[49] = 1'b0 | T42[33];
  assign T38[48] = 1'b0 | T42[32];
  assign T39[47] = shout_r[63] | 1'b0;
  assign T39[46] = shout_r[62] | 1'b0;
  assign T39[45] = shout_r[61] | 1'b0;
  assign T39[44] = shout_r[60] | 1'b0;
  assign T39[43] = shout_r[59] | 1'b0;
  assign T39[42] = shout_r[58] | 1'b0;
  assign T39[41] = shout_r[57] | 1'b0;
  assign T39[40] = shout_r[56] | 1'b0;
  assign T39[39] = shout_r[55] | 1'b0;
  assign T39[38] = shout_r[54] | 1'b0;
  assign T39[37] = shout_r[53] | 1'b0;
  assign T39[36] = shout_r[52] | 1'b0;
  assign T39[35] = shout_r[51] | 1'b0;
  assign T39[34] = shout_r[50] | 1'b0;
  assign T39[33] = shout_r[49] | 1'b0;
  assign T39[32] = shout_r[48] | 1'b0;
  assign T38_31 = shout_r[47] | 1'b0;
  assign T38_30 = shout_r[46] | 1'b0;
  assign T38_29 = shout_r[45] | 1'b0;
  assign T38_28 = shout_r[44] | 1'b0;
  assign T38_27 = shout_r[43] | 1'b0;
  assign T38_26 = shout_r[42] | 1'b0;
  assign T38_25 = shout_r[41] | 1'b0;
  assign T38_24 = shout_r[40] | 1'b0;
  assign T38_23 = shout_r[39] | 1'b0;
  assign T38_22 = shout_r[38] | 1'b0;
  assign T38_21 = shout_r[37] | 1'b0;
  assign T38_20 = shout_r[36] | 1'b0;
  assign T38_19 = shout_r[35] | 1'b0;
  assign T38_18 = shout_r[34] | 1'b0;
  assign T38_17 = shout_r[33] | 1'b0;
  assign T38_16 = shout_r[32] | 1'b0;
  assign shamt[5] = io_in2[5] & io_dw;
  assign N26 = ~T98;
  assign T53[63] = 1'b0 | T54[63];
  assign T53[62] = T57[63] | 1'b0;
  assign T53[61] = 1'b0 | T54_61;
  assign T53[60] = T55[62] | 1'b0;
  assign T53[59] = 1'b0 | T54_59;
  assign T53[58] = T55_60 | 1'b0;
  assign T53[57] = 1'b0 | T54_57;
  assign T53[56] = T55_58 | 1'b0;
  assign T53[55] = 1'b0 | T54_55;
  assign T53[54] = T55_56 | 1'b0;
  assign T53[53] = 1'b0 | T54_53;
  assign T53[52] = T55_54 | 1'b0;
  assign T53[51] = 1'b0 | T54_51;
  assign T53[50] = T55_52 | 1'b0;
  assign T53[49] = 1'b0 | T54_49;
  assign T53[48] = T55_50 | 1'b0;
  assign T53[47] = 1'b0 | T54_47;
  assign T53[46] = T55_48 | 1'b0;
  assign T53[45] = 1'b0 | T54_45;
  assign T53[44] = T55_46 | 1'b0;
  assign T53[43] = 1'b0 | T54_43;
  assign T53[42] = T55_44 | 1'b0;
  assign T53[41] = 1'b0 | T54_41;
  assign T53[40] = T55_42 | 1'b0;
  assign T53[39] = 1'b0 | T54_39;
  assign T53[38] = T55_40 | 1'b0;
  assign T53[37] = 1'b0 | T54_37;
  assign T53[36] = T55_38 | 1'b0;
  assign T53[35] = 1'b0 | T54_35;
  assign T53[34] = T55_36 | 1'b0;
  assign T53[33] = 1'b0 | T54_33;
  assign T53[32] = T55_34 | 1'b0;
  assign T53[31] = 1'b0 | T54_31;
  assign T53[30] = T55_32 | 1'b0;
  assign T53[29] = 1'b0 | T54_29;
  assign T53[28] = T55_30 | 1'b0;
  assign T53[27] = 1'b0 | T54_27;
  assign T53[26] = T55_28 | 1'b0;
  assign T53[25] = 1'b0 | T54_25;
  assign T53[24] = T55_26 | 1'b0;
  assign T53[23] = 1'b0 | T54_23;
  assign T53[22] = T55_24 | 1'b0;
  assign T53[21] = 1'b0 | T54_21;
  assign T53[20] = T55_22 | 1'b0;
  assign T53[19] = 1'b0 | T54_19;
  assign T53[18] = T55_20 | 1'b0;
  assign T53[17] = 1'b0 | T54_17;
  assign T53[16] = T55_18 | 1'b0;
  assign T53[15] = 1'b0 | T54_15;
  assign T53[14] = T55_16 | 1'b0;
  assign T53[13] = 1'b0 | T54_13;
  assign T53[12] = T55_14 | 1'b0;
  assign T53[11] = 1'b0 | T54_11;
  assign T53[10] = T55_12 | 1'b0;
  assign T53[9] = 1'b0 | T54_9;
  assign T53[8] = T55_10 | 1'b0;
  assign T53[7] = 1'b0 | T54_7;
  assign T53[6] = T55_8 | 1'b0;
  assign T53[5] = 1'b0 | T54_5;
  assign T53[4] = T55_6 | 1'b0;
  assign T53[3] = 1'b0 | T54_3;
  assign T53[2] = T55_4 | 1'b0;
  assign T53[1] = 1'b0 | T54_1;
  assign T53[0] = T55_2 | 1'b0;
  assign T57[63] = 1'b0 | T58[63];
  assign T54[63] = 1'b0 | T58[62];
  assign T55[62] = T61[63] | 1'b0;
  assign T54_61 = T61[62] | 1'b0;
  assign T55_60 = 1'b0 | T58_59;
  assign T54_59 = 1'b0 | T58_58;
  assign T55_58 = T59[61] | 1'b0;
  assign T54_57 = T59[60] | 1'b0;
  assign T55_56 = 1'b0 | T58_55;
  assign T54_55 = 1'b0 | T58_54;
  assign T55_54 = T59_57 | 1'b0;
  assign T54_53 = T59_56 | 1'b0;
  assign T55_52 = 1'b0 | T58_51;
  assign T54_51 = 1'b0 | T58_50;
  assign T55_50 = T59_53 | 1'b0;
  assign T54_49 = T59_52 | 1'b0;
  assign T55_48 = 1'b0 | T58_47;
  assign T54_47 = 1'b0 | T58_46;
  assign T55_46 = T59_49 | 1'b0;
  assign T54_45 = T59_48 | 1'b0;
  assign T55_44 = 1'b0 | T58_43;
  assign T54_43 = 1'b0 | T58_42;
  assign T55_42 = T59_45 | 1'b0;
  assign T54_41 = T59_44 | 1'b0;
  assign T55_40 = 1'b0 | T58_39;
  assign T54_39 = 1'b0 | T58_38;
  assign T55_38 = T59_41 | 1'b0;
  assign T54_37 = T59_40 | 1'b0;
  assign T55_36 = 1'b0 | T58_35;
  assign T54_35 = 1'b0 | T58_34;
  assign T55_34 = T59_37 | 1'b0;
  assign T54_33 = T59_36 | 1'b0;
  assign T55_32 = 1'b0 | T58_31;
  assign T54_31 = 1'b0 | T58_30;
  assign T55_30 = T59_33 | 1'b0;
  assign T54_29 = T59_32 | 1'b0;
  assign T55_28 = 1'b0 | T58_27;
  assign T54_27 = 1'b0 | T58_26;
  assign T55_26 = T59_29 | 1'b0;
  assign T54_25 = T59_28 | 1'b0;
  assign T55_24 = 1'b0 | T58_23;
  assign T54_23 = 1'b0 | T58_22;
  assign T55_22 = T59_25 | 1'b0;
  assign T54_21 = T59_24 | 1'b0;
  assign T55_20 = 1'b0 | T58_19;
  assign T54_19 = 1'b0 | T58_18;
  assign T55_18 = T59_21 | 1'b0;
  assign T54_17 = T59_20 | 1'b0;
  assign T55_16 = 1'b0 | T58_15;
  assign T54_15 = 1'b0 | T58_14;
  assign T55_14 = T59_17 | 1'b0;
  assign T54_13 = T59_16 | 1'b0;
  assign T55_12 = 1'b0 | T58_11;
  assign T54_11 = 1'b0 | T58_10;
  assign T55_10 = T59_13 | 1'b0;
  assign T54_9 = T59_12 | 1'b0;
  assign T55_8 = 1'b0 | T58_7;
  assign T54_7 = 1'b0 | T58_6;
  assign T55_6 = T59_9 | 1'b0;
  assign T54_5 = T59_8 | 1'b0;
  assign T55_4 = 1'b0 | T58_3;
  assign T54_3 = 1'b0 | T58_2;
  assign T55_2 = T59_5 | 1'b0;
  assign T54_1 = T59_4 | 1'b0;
  assign T61[63] = 1'b0 | T62[63];
  assign T61[62] = 1'b0 | T62[62];
  assign T58[63] = 1'b0 | T62[61];
  assign T58[62] = 1'b0 | T62[60];
  assign T59[61] = T65[63] | 1'b0;
  assign T59[60] = T65[62] | 1'b0;
  assign T58_59 = T65[61] | 1'b0;
  assign T58_58 = T65[60] | 1'b0;
  assign T59_57 = 1'b0 | T62_55;
  assign T59_56 = 1'b0 | T62_54;
  assign T58_55 = 1'b0 | T62_53;
  assign T58_54 = 1'b0 | T62_52;
  assign T59_53 = T63[59] | 1'b0;
  assign T59_52 = T63[58] | 1'b0;
  assign T58_51 = T63[57] | 1'b0;
  assign T58_50 = T63[56] | 1'b0;
  assign T59_49 = 1'b0 | T62_47;
  assign T59_48 = 1'b0 | T62_46;
  assign T58_47 = 1'b0 | T62_45;
  assign T58_46 = 1'b0 | T62_44;
  assign T59_45 = T63_51 | 1'b0;
  assign T59_44 = T63_50 | 1'b0;
  assign T58_43 = T63_49 | 1'b0;
  assign T58_42 = T63_48 | 1'b0;
  assign T59_41 = 1'b0 | T62_39;
  assign T59_40 = 1'b0 | T62_38;
  assign T58_39 = 1'b0 | T62_37;
  assign T58_38 = 1'b0 | T62_36;
  assign T59_37 = T63_43 | 1'b0;
  assign T59_36 = T63_42 | 1'b0;
  assign T58_35 = T63_41 | 1'b0;
  assign T58_34 = T63_40 | 1'b0;
  assign T59_33 = 1'b0 | T62_31;
  assign T59_32 = 1'b0 | T62_30;
  assign T58_31 = 1'b0 | T62_29;
  assign T58_30 = 1'b0 | T62_28;
  assign T59_29 = T63_35 | 1'b0;
  assign T59_28 = T63_34 | 1'b0;
  assign T58_27 = T63_33 | 1'b0;
  assign T58_26 = T63_32 | 1'b0;
  assign T59_25 = 1'b0 | T62_23;
  assign T59_24 = 1'b0 | T62_22;
  assign T58_23 = 1'b0 | T62_21;
  assign T58_22 = 1'b0 | T62_20;
  assign T59_21 = T63_27 | 1'b0;
  assign T59_20 = T63_26 | 1'b0;
  assign T58_19 = T63_25 | 1'b0;
  assign T58_18 = T63_24 | 1'b0;
  assign T59_17 = 1'b0 | T62_15;
  assign T59_16 = 1'b0 | T62_14;
  assign T58_15 = 1'b0 | T62_13;
  assign T58_14 = 1'b0 | T62_12;
  assign T59_13 = T63_19 | 1'b0;
  assign T59_12 = T63_18 | 1'b0;
  assign T58_11 = T63_17 | 1'b0;
  assign T58_10 = T63_16 | 1'b0;
  assign T59_9 = 1'b0 | T62_7;
  assign T59_8 = 1'b0 | T62_6;
  assign T58_7 = 1'b0 | T62_5;
  assign T58_6 = 1'b0 | T62_4;
  assign T59_5 = T63_11 | 1'b0;
  assign T59_4 = T63_10 | 1'b0;
  assign T58_3 = T63_9 | 1'b0;
  assign T58_2 = T63_8 | 1'b0;
  assign T65[63] = 1'b0 | T66[63];
  assign T65[62] = 1'b0 | T66[62];
  assign T65[61] = 1'b0 | T66[61];
  assign T65[60] = 1'b0 | T66[60];
  assign T62[63] = 1'b0 | T66[59];
  assign T62[62] = 1'b0 | T66[58];
  assign T62[61] = 1'b0 | T66[57];
  assign T62[60] = 1'b0 | T66[56];
  assign T63[59] = T69[63] | 1'b0;
  assign T63[58] = T69[62] | 1'b0;
  assign T63[57] = T69[61] | 1'b0;
  assign T63[56] = T69[60] | 1'b0;
  assign T62_55 = T69[59] | 1'b0;
  assign T62_54 = T69[58] | 1'b0;
  assign T62_53 = T69[57] | 1'b0;
  assign T62_52 = T69[56] | 1'b0;
  assign T63_51 = 1'b0 | T66_47;
  assign T63_50 = 1'b0 | T66_46;
  assign T63_49 = 1'b0 | T66_45;
  assign T63_48 = 1'b0 | T66_44;
  assign T62_47 = 1'b0 | T66_43;
  assign T62_46 = 1'b0 | T66_42;
  assign T62_45 = 1'b0 | T66_41;
  assign T62_44 = 1'b0 | T66_40;
  assign T63_43 = T67[55] | 1'b0;
  assign T63_42 = T67[54] | 1'b0;
  assign T63_41 = T67[53] | 1'b0;
  assign T63_40 = T67[52] | 1'b0;
  assign T62_39 = T67[51] | 1'b0;
  assign T62_38 = T67[50] | 1'b0;
  assign T62_37 = T67[49] | 1'b0;
  assign T62_36 = T67[48] | 1'b0;
  assign T63_35 = 1'b0 | T66_31;
  assign T63_34 = 1'b0 | T66_30;
  assign T63_33 = 1'b0 | T66_29;
  assign T63_32 = 1'b0 | T66_28;
  assign T62_31 = 1'b0 | T66_27;
  assign T62_30 = 1'b0 | T66_26;
  assign T62_29 = 1'b0 | T66_25;
  assign T62_28 = 1'b0 | T66_24;
  assign T63_27 = T67_39 | 1'b0;
  assign T63_26 = T67_38 | 1'b0;
  assign T63_25 = T67_37 | 1'b0;
  assign T63_24 = T67_36 | 1'b0;
  assign T62_23 = T67_35 | 1'b0;
  assign T62_22 = T67_34 | 1'b0;
  assign T62_21 = T67_33 | 1'b0;
  assign T62_20 = T67_32 | 1'b0;
  assign T63_19 = 1'b0 | T66_15;
  assign T63_18 = 1'b0 | T66_14;
  assign T63_17 = 1'b0 | T66_13;
  assign T63_16 = 1'b0 | T66_12;
  assign T62_15 = 1'b0 | T66_11;
  assign T62_14 = 1'b0 | T66_10;
  assign T62_13 = 1'b0 | T66_9;
  assign T62_12 = 1'b0 | T66_8;
  assign T63_11 = T67_23 | 1'b0;
  assign T63_10 = T67_22 | 1'b0;
  assign T63_9 = T67_21 | 1'b0;
  assign T63_8 = T67_20 | 1'b0;
  assign T62_7 = T67_19 | 1'b0;
  assign T62_6 = T67_18 | 1'b0;
  assign T62_5 = T67_17 | 1'b0;
  assign T62_4 = T67_16 | 1'b0;
  assign T69[63] = 1'b0 | T70[63];
  assign T69[62] = 1'b0 | T70[62];
  assign T69[61] = 1'b0 | T70[61];
  assign T69[60] = 1'b0 | T70[60];
  assign T69[59] = 1'b0 | T70[59];
  assign T69[58] = 1'b0 | T70[58];
  assign T69[57] = 1'b0 | T70[57];
  assign T69[56] = 1'b0 | T70[56];
  assign T66[63] = 1'b0 | T70[55];
  assign T66[62] = 1'b0 | T70[54];
  assign T66[61] = 1'b0 | T70[53];
  assign T66[60] = 1'b0 | T70[52];
  assign T66[59] = 1'b0 | T70[51];
  assign T66[58] = 1'b0 | T70[50];
  assign T66[57] = 1'b0 | T70[49];
  assign T66[56] = 1'b0 | T70[48];
  assign T67[55] = T73[63] | 1'b0;
  assign T67[54] = T73[62] | 1'b0;
  assign T67[53] = T73[61] | 1'b0;
  assign T67[52] = T73[60] | 1'b0;
  assign T67[51] = T73[59] | 1'b0;
  assign T67[50] = T73[58] | 1'b0;
  assign T67[49] = T73[57] | 1'b0;
  assign T67[48] = T73[56] | 1'b0;
  assign T66_47 = T73[55] | 1'b0;
  assign T66_46 = T73[54] | 1'b0;
  assign T66_45 = T73[53] | 1'b0;
  assign T66_44 = T73[52] | 1'b0;
  assign T66_43 = T73[51] | 1'b0;
  assign T66_42 = T73[50] | 1'b0;
  assign T66_41 = T73[49] | 1'b0;
  assign T66_40 = T73[48] | 1'b0;
  assign T67_39 = 1'b0 | T70_31;
  assign T67_38 = 1'b0 | T70_30;
  assign T67_37 = 1'b0 | T70_29;
  assign T67_36 = 1'b0 | T70_28;
  assign T67_35 = 1'b0 | T70_27;
  assign T67_34 = 1'b0 | T70_26;
  assign T67_33 = 1'b0 | T70_25;
  assign T67_32 = 1'b0 | T70_24;
  assign T66_31 = 1'b0 | T70_23;
  assign T66_30 = 1'b0 | T70_22;
  assign T66_29 = 1'b0 | T70_21;
  assign T66_28 = 1'b0 | T70_20;
  assign T66_27 = 1'b0 | T70_19;
  assign T66_26 = 1'b0 | T70_18;
  assign T66_25 = 1'b0 | T70_17;
  assign T66_24 = 1'b0 | T70_16;
  assign T67_23 = T71[47] | 1'b0;
  assign T67_22 = T71[46] | 1'b0;
  assign T67_21 = T71[45] | 1'b0;
  assign T67_20 = T71[44] | 1'b0;
  assign T67_19 = T71[43] | 1'b0;
  assign T67_18 = T71[42] | 1'b0;
  assign T67_17 = T71[41] | 1'b0;
  assign T67_16 = T71[40] | 1'b0;
  assign T66_15 = T71[39] | 1'b0;
  assign T66_14 = T71[38] | 1'b0;
  assign T66_13 = T71[37] | 1'b0;
  assign T66_12 = T71[36] | 1'b0;
  assign T66_11 = T71[35] | 1'b0;
  assign T66_10 = T71[34] | 1'b0;
  assign T66_9 = T71[33] | 1'b0;
  assign T66_8 = T71[32] | 1'b0;
  assign T73[63] = 1'b0 | io_in1[31];
  assign T73[62] = 1'b0 | io_in1[30];
  assign T73[61] = 1'b0 | io_in1[29];
  assign T73[60] = 1'b0 | io_in1[28];
  assign T73[59] = 1'b0 | io_in1[27];
  assign T73[58] = 1'b0 | io_in1[26];
  assign T73[57] = 1'b0 | io_in1[25];
  assign T73[56] = 1'b0 | io_in1[24];
  assign T73[55] = 1'b0 | io_in1[23];
  assign T73[54] = 1'b0 | io_in1[22];
  assign T73[53] = 1'b0 | io_in1[21];
  assign T73[52] = 1'b0 | io_in1[20];
  assign T73[51] = 1'b0 | io_in1[19];
  assign T73[50] = 1'b0 | io_in1[18];
  assign T73[49] = 1'b0 | io_in1[17];
  assign T73[48] = 1'b0 | io_in1[16];
  assign T70[63] = 1'b0 | io_in1[15];
  assign T70[62] = 1'b0 | io_in1[14];
  assign T70[61] = 1'b0 | io_in1[13];
  assign T70[60] = 1'b0 | io_in1[12];
  assign T70[59] = 1'b0 | io_in1[11];
  assign T70[58] = 1'b0 | io_in1[10];
  assign T70[57] = 1'b0 | io_in1[9];
  assign T70[56] = 1'b0 | io_in1[8];
  assign T70[55] = 1'b0 | io_in1[7];
  assign T70[54] = 1'b0 | io_in1[6];
  assign T70[53] = 1'b0 | io_in1[5];
  assign T70[52] = 1'b0 | io_in1[4];
  assign T70[51] = 1'b0 | io_in1[3];
  assign T70[50] = 1'b0 | io_in1[2];
  assign T70[49] = 1'b0 | io_in1[1];
  assign T70[48] = 1'b0 | io_in1[0];
  assign T71[47] = T77[31] | 1'b0;
  assign T71[46] = T77[30] | 1'b0;
  assign T71[45] = T77[29] | 1'b0;
  assign T71[44] = T77[28] | 1'b0;
  assign T71[43] = T77[27] | 1'b0;
  assign T71[42] = T77[26] | 1'b0;
  assign T71[41] = T77[25] | 1'b0;
  assign T71[40] = T77[24] | 1'b0;
  assign T71[39] = T77[23] | 1'b0;
  assign T71[38] = T77[22] | 1'b0;
  assign T71[37] = T77[21] | 1'b0;
  assign T71[36] = T77[20] | 1'b0;
  assign T71[35] = T77[19] | 1'b0;
  assign T71[34] = T77[18] | 1'b0;
  assign T71[33] = T77[17] | 1'b0;
  assign T71[32] = T77[16] | 1'b0;
  assign T70_31 = T77[15] | 1'b0;
  assign T70_30 = T77[14] | 1'b0;
  assign T70_29 = T77[13] | 1'b0;
  assign T70_28 = T77[12] | 1'b0;
  assign T70_27 = T77[11] | 1'b0;
  assign T70_26 = T77[10] | 1'b0;
  assign T70_25 = T77[9] | 1'b0;
  assign T70_24 = T77[8] | 1'b0;
  assign T70_23 = T77[7] | 1'b0;
  assign T70_22 = T77[6] | 1'b0;
  assign T70_21 = T77[5] | 1'b0;
  assign T70_20 = T77[4] | 1'b0;
  assign T70_19 = T77[3] | 1'b0;
  assign T70_18 = T77[2] | 1'b0;
  assign T70_17 = T77[1] | 1'b0;
  assign T70_16 = T77[0] | 1'b0;
  assign T153[0] = io_fn[3] & io_in1[31];
  assign T98 = N117 | N119;
  assign T51[64] = io_fn[3] & T51[63];
  assign N27 = ~T118;
  assign T118 = N117 | N119;
  assign T121[63] = 1'b0 | lg[63];
  assign T121[62] = 1'b0 | lg[62];
  assign T121[61] = 1'b0 | lg[61];
  assign T121[60] = 1'b0 | lg[60];
  assign T121[59] = 1'b0 | lg[59];
  assign T121[58] = 1'b0 | lg[58];
  assign T121[57] = 1'b0 | lg[57];
  assign T121[56] = 1'b0 | lg[56];
  assign T121[55] = 1'b0 | lg[55];
  assign T121[54] = 1'b0 | lg[54];
  assign T121[53] = 1'b0 | lg[53];
  assign T121[52] = 1'b0 | lg[52];
  assign T121[51] = 1'b0 | lg[51];
  assign T121[50] = 1'b0 | lg[50];
  assign T121[49] = 1'b0 | lg[49];
  assign T121[48] = 1'b0 | lg[48];
  assign T121[47] = 1'b0 | lg[47];
  assign T121[46] = 1'b0 | lg[46];
  assign T121[45] = 1'b0 | lg[45];
  assign T121[44] = 1'b0 | lg[44];
  assign T121[43] = 1'b0 | lg[43];
  assign T121[42] = 1'b0 | lg[42];
  assign T121[41] = 1'b0 | lg[41];
  assign T121[40] = 1'b0 | lg[40];
  assign T121[39] = 1'b0 | lg[39];
  assign T121[38] = 1'b0 | lg[38];
  assign T121[37] = 1'b0 | lg[37];
  assign T121[36] = 1'b0 | lg[36];
  assign T121[35] = 1'b0 | lg[35];
  assign T121[34] = 1'b0 | lg[34];
  assign T121[33] = 1'b0 | lg[33];
  assign T121[32] = 1'b0 | lg[32];
  assign T121[31] = 1'b0 | lg[31];
  assign T121[30] = 1'b0 | lg[30];
  assign T121[29] = 1'b0 | lg[29];
  assign T121[28] = 1'b0 | lg[28];
  assign T121[27] = 1'b0 | lg[27];
  assign T121[26] = 1'b0 | lg[26];
  assign T121[25] = 1'b0 | lg[25];
  assign T121[24] = 1'b0 | lg[24];
  assign T121[23] = 1'b0 | lg[23];
  assign T121[22] = 1'b0 | lg[22];
  assign T121[21] = 1'b0 | lg[21];
  assign T121[20] = 1'b0 | lg[20];
  assign T121[19] = 1'b0 | lg[19];
  assign T121[18] = 1'b0 | lg[18];
  assign T121[17] = 1'b0 | lg[17];
  assign T121[16] = 1'b0 | lg[16];
  assign T121[15] = 1'b0 | lg[15];
  assign T121[14] = 1'b0 | lg[14];
  assign T121[13] = 1'b0 | lg[13];
  assign T121[12] = 1'b0 | lg[12];
  assign T121[11] = 1'b0 | lg[11];
  assign T121[10] = 1'b0 | lg[10];
  assign T121[9] = 1'b0 | lg[9];
  assign T121[8] = 1'b0 | lg[8];
  assign T121[7] = 1'b0 | lg[7];
  assign T121[6] = 1'b0 | lg[6];
  assign T121[5] = 1'b0 | lg[5];
  assign T121[4] = 1'b0 | lg[4];
  assign T121[3] = 1'b0 | lg[3];
  assign T121[2] = 1'b0 | lg[2];
  assign T121[1] = 1'b0 | lg[1];
  assign T121[0] = T160[0] | lg[0];
  assign lg[63] = T127[63] | T122[63];
  assign lg[62] = T127[62] | T122[62];
  assign lg[61] = T127[61] | T122[61];
  assign lg[60] = T127[60] | T122[60];
  assign lg[59] = T127[59] | T122[59];
  assign lg[58] = T127[58] | T122[58];
  assign lg[57] = T127[57] | T122[57];
  assign lg[56] = T127[56] | T122[56];
  assign lg[55] = T127[55] | T122[55];
  assign lg[54] = T127[54] | T122[54];
  assign lg[53] = T127[53] | T122[53];
  assign lg[52] = T127[52] | T122[52];
  assign lg[51] = T127[51] | T122[51];
  assign lg[50] = T127[50] | T122[50];
  assign lg[49] = T127[49] | T122[49];
  assign lg[48] = T127[48] | T122[48];
  assign lg[47] = T127[47] | T122[47];
  assign lg[46] = T127[46] | T122[46];
  assign lg[45] = T127[45] | T122[45];
  assign lg[44] = T127[44] | T122[44];
  assign lg[43] = T127[43] | T122[43];
  assign lg[42] = T127[42] | T122[42];
  assign lg[41] = T127[41] | T122[41];
  assign lg[40] = T127[40] | T122[40];
  assign lg[39] = T127[39] | T122[39];
  assign lg[38] = T127[38] | T122[38];
  assign lg[37] = T127[37] | T122[37];
  assign lg[36] = T127[36] | T122[36];
  assign lg[35] = T127[35] | T122[35];
  assign lg[34] = T127[34] | T122[34];
  assign lg[33] = T127[33] | T122[33];
  assign lg[32] = T127[32] | T122[32];
  assign lg[31] = T127[31] | T122[31];
  assign lg[30] = T127[30] | T122[30];
  assign lg[29] = T127[29] | T122[29];
  assign lg[28] = T127[28] | T122[28];
  assign lg[27] = T127[27] | T122[27];
  assign lg[26] = T127[26] | T122[26];
  assign lg[25] = T127[25] | T122[25];
  assign lg[24] = T127[24] | T122[24];
  assign lg[23] = T127[23] | T122[23];
  assign lg[22] = T127[22] | T122[22];
  assign lg[21] = T127[21] | T122[21];
  assign lg[20] = T127[20] | T122[20];
  assign lg[19] = T127[19] | T122[19];
  assign lg[18] = T127[18] | T122[18];
  assign lg[17] = T127[17] | T122[17];
  assign lg[16] = T127[16] | T122[16];
  assign lg[15] = T127[15] | T122[15];
  assign lg[14] = T127[14] | T122[14];
  assign lg[13] = T127[13] | T122[13];
  assign lg[12] = T127[12] | T122[12];
  assign lg[11] = T127[11] | T122[11];
  assign lg[10] = T127[10] | T122[10];
  assign lg[9] = T127[9] | T122[9];
  assign lg[8] = T127[8] | T122[8];
  assign lg[7] = T127[7] | T122[7];
  assign lg[6] = T127[6] | T122[6];
  assign lg[5] = T127[5] | T122[5];
  assign lg[4] = T127[4] | T122[4];
  assign lg[3] = T127[3] | T122[3];
  assign lg[2] = T127[2] | T122[2];
  assign lg[1] = T127[1] | T122[1];
  assign lg[0] = T127[0] | T122[0];
  assign N28 = ~T124;
  assign T123[63] = io_in1[63] & io_in2[63];
  assign T123[62] = io_in1[62] & io_in2[62];
  assign T123[61] = io_in1[61] & io_in2[61];
  assign T123[60] = io_in1[60] & io_in2[60];
  assign T123[59] = io_in1[59] & io_in2[59];
  assign T123[58] = io_in1[58] & io_in2[58];
  assign T123[57] = io_in1[57] & io_in2[57];
  assign T123[56] = io_in1[56] & io_in2[56];
  assign T123[55] = io_in1[55] & io_in2[55];
  assign T123[54] = io_in1[54] & io_in2[54];
  assign T123[53] = io_in1[53] & io_in2[53];
  assign T123[52] = io_in1[52] & io_in2[52];
  assign T123[51] = io_in1[51] & io_in2[51];
  assign T123[50] = io_in1[50] & io_in2[50];
  assign T123[49] = io_in1[49] & io_in2[49];
  assign T123[48] = io_in1[48] & io_in2[48];
  assign T123[47] = io_in1[47] & io_in2[47];
  assign T123[46] = io_in1[46] & io_in2[46];
  assign T123[45] = io_in1[45] & io_in2[45];
  assign T123[44] = io_in1[44] & io_in2[44];
  assign T123[43] = io_in1[43] & io_in2[43];
  assign T123[42] = io_in1[42] & io_in2[42];
  assign T123[41] = io_in1[41] & io_in2[41];
  assign T123[40] = io_in1[40] & io_in2[40];
  assign T123[39] = io_in1[39] & io_in2[39];
  assign T123[38] = io_in1[38] & io_in2[38];
  assign T123[37] = io_in1[37] & io_in2[37];
  assign T123[36] = io_in1[36] & io_in2[36];
  assign T123[35] = io_in1[35] & io_in2[35];
  assign T123[34] = io_in1[34] & io_in2[34];
  assign T123[33] = io_in1[33] & io_in2[33];
  assign T123[32] = io_in1[32] & io_in2[32];
  assign T123[31] = io_in1[31] & io_in2[31];
  assign T123[30] = io_in1[30] & io_in2[30];
  assign T123[29] = io_in1[29] & io_in2[29];
  assign T123[28] = io_in1[28] & io_in2[28];
  assign T123[27] = io_in1[27] & io_in2[27];
  assign T123[26] = io_in1[26] & io_in2[26];
  assign T123[25] = io_in1[25] & io_in2[25];
  assign T123[24] = io_in1[24] & io_in2[24];
  assign T123[23] = io_in1[23] & io_in2[23];
  assign T123[22] = io_in1[22] & io_in2[22];
  assign T123[21] = io_in1[21] & io_in2[21];
  assign T123[20] = io_in1[20] & io_in2[20];
  assign T123[19] = io_in1[19] & io_in2[19];
  assign T123[18] = io_in1[18] & io_in2[18];
  assign T123[17] = io_in1[17] & io_in2[17];
  assign T123[16] = io_in1[16] & io_in2[16];
  assign T123[15] = io_in1[15] & io_in2[15];
  assign T123[14] = io_in1[14] & io_in2[14];
  assign T123[13] = io_in1[13] & io_in2[13];
  assign T123[12] = io_in1[12] & io_in2[12];
  assign T123[11] = io_in1[11] & io_in2[11];
  assign T123[10] = io_in1[10] & io_in2[10];
  assign T123[9] = io_in1[9] & io_in2[9];
  assign T123[8] = io_in1[8] & io_in2[8];
  assign T123[7] = io_in1[7] & io_in2[7];
  assign T123[6] = io_in1[6] & io_in2[6];
  assign T123[5] = io_in1[5] & io_in2[5];
  assign T123[4] = io_in1[4] & io_in2[4];
  assign T123[3] = io_in1[3] & io_in2[3];
  assign T123[2] = io_in1[2] & io_in2[2];
  assign T123[1] = io_in1[1] & io_in2[1];
  assign T123[0] = io_in1[0] & io_in2[0];
  assign T124 = N124 | N126;
  assign N29 = ~T128;
  assign T128 = N121 | N124;
  assign T160[0] = T132 & io_cmp_out;
  assign T132 = T134 | T133;
  assign T134 = N43 | N46;
  assign T137 = N34 | N40;

endmodule