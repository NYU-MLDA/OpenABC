module bsg_mem_1r1w_synth_width_p101_els_p8_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [100:0] w_data_i;
  input [2:0] r_addr_i;
  output [100:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [100:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53;
  wire [807:0] mem;
  reg mem_807_sv2v_reg,mem_806_sv2v_reg,mem_805_sv2v_reg,mem_804_sv2v_reg,
  mem_803_sv2v_reg,mem_802_sv2v_reg,mem_801_sv2v_reg,mem_800_sv2v_reg,mem_799_sv2v_reg,
  mem_798_sv2v_reg,mem_797_sv2v_reg,mem_796_sv2v_reg,mem_795_sv2v_reg,mem_794_sv2v_reg,
  mem_793_sv2v_reg,mem_792_sv2v_reg,mem_791_sv2v_reg,mem_790_sv2v_reg,
  mem_789_sv2v_reg,mem_788_sv2v_reg,mem_787_sv2v_reg,mem_786_sv2v_reg,mem_785_sv2v_reg,
  mem_784_sv2v_reg,mem_783_sv2v_reg,mem_782_sv2v_reg,mem_781_sv2v_reg,mem_780_sv2v_reg,
  mem_779_sv2v_reg,mem_778_sv2v_reg,mem_777_sv2v_reg,mem_776_sv2v_reg,
  mem_775_sv2v_reg,mem_774_sv2v_reg,mem_773_sv2v_reg,mem_772_sv2v_reg,mem_771_sv2v_reg,
  mem_770_sv2v_reg,mem_769_sv2v_reg,mem_768_sv2v_reg,mem_767_sv2v_reg,mem_766_sv2v_reg,
  mem_765_sv2v_reg,mem_764_sv2v_reg,mem_763_sv2v_reg,mem_762_sv2v_reg,mem_761_sv2v_reg,
  mem_760_sv2v_reg,mem_759_sv2v_reg,mem_758_sv2v_reg,mem_757_sv2v_reg,
  mem_756_sv2v_reg,mem_755_sv2v_reg,mem_754_sv2v_reg,mem_753_sv2v_reg,mem_752_sv2v_reg,
  mem_751_sv2v_reg,mem_750_sv2v_reg,mem_749_sv2v_reg,mem_748_sv2v_reg,mem_747_sv2v_reg,
  mem_746_sv2v_reg,mem_745_sv2v_reg,mem_744_sv2v_reg,mem_743_sv2v_reg,
  mem_742_sv2v_reg,mem_741_sv2v_reg,mem_740_sv2v_reg,mem_739_sv2v_reg,mem_738_sv2v_reg,
  mem_737_sv2v_reg,mem_736_sv2v_reg,mem_735_sv2v_reg,mem_734_sv2v_reg,mem_733_sv2v_reg,
  mem_732_sv2v_reg,mem_731_sv2v_reg,mem_730_sv2v_reg,mem_729_sv2v_reg,mem_728_sv2v_reg,
  mem_727_sv2v_reg,mem_726_sv2v_reg,mem_725_sv2v_reg,mem_724_sv2v_reg,
  mem_723_sv2v_reg,mem_722_sv2v_reg,mem_721_sv2v_reg,mem_720_sv2v_reg,mem_719_sv2v_reg,
  mem_718_sv2v_reg,mem_717_sv2v_reg,mem_716_sv2v_reg,mem_715_sv2v_reg,mem_714_sv2v_reg,
  mem_713_sv2v_reg,mem_712_sv2v_reg,mem_711_sv2v_reg,mem_710_sv2v_reg,
  mem_709_sv2v_reg,mem_708_sv2v_reg,mem_707_sv2v_reg,mem_706_sv2v_reg,mem_705_sv2v_reg,
  mem_704_sv2v_reg,mem_703_sv2v_reg,mem_702_sv2v_reg,mem_701_sv2v_reg,mem_700_sv2v_reg,
  mem_699_sv2v_reg,mem_698_sv2v_reg,mem_697_sv2v_reg,mem_696_sv2v_reg,
  mem_695_sv2v_reg,mem_694_sv2v_reg,mem_693_sv2v_reg,mem_692_sv2v_reg,mem_691_sv2v_reg,
  mem_690_sv2v_reg,mem_689_sv2v_reg,mem_688_sv2v_reg,mem_687_sv2v_reg,mem_686_sv2v_reg,
  mem_685_sv2v_reg,mem_684_sv2v_reg,mem_683_sv2v_reg,mem_682_sv2v_reg,mem_681_sv2v_reg,
  mem_680_sv2v_reg,mem_679_sv2v_reg,mem_678_sv2v_reg,mem_677_sv2v_reg,
  mem_676_sv2v_reg,mem_675_sv2v_reg,mem_674_sv2v_reg,mem_673_sv2v_reg,mem_672_sv2v_reg,
  mem_671_sv2v_reg,mem_670_sv2v_reg,mem_669_sv2v_reg,mem_668_sv2v_reg,mem_667_sv2v_reg,
  mem_666_sv2v_reg,mem_665_sv2v_reg,mem_664_sv2v_reg,mem_663_sv2v_reg,
  mem_662_sv2v_reg,mem_661_sv2v_reg,mem_660_sv2v_reg,mem_659_sv2v_reg,mem_658_sv2v_reg,
  mem_657_sv2v_reg,mem_656_sv2v_reg,mem_655_sv2v_reg,mem_654_sv2v_reg,mem_653_sv2v_reg,
  mem_652_sv2v_reg,mem_651_sv2v_reg,mem_650_sv2v_reg,mem_649_sv2v_reg,mem_648_sv2v_reg,
  mem_647_sv2v_reg,mem_646_sv2v_reg,mem_645_sv2v_reg,mem_644_sv2v_reg,
  mem_643_sv2v_reg,mem_642_sv2v_reg,mem_641_sv2v_reg,mem_640_sv2v_reg,mem_639_sv2v_reg,
  mem_638_sv2v_reg,mem_637_sv2v_reg,mem_636_sv2v_reg,mem_635_sv2v_reg,mem_634_sv2v_reg,
  mem_633_sv2v_reg,mem_632_sv2v_reg,mem_631_sv2v_reg,mem_630_sv2v_reg,
  mem_629_sv2v_reg,mem_628_sv2v_reg,mem_627_sv2v_reg,mem_626_sv2v_reg,mem_625_sv2v_reg,
  mem_624_sv2v_reg,mem_623_sv2v_reg,mem_622_sv2v_reg,mem_621_sv2v_reg,mem_620_sv2v_reg,
  mem_619_sv2v_reg,mem_618_sv2v_reg,mem_617_sv2v_reg,mem_616_sv2v_reg,
  mem_615_sv2v_reg,mem_614_sv2v_reg,mem_613_sv2v_reg,mem_612_sv2v_reg,mem_611_sv2v_reg,
  mem_610_sv2v_reg,mem_609_sv2v_reg,mem_608_sv2v_reg,mem_607_sv2v_reg,mem_606_sv2v_reg,
  mem_605_sv2v_reg,mem_604_sv2v_reg,mem_603_sv2v_reg,mem_602_sv2v_reg,mem_601_sv2v_reg,
  mem_600_sv2v_reg,mem_599_sv2v_reg,mem_598_sv2v_reg,mem_597_sv2v_reg,
  mem_596_sv2v_reg,mem_595_sv2v_reg,mem_594_sv2v_reg,mem_593_sv2v_reg,mem_592_sv2v_reg,
  mem_591_sv2v_reg,mem_590_sv2v_reg,mem_589_sv2v_reg,mem_588_sv2v_reg,mem_587_sv2v_reg,
  mem_586_sv2v_reg,mem_585_sv2v_reg,mem_584_sv2v_reg,mem_583_sv2v_reg,
  mem_582_sv2v_reg,mem_581_sv2v_reg,mem_580_sv2v_reg,mem_579_sv2v_reg,mem_578_sv2v_reg,
  mem_577_sv2v_reg,mem_576_sv2v_reg,mem_575_sv2v_reg,mem_574_sv2v_reg,mem_573_sv2v_reg,
  mem_572_sv2v_reg,mem_571_sv2v_reg,mem_570_sv2v_reg,mem_569_sv2v_reg,mem_568_sv2v_reg,
  mem_567_sv2v_reg,mem_566_sv2v_reg,mem_565_sv2v_reg,mem_564_sv2v_reg,
  mem_563_sv2v_reg,mem_562_sv2v_reg,mem_561_sv2v_reg,mem_560_sv2v_reg,mem_559_sv2v_reg,
  mem_558_sv2v_reg,mem_557_sv2v_reg,mem_556_sv2v_reg,mem_555_sv2v_reg,mem_554_sv2v_reg,
  mem_553_sv2v_reg,mem_552_sv2v_reg,mem_551_sv2v_reg,mem_550_sv2v_reg,
  mem_549_sv2v_reg,mem_548_sv2v_reg,mem_547_sv2v_reg,mem_546_sv2v_reg,mem_545_sv2v_reg,
  mem_544_sv2v_reg,mem_543_sv2v_reg,mem_542_sv2v_reg,mem_541_sv2v_reg,mem_540_sv2v_reg,
  mem_539_sv2v_reg,mem_538_sv2v_reg,mem_537_sv2v_reg,mem_536_sv2v_reg,
  mem_535_sv2v_reg,mem_534_sv2v_reg,mem_533_sv2v_reg,mem_532_sv2v_reg,mem_531_sv2v_reg,
  mem_530_sv2v_reg,mem_529_sv2v_reg,mem_528_sv2v_reg,mem_527_sv2v_reg,mem_526_sv2v_reg,
  mem_525_sv2v_reg,mem_524_sv2v_reg,mem_523_sv2v_reg,mem_522_sv2v_reg,mem_521_sv2v_reg,
  mem_520_sv2v_reg,mem_519_sv2v_reg,mem_518_sv2v_reg,mem_517_sv2v_reg,
  mem_516_sv2v_reg,mem_515_sv2v_reg,mem_514_sv2v_reg,mem_513_sv2v_reg,mem_512_sv2v_reg,
  mem_511_sv2v_reg,mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,mem_507_sv2v_reg,
  mem_506_sv2v_reg,mem_505_sv2v_reg,mem_504_sv2v_reg,mem_503_sv2v_reg,
  mem_502_sv2v_reg,mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,mem_498_sv2v_reg,
  mem_497_sv2v_reg,mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,mem_493_sv2v_reg,
  mem_492_sv2v_reg,mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,mem_488_sv2v_reg,
  mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,mem_484_sv2v_reg,
  mem_483_sv2v_reg,mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,mem_479_sv2v_reg,
  mem_478_sv2v_reg,mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,mem_474_sv2v_reg,
  mem_473_sv2v_reg,mem_472_sv2v_reg,mem_471_sv2v_reg,mem_470_sv2v_reg,
  mem_469_sv2v_reg,mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,mem_465_sv2v_reg,
  mem_464_sv2v_reg,mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,mem_460_sv2v_reg,
  mem_459_sv2v_reg,mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,
  mem_455_sv2v_reg,mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,mem_451_sv2v_reg,
  mem_450_sv2v_reg,mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,mem_446_sv2v_reg,
  mem_445_sv2v_reg,mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,mem_441_sv2v_reg,
  mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,
  mem_436_sv2v_reg,mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,
  mem_431_sv2v_reg,mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,mem_427_sv2v_reg,
  mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,mem_423_sv2v_reg,
  mem_422_sv2v_reg,mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,
  mem_417_sv2v_reg,mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,mem_413_sv2v_reg,
  mem_412_sv2v_reg,mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,mem_408_sv2v_reg,
  mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,
  mem_403_sv2v_reg,mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,mem_399_sv2v_reg,
  mem_398_sv2v_reg,mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,mem_394_sv2v_reg,
  mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,mem_390_sv2v_reg,
  mem_389_sv2v_reg,mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,
  mem_384_sv2v_reg,mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,mem_380_sv2v_reg,
  mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,
  mem_375_sv2v_reg,mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,
  mem_370_sv2v_reg,mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,mem_366_sv2v_reg,
  mem_365_sv2v_reg,mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,mem_361_sv2v_reg,
  mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,
  mem_356_sv2v_reg,mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,
  mem_351_sv2v_reg,mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,mem_347_sv2v_reg,
  mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,mem_343_sv2v_reg,
  mem_342_sv2v_reg,mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,
  mem_337_sv2v_reg,mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,mem_333_sv2v_reg,
  mem_332_sv2v_reg,mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,mem_328_sv2v_reg,
  mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,
  mem_323_sv2v_reg,mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,mem_319_sv2v_reg,
  mem_318_sv2v_reg,mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,mem_314_sv2v_reg,
  mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,mem_310_sv2v_reg,
  mem_309_sv2v_reg,mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,
  mem_304_sv2v_reg,mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,mem_300_sv2v_reg,
  mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,
  mem_295_sv2v_reg,mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,
  mem_290_sv2v_reg,mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,mem_286_sv2v_reg,
  mem_285_sv2v_reg,mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,mem_281_sv2v_reg,
  mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,
  mem_276_sv2v_reg,mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,
  mem_271_sv2v_reg,mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,mem_267_sv2v_reg,
  mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,mem_263_sv2v_reg,
  mem_262_sv2v_reg,mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,
  mem_257_sv2v_reg,mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,mem_253_sv2v_reg,
  mem_252_sv2v_reg,mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,mem_248_sv2v_reg,
  mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,
  mem_243_sv2v_reg,mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,mem_239_sv2v_reg,
  mem_238_sv2v_reg,mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,mem_234_sv2v_reg,
  mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,
  mem_229_sv2v_reg,mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,
  mem_224_sv2v_reg,mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,mem_220_sv2v_reg,
  mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,
  mem_215_sv2v_reg,mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,
  mem_210_sv2v_reg,mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,mem_206_sv2v_reg,
  mem_205_sv2v_reg,mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,mem_201_sv2v_reg,
  mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,
  mem_196_sv2v_reg,mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,
  mem_191_sv2v_reg,mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,mem_187_sv2v_reg,
  mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,
  mem_182_sv2v_reg,mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,
  mem_177_sv2v_reg,mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,mem_173_sv2v_reg,
  mem_172_sv2v_reg,mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,mem_168_sv2v_reg,
  mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,
  mem_163_sv2v_reg,mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,mem_159_sv2v_reg,
  mem_158_sv2v_reg,mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,mem_154_sv2v_reg,
  mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,
  mem_149_sv2v_reg,mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,
  mem_144_sv2v_reg,mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,mem_140_sv2v_reg,
  mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,
  mem_135_sv2v_reg,mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,
  mem_130_sv2v_reg,mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,mem_126_sv2v_reg,
  mem_125_sv2v_reg,mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,mem_121_sv2v_reg,
  mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,
  mem_116_sv2v_reg,mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,
  mem_111_sv2v_reg,mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,mem_107_sv2v_reg,
  mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,
  mem_102_sv2v_reg,mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,
  mem_97_sv2v_reg,mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,
  mem_92_sv2v_reg,mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,
  mem_87_sv2v_reg,mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,
  mem_82_sv2v_reg,mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,
  mem_77_sv2v_reg,mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,
  mem_72_sv2v_reg,mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,
  mem_67_sv2v_reg,mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,
  mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,
  mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,
  mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,
  mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,
  mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,
  mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,
  mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,
  mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,
  mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,
  mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,
  mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,
  mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,
  mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[100] = (N17)? mem[100] : 
                         (N19)? mem[201] : 
                         (N21)? mem[302] : 
                         (N23)? mem[403] : 
                         (N18)? mem[504] : 
                         (N20)? mem[605] : 
                         (N22)? mem[706] : 
                         (N24)? mem[807] : 1'b0;
  assign r_data_o[99] = (N17)? mem[99] : 
                        (N19)? mem[200] : 
                        (N21)? mem[301] : 
                        (N23)? mem[402] : 
                        (N18)? mem[503] : 
                        (N20)? mem[604] : 
                        (N22)? mem[705] : 
                        (N24)? mem[806] : 1'b0;
  assign r_data_o[98] = (N17)? mem[98] : 
                        (N19)? mem[199] : 
                        (N21)? mem[300] : 
                        (N23)? mem[401] : 
                        (N18)? mem[502] : 
                        (N20)? mem[603] : 
                        (N22)? mem[704] : 
                        (N24)? mem[805] : 1'b0;
  assign r_data_o[97] = (N17)? mem[97] : 
                        (N19)? mem[198] : 
                        (N21)? mem[299] : 
                        (N23)? mem[400] : 
                        (N18)? mem[501] : 
                        (N20)? mem[602] : 
                        (N22)? mem[703] : 
                        (N24)? mem[804] : 1'b0;
  assign r_data_o[96] = (N17)? mem[96] : 
                        (N19)? mem[197] : 
                        (N21)? mem[298] : 
                        (N23)? mem[399] : 
                        (N18)? mem[500] : 
                        (N20)? mem[601] : 
                        (N22)? mem[702] : 
                        (N24)? mem[803] : 1'b0;
  assign r_data_o[95] = (N17)? mem[95] : 
                        (N19)? mem[196] : 
                        (N21)? mem[297] : 
                        (N23)? mem[398] : 
                        (N18)? mem[499] : 
                        (N20)? mem[600] : 
                        (N22)? mem[701] : 
                        (N24)? mem[802] : 1'b0;
  assign r_data_o[94] = (N17)? mem[94] : 
                        (N19)? mem[195] : 
                        (N21)? mem[296] : 
                        (N23)? mem[397] : 
                        (N18)? mem[498] : 
                        (N20)? mem[599] : 
                        (N22)? mem[700] : 
                        (N24)? mem[801] : 1'b0;
  assign r_data_o[93] = (N17)? mem[93] : 
                        (N19)? mem[194] : 
                        (N21)? mem[295] : 
                        (N23)? mem[396] : 
                        (N18)? mem[497] : 
                        (N20)? mem[598] : 
                        (N22)? mem[699] : 
                        (N24)? mem[800] : 1'b0;
  assign r_data_o[92] = (N17)? mem[92] : 
                        (N19)? mem[193] : 
                        (N21)? mem[294] : 
                        (N23)? mem[395] : 
                        (N18)? mem[496] : 
                        (N20)? mem[597] : 
                        (N22)? mem[698] : 
                        (N24)? mem[799] : 1'b0;
  assign r_data_o[91] = (N17)? mem[91] : 
                        (N19)? mem[192] : 
                        (N21)? mem[293] : 
                        (N23)? mem[394] : 
                        (N18)? mem[495] : 
                        (N20)? mem[596] : 
                        (N22)? mem[697] : 
                        (N24)? mem[798] : 1'b0;
  assign r_data_o[90] = (N17)? mem[90] : 
                        (N19)? mem[191] : 
                        (N21)? mem[292] : 
                        (N23)? mem[393] : 
                        (N18)? mem[494] : 
                        (N20)? mem[595] : 
                        (N22)? mem[696] : 
                        (N24)? mem[797] : 1'b0;
  assign r_data_o[89] = (N17)? mem[89] : 
                        (N19)? mem[190] : 
                        (N21)? mem[291] : 
                        (N23)? mem[392] : 
                        (N18)? mem[493] : 
                        (N20)? mem[594] : 
                        (N22)? mem[695] : 
                        (N24)? mem[796] : 1'b0;
  assign r_data_o[88] = (N17)? mem[88] : 
                        (N19)? mem[189] : 
                        (N21)? mem[290] : 
                        (N23)? mem[391] : 
                        (N18)? mem[492] : 
                        (N20)? mem[593] : 
                        (N22)? mem[694] : 
                        (N24)? mem[795] : 1'b0;
  assign r_data_o[87] = (N17)? mem[87] : 
                        (N19)? mem[188] : 
                        (N21)? mem[289] : 
                        (N23)? mem[390] : 
                        (N18)? mem[491] : 
                        (N20)? mem[592] : 
                        (N22)? mem[693] : 
                        (N24)? mem[794] : 1'b0;
  assign r_data_o[86] = (N17)? mem[86] : 
                        (N19)? mem[187] : 
                        (N21)? mem[288] : 
                        (N23)? mem[389] : 
                        (N18)? mem[490] : 
                        (N20)? mem[591] : 
                        (N22)? mem[692] : 
                        (N24)? mem[793] : 1'b0;
  assign r_data_o[85] = (N17)? mem[85] : 
                        (N19)? mem[186] : 
                        (N21)? mem[287] : 
                        (N23)? mem[388] : 
                        (N18)? mem[489] : 
                        (N20)? mem[590] : 
                        (N22)? mem[691] : 
                        (N24)? mem[792] : 1'b0;
  assign r_data_o[84] = (N17)? mem[84] : 
                        (N19)? mem[185] : 
                        (N21)? mem[286] : 
                        (N23)? mem[387] : 
                        (N18)? mem[488] : 
                        (N20)? mem[589] : 
                        (N22)? mem[690] : 
                        (N24)? mem[791] : 1'b0;
  assign r_data_o[83] = (N17)? mem[83] : 
                        (N19)? mem[184] : 
                        (N21)? mem[285] : 
                        (N23)? mem[386] : 
                        (N18)? mem[487] : 
                        (N20)? mem[588] : 
                        (N22)? mem[689] : 
                        (N24)? mem[790] : 1'b0;
  assign r_data_o[82] = (N17)? mem[82] : 
                        (N19)? mem[183] : 
                        (N21)? mem[284] : 
                        (N23)? mem[385] : 
                        (N18)? mem[486] : 
                        (N20)? mem[587] : 
                        (N22)? mem[688] : 
                        (N24)? mem[789] : 1'b0;
  assign r_data_o[81] = (N17)? mem[81] : 
                        (N19)? mem[182] : 
                        (N21)? mem[283] : 
                        (N23)? mem[384] : 
                        (N18)? mem[485] : 
                        (N20)? mem[586] : 
                        (N22)? mem[687] : 
                        (N24)? mem[788] : 1'b0;
  assign r_data_o[80] = (N17)? mem[80] : 
                        (N19)? mem[181] : 
                        (N21)? mem[282] : 
                        (N23)? mem[383] : 
                        (N18)? mem[484] : 
                        (N20)? mem[585] : 
                        (N22)? mem[686] : 
                        (N24)? mem[787] : 1'b0;
  assign r_data_o[79] = (N17)? mem[79] : 
                        (N19)? mem[180] : 
                        (N21)? mem[281] : 
                        (N23)? mem[382] : 
                        (N18)? mem[483] : 
                        (N20)? mem[584] : 
                        (N22)? mem[685] : 
                        (N24)? mem[786] : 1'b0;
  assign r_data_o[78] = (N17)? mem[78] : 
                        (N19)? mem[179] : 
                        (N21)? mem[280] : 
                        (N23)? mem[381] : 
                        (N18)? mem[482] : 
                        (N20)? mem[583] : 
                        (N22)? mem[684] : 
                        (N24)? mem[785] : 1'b0;
  assign r_data_o[77] = (N17)? mem[77] : 
                        (N19)? mem[178] : 
                        (N21)? mem[279] : 
                        (N23)? mem[380] : 
                        (N18)? mem[481] : 
                        (N20)? mem[582] : 
                        (N22)? mem[683] : 
                        (N24)? mem[784] : 1'b0;
  assign r_data_o[76] = (N17)? mem[76] : 
                        (N19)? mem[177] : 
                        (N21)? mem[278] : 
                        (N23)? mem[379] : 
                        (N18)? mem[480] : 
                        (N20)? mem[581] : 
                        (N22)? mem[682] : 
                        (N24)? mem[783] : 1'b0;
  assign r_data_o[75] = (N17)? mem[75] : 
                        (N19)? mem[176] : 
                        (N21)? mem[277] : 
                        (N23)? mem[378] : 
                        (N18)? mem[479] : 
                        (N20)? mem[580] : 
                        (N22)? mem[681] : 
                        (N24)? mem[782] : 1'b0;
  assign r_data_o[74] = (N17)? mem[74] : 
                        (N19)? mem[175] : 
                        (N21)? mem[276] : 
                        (N23)? mem[377] : 
                        (N18)? mem[478] : 
                        (N20)? mem[579] : 
                        (N22)? mem[680] : 
                        (N24)? mem[781] : 1'b0;
  assign r_data_o[73] = (N17)? mem[73] : 
                        (N19)? mem[174] : 
                        (N21)? mem[275] : 
                        (N23)? mem[376] : 
                        (N18)? mem[477] : 
                        (N20)? mem[578] : 
                        (N22)? mem[679] : 
                        (N24)? mem[780] : 1'b0;
  assign r_data_o[72] = (N17)? mem[72] : 
                        (N19)? mem[173] : 
                        (N21)? mem[274] : 
                        (N23)? mem[375] : 
                        (N18)? mem[476] : 
                        (N20)? mem[577] : 
                        (N22)? mem[678] : 
                        (N24)? mem[779] : 1'b0;
  assign r_data_o[71] = (N17)? mem[71] : 
                        (N19)? mem[172] : 
                        (N21)? mem[273] : 
                        (N23)? mem[374] : 
                        (N18)? mem[475] : 
                        (N20)? mem[576] : 
                        (N22)? mem[677] : 
                        (N24)? mem[778] : 1'b0;
  assign r_data_o[70] = (N17)? mem[70] : 
                        (N19)? mem[171] : 
                        (N21)? mem[272] : 
                        (N23)? mem[373] : 
                        (N18)? mem[474] : 
                        (N20)? mem[575] : 
                        (N22)? mem[676] : 
                        (N24)? mem[777] : 1'b0;
  assign r_data_o[69] = (N17)? mem[69] : 
                        (N19)? mem[170] : 
                        (N21)? mem[271] : 
                        (N23)? mem[372] : 
                        (N18)? mem[473] : 
                        (N20)? mem[574] : 
                        (N22)? mem[675] : 
                        (N24)? mem[776] : 1'b0;
  assign r_data_o[68] = (N17)? mem[68] : 
                        (N19)? mem[169] : 
                        (N21)? mem[270] : 
                        (N23)? mem[371] : 
                        (N18)? mem[472] : 
                        (N20)? mem[573] : 
                        (N22)? mem[674] : 
                        (N24)? mem[775] : 1'b0;
  assign r_data_o[67] = (N17)? mem[67] : 
                        (N19)? mem[168] : 
                        (N21)? mem[269] : 
                        (N23)? mem[370] : 
                        (N18)? mem[471] : 
                        (N20)? mem[572] : 
                        (N22)? mem[673] : 
                        (N24)? mem[774] : 1'b0;
  assign r_data_o[66] = (N17)? mem[66] : 
                        (N19)? mem[167] : 
                        (N21)? mem[268] : 
                        (N23)? mem[369] : 
                        (N18)? mem[470] : 
                        (N20)? mem[571] : 
                        (N22)? mem[672] : 
                        (N24)? mem[773] : 1'b0;
  assign r_data_o[65] = (N17)? mem[65] : 
                        (N19)? mem[166] : 
                        (N21)? mem[267] : 
                        (N23)? mem[368] : 
                        (N18)? mem[469] : 
                        (N20)? mem[570] : 
                        (N22)? mem[671] : 
                        (N24)? mem[772] : 1'b0;
  assign r_data_o[64] = (N17)? mem[64] : 
                        (N19)? mem[165] : 
                        (N21)? mem[266] : 
                        (N23)? mem[367] : 
                        (N18)? mem[468] : 
                        (N20)? mem[569] : 
                        (N22)? mem[670] : 
                        (N24)? mem[771] : 1'b0;
  assign r_data_o[63] = (N17)? mem[63] : 
                        (N19)? mem[164] : 
                        (N21)? mem[265] : 
                        (N23)? mem[366] : 
                        (N18)? mem[467] : 
                        (N20)? mem[568] : 
                        (N22)? mem[669] : 
                        (N24)? mem[770] : 1'b0;
  assign r_data_o[62] = (N17)? mem[62] : 
                        (N19)? mem[163] : 
                        (N21)? mem[264] : 
                        (N23)? mem[365] : 
                        (N18)? mem[466] : 
                        (N20)? mem[567] : 
                        (N22)? mem[668] : 
                        (N24)? mem[769] : 1'b0;
  assign r_data_o[61] = (N17)? mem[61] : 
                        (N19)? mem[162] : 
                        (N21)? mem[263] : 
                        (N23)? mem[364] : 
                        (N18)? mem[465] : 
                        (N20)? mem[566] : 
                        (N22)? mem[667] : 
                        (N24)? mem[768] : 1'b0;
  assign r_data_o[60] = (N17)? mem[60] : 
                        (N19)? mem[161] : 
                        (N21)? mem[262] : 
                        (N23)? mem[363] : 
                        (N18)? mem[464] : 
                        (N20)? mem[565] : 
                        (N22)? mem[666] : 
                        (N24)? mem[767] : 1'b0;
  assign r_data_o[59] = (N17)? mem[59] : 
                        (N19)? mem[160] : 
                        (N21)? mem[261] : 
                        (N23)? mem[362] : 
                        (N18)? mem[463] : 
                        (N20)? mem[564] : 
                        (N22)? mem[665] : 
                        (N24)? mem[766] : 1'b0;
  assign r_data_o[58] = (N17)? mem[58] : 
                        (N19)? mem[159] : 
                        (N21)? mem[260] : 
                        (N23)? mem[361] : 
                        (N18)? mem[462] : 
                        (N20)? mem[563] : 
                        (N22)? mem[664] : 
                        (N24)? mem[765] : 1'b0;
  assign r_data_o[57] = (N17)? mem[57] : 
                        (N19)? mem[158] : 
                        (N21)? mem[259] : 
                        (N23)? mem[360] : 
                        (N18)? mem[461] : 
                        (N20)? mem[562] : 
                        (N22)? mem[663] : 
                        (N24)? mem[764] : 1'b0;
  assign r_data_o[56] = (N17)? mem[56] : 
                        (N19)? mem[157] : 
                        (N21)? mem[258] : 
                        (N23)? mem[359] : 
                        (N18)? mem[460] : 
                        (N20)? mem[561] : 
                        (N22)? mem[662] : 
                        (N24)? mem[763] : 1'b0;
  assign r_data_o[55] = (N17)? mem[55] : 
                        (N19)? mem[156] : 
                        (N21)? mem[257] : 
                        (N23)? mem[358] : 
                        (N18)? mem[459] : 
                        (N20)? mem[560] : 
                        (N22)? mem[661] : 
                        (N24)? mem[762] : 1'b0;
  assign r_data_o[54] = (N17)? mem[54] : 
                        (N19)? mem[155] : 
                        (N21)? mem[256] : 
                        (N23)? mem[357] : 
                        (N18)? mem[458] : 
                        (N20)? mem[559] : 
                        (N22)? mem[660] : 
                        (N24)? mem[761] : 1'b0;
  assign r_data_o[53] = (N17)? mem[53] : 
                        (N19)? mem[154] : 
                        (N21)? mem[255] : 
                        (N23)? mem[356] : 
                        (N18)? mem[457] : 
                        (N20)? mem[558] : 
                        (N22)? mem[659] : 
                        (N24)? mem[760] : 1'b0;
  assign r_data_o[52] = (N17)? mem[52] : 
                        (N19)? mem[153] : 
                        (N21)? mem[254] : 
                        (N23)? mem[355] : 
                        (N18)? mem[456] : 
                        (N20)? mem[557] : 
                        (N22)? mem[658] : 
                        (N24)? mem[759] : 1'b0;
  assign r_data_o[51] = (N17)? mem[51] : 
                        (N19)? mem[152] : 
                        (N21)? mem[253] : 
                        (N23)? mem[354] : 
                        (N18)? mem[455] : 
                        (N20)? mem[556] : 
                        (N22)? mem[657] : 
                        (N24)? mem[758] : 1'b0;
  assign r_data_o[50] = (N17)? mem[50] : 
                        (N19)? mem[151] : 
                        (N21)? mem[252] : 
                        (N23)? mem[353] : 
                        (N18)? mem[454] : 
                        (N20)? mem[555] : 
                        (N22)? mem[656] : 
                        (N24)? mem[757] : 1'b0;
  assign r_data_o[49] = (N17)? mem[49] : 
                        (N19)? mem[150] : 
                        (N21)? mem[251] : 
                        (N23)? mem[352] : 
                        (N18)? mem[453] : 
                        (N20)? mem[554] : 
                        (N22)? mem[655] : 
                        (N24)? mem[756] : 1'b0;
  assign r_data_o[48] = (N17)? mem[48] : 
                        (N19)? mem[149] : 
                        (N21)? mem[250] : 
                        (N23)? mem[351] : 
                        (N18)? mem[452] : 
                        (N20)? mem[553] : 
                        (N22)? mem[654] : 
                        (N24)? mem[755] : 1'b0;
  assign r_data_o[47] = (N17)? mem[47] : 
                        (N19)? mem[148] : 
                        (N21)? mem[249] : 
                        (N23)? mem[350] : 
                        (N18)? mem[451] : 
                        (N20)? mem[552] : 
                        (N22)? mem[653] : 
                        (N24)? mem[754] : 1'b0;
  assign r_data_o[46] = (N17)? mem[46] : 
                        (N19)? mem[147] : 
                        (N21)? mem[248] : 
                        (N23)? mem[349] : 
                        (N18)? mem[450] : 
                        (N20)? mem[551] : 
                        (N22)? mem[652] : 
                        (N24)? mem[753] : 1'b0;
  assign r_data_o[45] = (N17)? mem[45] : 
                        (N19)? mem[146] : 
                        (N21)? mem[247] : 
                        (N23)? mem[348] : 
                        (N18)? mem[449] : 
                        (N20)? mem[550] : 
                        (N22)? mem[651] : 
                        (N24)? mem[752] : 1'b0;
  assign r_data_o[44] = (N17)? mem[44] : 
                        (N19)? mem[145] : 
                        (N21)? mem[246] : 
                        (N23)? mem[347] : 
                        (N18)? mem[448] : 
                        (N20)? mem[549] : 
                        (N22)? mem[650] : 
                        (N24)? mem[751] : 1'b0;
  assign r_data_o[43] = (N17)? mem[43] : 
                        (N19)? mem[144] : 
                        (N21)? mem[245] : 
                        (N23)? mem[346] : 
                        (N18)? mem[447] : 
                        (N20)? mem[548] : 
                        (N22)? mem[649] : 
                        (N24)? mem[750] : 1'b0;
  assign r_data_o[42] = (N17)? mem[42] : 
                        (N19)? mem[143] : 
                        (N21)? mem[244] : 
                        (N23)? mem[345] : 
                        (N18)? mem[446] : 
                        (N20)? mem[547] : 
                        (N22)? mem[648] : 
                        (N24)? mem[749] : 1'b0;
  assign r_data_o[41] = (N17)? mem[41] : 
                        (N19)? mem[142] : 
                        (N21)? mem[243] : 
                        (N23)? mem[344] : 
                        (N18)? mem[445] : 
                        (N20)? mem[546] : 
                        (N22)? mem[647] : 
                        (N24)? mem[748] : 1'b0;
  assign r_data_o[40] = (N17)? mem[40] : 
                        (N19)? mem[141] : 
                        (N21)? mem[242] : 
                        (N23)? mem[343] : 
                        (N18)? mem[444] : 
                        (N20)? mem[545] : 
                        (N22)? mem[646] : 
                        (N24)? mem[747] : 1'b0;
  assign r_data_o[39] = (N17)? mem[39] : 
                        (N19)? mem[140] : 
                        (N21)? mem[241] : 
                        (N23)? mem[342] : 
                        (N18)? mem[443] : 
                        (N20)? mem[544] : 
                        (N22)? mem[645] : 
                        (N24)? mem[746] : 1'b0;
  assign r_data_o[38] = (N17)? mem[38] : 
                        (N19)? mem[139] : 
                        (N21)? mem[240] : 
                        (N23)? mem[341] : 
                        (N18)? mem[442] : 
                        (N20)? mem[543] : 
                        (N22)? mem[644] : 
                        (N24)? mem[745] : 1'b0;
  assign r_data_o[37] = (N17)? mem[37] : 
                        (N19)? mem[138] : 
                        (N21)? mem[239] : 
                        (N23)? mem[340] : 
                        (N18)? mem[441] : 
                        (N20)? mem[542] : 
                        (N22)? mem[643] : 
                        (N24)? mem[744] : 1'b0;
  assign r_data_o[36] = (N17)? mem[36] : 
                        (N19)? mem[137] : 
                        (N21)? mem[238] : 
                        (N23)? mem[339] : 
                        (N18)? mem[440] : 
                        (N20)? mem[541] : 
                        (N22)? mem[642] : 
                        (N24)? mem[743] : 1'b0;
  assign r_data_o[35] = (N17)? mem[35] : 
                        (N19)? mem[136] : 
                        (N21)? mem[237] : 
                        (N23)? mem[338] : 
                        (N18)? mem[439] : 
                        (N20)? mem[540] : 
                        (N22)? mem[641] : 
                        (N24)? mem[742] : 1'b0;
  assign r_data_o[34] = (N17)? mem[34] : 
                        (N19)? mem[135] : 
                        (N21)? mem[236] : 
                        (N23)? mem[337] : 
                        (N18)? mem[438] : 
                        (N20)? mem[539] : 
                        (N22)? mem[640] : 
                        (N24)? mem[741] : 1'b0;
  assign r_data_o[33] = (N17)? mem[33] : 
                        (N19)? mem[134] : 
                        (N21)? mem[235] : 
                        (N23)? mem[336] : 
                        (N18)? mem[437] : 
                        (N20)? mem[538] : 
                        (N22)? mem[639] : 
                        (N24)? mem[740] : 1'b0;
  assign r_data_o[32] = (N17)? mem[32] : 
                        (N19)? mem[133] : 
                        (N21)? mem[234] : 
                        (N23)? mem[335] : 
                        (N18)? mem[436] : 
                        (N20)? mem[537] : 
                        (N22)? mem[638] : 
                        (N24)? mem[739] : 1'b0;
  assign r_data_o[31] = (N17)? mem[31] : 
                        (N19)? mem[132] : 
                        (N21)? mem[233] : 
                        (N23)? mem[334] : 
                        (N18)? mem[435] : 
                        (N20)? mem[536] : 
                        (N22)? mem[637] : 
                        (N24)? mem[738] : 1'b0;
  assign r_data_o[30] = (N17)? mem[30] : 
                        (N19)? mem[131] : 
                        (N21)? mem[232] : 
                        (N23)? mem[333] : 
                        (N18)? mem[434] : 
                        (N20)? mem[535] : 
                        (N22)? mem[636] : 
                        (N24)? mem[737] : 1'b0;
  assign r_data_o[29] = (N17)? mem[29] : 
                        (N19)? mem[130] : 
                        (N21)? mem[231] : 
                        (N23)? mem[332] : 
                        (N18)? mem[433] : 
                        (N20)? mem[534] : 
                        (N22)? mem[635] : 
                        (N24)? mem[736] : 1'b0;
  assign r_data_o[28] = (N17)? mem[28] : 
                        (N19)? mem[129] : 
                        (N21)? mem[230] : 
                        (N23)? mem[331] : 
                        (N18)? mem[432] : 
                        (N20)? mem[533] : 
                        (N22)? mem[634] : 
                        (N24)? mem[735] : 1'b0;
  assign r_data_o[27] = (N17)? mem[27] : 
                        (N19)? mem[128] : 
                        (N21)? mem[229] : 
                        (N23)? mem[330] : 
                        (N18)? mem[431] : 
                        (N20)? mem[532] : 
                        (N22)? mem[633] : 
                        (N24)? mem[734] : 1'b0;
  assign r_data_o[26] = (N17)? mem[26] : 
                        (N19)? mem[127] : 
                        (N21)? mem[228] : 
                        (N23)? mem[329] : 
                        (N18)? mem[430] : 
                        (N20)? mem[531] : 
                        (N22)? mem[632] : 
                        (N24)? mem[733] : 1'b0;
  assign r_data_o[25] = (N17)? mem[25] : 
                        (N19)? mem[126] : 
                        (N21)? mem[227] : 
                        (N23)? mem[328] : 
                        (N18)? mem[429] : 
                        (N20)? mem[530] : 
                        (N22)? mem[631] : 
                        (N24)? mem[732] : 1'b0;
  assign r_data_o[24] = (N17)? mem[24] : 
                        (N19)? mem[125] : 
                        (N21)? mem[226] : 
                        (N23)? mem[327] : 
                        (N18)? mem[428] : 
                        (N20)? mem[529] : 
                        (N22)? mem[630] : 
                        (N24)? mem[731] : 1'b0;
  assign r_data_o[23] = (N17)? mem[23] : 
                        (N19)? mem[124] : 
                        (N21)? mem[225] : 
                        (N23)? mem[326] : 
                        (N18)? mem[427] : 
                        (N20)? mem[528] : 
                        (N22)? mem[629] : 
                        (N24)? mem[730] : 1'b0;
  assign r_data_o[22] = (N17)? mem[22] : 
                        (N19)? mem[123] : 
                        (N21)? mem[224] : 
                        (N23)? mem[325] : 
                        (N18)? mem[426] : 
                        (N20)? mem[527] : 
                        (N22)? mem[628] : 
                        (N24)? mem[729] : 1'b0;
  assign r_data_o[21] = (N17)? mem[21] : 
                        (N19)? mem[122] : 
                        (N21)? mem[223] : 
                        (N23)? mem[324] : 
                        (N18)? mem[425] : 
                        (N20)? mem[526] : 
                        (N22)? mem[627] : 
                        (N24)? mem[728] : 1'b0;
  assign r_data_o[20] = (N17)? mem[20] : 
                        (N19)? mem[121] : 
                        (N21)? mem[222] : 
                        (N23)? mem[323] : 
                        (N18)? mem[424] : 
                        (N20)? mem[525] : 
                        (N22)? mem[626] : 
                        (N24)? mem[727] : 1'b0;
  assign r_data_o[19] = (N17)? mem[19] : 
                        (N19)? mem[120] : 
                        (N21)? mem[221] : 
                        (N23)? mem[322] : 
                        (N18)? mem[423] : 
                        (N20)? mem[524] : 
                        (N22)? mem[625] : 
                        (N24)? mem[726] : 1'b0;
  assign r_data_o[18] = (N17)? mem[18] : 
                        (N19)? mem[119] : 
                        (N21)? mem[220] : 
                        (N23)? mem[321] : 
                        (N18)? mem[422] : 
                        (N20)? mem[523] : 
                        (N22)? mem[624] : 
                        (N24)? mem[725] : 1'b0;
  assign r_data_o[17] = (N17)? mem[17] : 
                        (N19)? mem[118] : 
                        (N21)? mem[219] : 
                        (N23)? mem[320] : 
                        (N18)? mem[421] : 
                        (N20)? mem[522] : 
                        (N22)? mem[623] : 
                        (N24)? mem[724] : 1'b0;
  assign r_data_o[16] = (N17)? mem[16] : 
                        (N19)? mem[117] : 
                        (N21)? mem[218] : 
                        (N23)? mem[319] : 
                        (N18)? mem[420] : 
                        (N20)? mem[521] : 
                        (N22)? mem[622] : 
                        (N24)? mem[723] : 1'b0;
  assign r_data_o[15] = (N17)? mem[15] : 
                        (N19)? mem[116] : 
                        (N21)? mem[217] : 
                        (N23)? mem[318] : 
                        (N18)? mem[419] : 
                        (N20)? mem[520] : 
                        (N22)? mem[621] : 
                        (N24)? mem[722] : 1'b0;
  assign r_data_o[14] = (N17)? mem[14] : 
                        (N19)? mem[115] : 
                        (N21)? mem[216] : 
                        (N23)? mem[317] : 
                        (N18)? mem[418] : 
                        (N20)? mem[519] : 
                        (N22)? mem[620] : 
                        (N24)? mem[721] : 1'b0;
  assign r_data_o[13] = (N17)? mem[13] : 
                        (N19)? mem[114] : 
                        (N21)? mem[215] : 
                        (N23)? mem[316] : 
                        (N18)? mem[417] : 
                        (N20)? mem[518] : 
                        (N22)? mem[619] : 
                        (N24)? mem[720] : 1'b0;
  assign r_data_o[12] = (N17)? mem[12] : 
                        (N19)? mem[113] : 
                        (N21)? mem[214] : 
                        (N23)? mem[315] : 
                        (N18)? mem[416] : 
                        (N20)? mem[517] : 
                        (N22)? mem[618] : 
                        (N24)? mem[719] : 1'b0;
  assign r_data_o[11] = (N17)? mem[11] : 
                        (N19)? mem[112] : 
                        (N21)? mem[213] : 
                        (N23)? mem[314] : 
                        (N18)? mem[415] : 
                        (N20)? mem[516] : 
                        (N22)? mem[617] : 
                        (N24)? mem[718] : 1'b0;
  assign r_data_o[10] = (N17)? mem[10] : 
                        (N19)? mem[111] : 
                        (N21)? mem[212] : 
                        (N23)? mem[313] : 
                        (N18)? mem[414] : 
                        (N20)? mem[515] : 
                        (N22)? mem[616] : 
                        (N24)? mem[717] : 1'b0;
  assign r_data_o[9] = (N17)? mem[9] : 
                       (N19)? mem[110] : 
                       (N21)? mem[211] : 
                       (N23)? mem[312] : 
                       (N18)? mem[413] : 
                       (N20)? mem[514] : 
                       (N22)? mem[615] : 
                       (N24)? mem[716] : 1'b0;
  assign r_data_o[8] = (N17)? mem[8] : 
                       (N19)? mem[109] : 
                       (N21)? mem[210] : 
                       (N23)? mem[311] : 
                       (N18)? mem[412] : 
                       (N20)? mem[513] : 
                       (N22)? mem[614] : 
                       (N24)? mem[715] : 1'b0;
  assign r_data_o[7] = (N17)? mem[7] : 
                       (N19)? mem[108] : 
                       (N21)? mem[209] : 
                       (N23)? mem[310] : 
                       (N18)? mem[411] : 
                       (N20)? mem[512] : 
                       (N22)? mem[613] : 
                       (N24)? mem[714] : 1'b0;
  assign r_data_o[6] = (N17)? mem[6] : 
                       (N19)? mem[107] : 
                       (N21)? mem[208] : 
                       (N23)? mem[309] : 
                       (N18)? mem[410] : 
                       (N20)? mem[511] : 
                       (N22)? mem[612] : 
                       (N24)? mem[713] : 1'b0;
  assign r_data_o[5] = (N17)? mem[5] : 
                       (N19)? mem[106] : 
                       (N21)? mem[207] : 
                       (N23)? mem[308] : 
                       (N18)? mem[409] : 
                       (N20)? mem[510] : 
                       (N22)? mem[611] : 
                       (N24)? mem[712] : 1'b0;
  assign r_data_o[4] = (N17)? mem[4] : 
                       (N19)? mem[105] : 
                       (N21)? mem[206] : 
                       (N23)? mem[307] : 
                       (N18)? mem[408] : 
                       (N20)? mem[509] : 
                       (N22)? mem[610] : 
                       (N24)? mem[711] : 1'b0;
  assign r_data_o[3] = (N17)? mem[3] : 
                       (N19)? mem[104] : 
                       (N21)? mem[205] : 
                       (N23)? mem[306] : 
                       (N18)? mem[407] : 
                       (N20)? mem[508] : 
                       (N22)? mem[609] : 
                       (N24)? mem[710] : 1'b0;
  assign r_data_o[2] = (N17)? mem[2] : 
                       (N19)? mem[103] : 
                       (N21)? mem[204] : 
                       (N23)? mem[305] : 
                       (N18)? mem[406] : 
                       (N20)? mem[507] : 
                       (N22)? mem[608] : 
                       (N24)? mem[709] : 1'b0;
  assign r_data_o[1] = (N17)? mem[1] : 
                       (N19)? mem[102] : 
                       (N21)? mem[203] : 
                       (N23)? mem[304] : 
                       (N18)? mem[405] : 
                       (N20)? mem[506] : 
                       (N22)? mem[607] : 
                       (N24)? mem[708] : 1'b0;
  assign r_data_o[0] = (N17)? mem[0] : 
                       (N19)? mem[101] : 
                       (N21)? mem[202] : 
                       (N23)? mem[303] : 
                       (N18)? mem[404] : 
                       (N20)? mem[505] : 
                       (N22)? mem[606] : 
                       (N24)? mem[707] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_807_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_806_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_805_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_804_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_803_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_802_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_801_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_800_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_799_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_798_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_797_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_796_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_795_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_794_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_793_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_792_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_791_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_790_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_789_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_788_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_787_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_786_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_785_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_784_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_783_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_782_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_781_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_780_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_779_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_778_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_777_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_776_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_775_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_774_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_773_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_772_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_771_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_770_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_769_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_768_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_767_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_766_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_765_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_764_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_763_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_762_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_761_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_760_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_759_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_758_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_757_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_756_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_755_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_754_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_753_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_752_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_751_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_750_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_749_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_748_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_747_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_746_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_745_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_744_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_743_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_742_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_741_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_740_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_739_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_738_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_737_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_736_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_735_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_734_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_733_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_732_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_731_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_730_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_729_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_728_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_727_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_726_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_725_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_724_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_723_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_722_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_721_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_720_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_719_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_718_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_717_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_716_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_715_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_714_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_713_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_712_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_711_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_710_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_709_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N49) begin
      mem_708_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N48) begin
      mem_707_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_706_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_705_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_704_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_703_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_702_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_701_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_700_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_699_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_698_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_697_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_696_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_695_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_694_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_693_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_692_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_691_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_690_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_689_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_688_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_687_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_686_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_685_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_684_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_683_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_682_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_681_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_680_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_679_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_678_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_677_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_676_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_675_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_674_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_673_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_672_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_671_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_670_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_669_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_668_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_667_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_666_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_665_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_664_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_663_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_662_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_661_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_660_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_659_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_658_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_657_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_656_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_655_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_654_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_653_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_652_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_651_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_650_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_649_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_648_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_647_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_646_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_645_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_644_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_643_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_642_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_641_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_640_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_639_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_638_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_637_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_636_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_635_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_634_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_633_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_632_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_631_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_630_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_629_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_628_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_627_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_626_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_625_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_624_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_623_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_622_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_621_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_620_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_619_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_618_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_617_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_616_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_615_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_614_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_613_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_612_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_611_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_610_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_609_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_608_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N47) begin
      mem_607_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N46) begin
      mem_606_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_605_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_604_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_603_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_602_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_601_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_600_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_599_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_598_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_597_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_596_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_595_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_594_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_593_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_592_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_591_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_590_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_589_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_588_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_587_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_586_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_585_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_584_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_583_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_582_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_581_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_580_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_579_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_578_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_577_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_576_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_575_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_574_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_573_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_572_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_571_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_570_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_569_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_568_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_567_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_566_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_565_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_564_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_563_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_562_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_561_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_560_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_559_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_558_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_557_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_556_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_555_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_554_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_553_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_552_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_551_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_550_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_549_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_548_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_547_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_546_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_545_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_544_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_543_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_542_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_541_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_540_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_539_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_538_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_537_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_536_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_535_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_534_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_533_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_532_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_531_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_530_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_529_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_528_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_527_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_526_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_525_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_524_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_523_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_522_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_521_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_520_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_519_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_518_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_517_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_516_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_515_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_514_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_513_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_512_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_511_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_510_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_509_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_508_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_507_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N45) begin
      mem_506_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N44) begin
      mem_505_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_504_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_503_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_502_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_501_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_500_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_499_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_498_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_497_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_496_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_495_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_494_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_493_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_492_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_491_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_490_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_489_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_488_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_487_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_486_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_485_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_484_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_483_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_482_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_481_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_480_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_479_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_478_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_477_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_476_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_475_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_474_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_473_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_472_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_471_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_470_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_469_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_468_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_467_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_466_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_465_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_464_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_463_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_462_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_461_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_460_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_459_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_458_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_457_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_456_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_455_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_454_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_453_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_452_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_451_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_450_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_449_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_448_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_447_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_446_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_445_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_444_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_443_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_442_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_441_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_440_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_439_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_438_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_437_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_436_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_435_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_434_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_433_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_432_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_431_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_430_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_429_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_428_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_427_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_426_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_425_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_424_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_423_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_422_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_421_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_420_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_419_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_418_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_417_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_416_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_415_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_414_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_413_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_412_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_411_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_410_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_409_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_408_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_407_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_406_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N43) begin
      mem_405_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N42) begin
      mem_404_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_403_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_402_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_401_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_400_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_399_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_398_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_397_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_396_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_395_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_394_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_393_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_392_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_391_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_390_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_389_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_388_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_387_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_386_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_385_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_384_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_383_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_382_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_381_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_380_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_379_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_378_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_377_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_376_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_375_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_374_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_373_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_372_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_371_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_370_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_369_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_368_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_367_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_366_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_365_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_364_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_363_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_362_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_361_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_360_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_359_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_358_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_357_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_356_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_355_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_354_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_353_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_352_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_351_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_350_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_349_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_348_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_347_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_346_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_345_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_344_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_343_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_342_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_341_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_340_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_339_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_338_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_337_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_336_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_335_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_334_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_333_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_332_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_331_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_330_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_329_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_328_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_327_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_326_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_325_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_324_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_323_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_322_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_321_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_320_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_319_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_318_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_317_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_316_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_315_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_314_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_313_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_312_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_311_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_310_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_309_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_308_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_307_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_306_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_305_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_304_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_303_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_302_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_301_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_300_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_299_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_298_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_297_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_296_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_295_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_294_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_293_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_292_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_291_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_290_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_289_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_288_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_287_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_286_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_285_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_284_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_283_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_282_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_281_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_280_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_279_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_278_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_277_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_276_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_275_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_274_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_273_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_272_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_271_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_270_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_269_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_268_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_267_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_266_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_265_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_264_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_263_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_262_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_261_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_260_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_259_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_258_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_257_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_256_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_255_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_254_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_253_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_252_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_251_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_250_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_249_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_248_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_247_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_246_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_245_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_244_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_243_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_242_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_241_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_240_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_239_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_238_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_237_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_236_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_235_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_234_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_233_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_232_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_231_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_230_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_229_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_228_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_227_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_226_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_225_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_224_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_223_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_222_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_221_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_220_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_219_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_218_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_217_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_216_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_215_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_214_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_213_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_212_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_211_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_210_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_209_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_208_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_207_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_206_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_205_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_204_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_203_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_202_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_201_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_200_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_199_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_198_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_197_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_196_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_195_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_194_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_193_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_192_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_191_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_190_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_189_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_188_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_187_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_186_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_185_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_184_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_183_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_182_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_181_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_180_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_179_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_178_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_177_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_176_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_175_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_174_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_173_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_172_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_171_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_170_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_169_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_168_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_167_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_166_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_165_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_164_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_163_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_162_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_161_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_160_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_159_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_158_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_157_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_156_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_155_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_154_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_153_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_152_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_151_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_150_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_149_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_148_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_147_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_146_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_145_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_144_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_143_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_142_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_141_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_140_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_139_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_138_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_137_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_136_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_135_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_134_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_133_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_132_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_131_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_130_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_129_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_128_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_127_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_126_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_125_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_124_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_123_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_122_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_121_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_120_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_119_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_118_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_117_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_116_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_115_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_114_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_113_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_112_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_111_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_110_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_109_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_108_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_107_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_106_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_105_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_104_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_103_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_102_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_101_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_100_sv2v_reg <= w_data_i[100];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_99_sv2v_reg <= w_data_i[99];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_98_sv2v_reg <= w_data_i[98];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_97_sv2v_reg <= w_data_i[97];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_96_sv2v_reg <= w_data_i[96];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_95_sv2v_reg <= w_data_i[95];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_94_sv2v_reg <= w_data_i[94];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_93_sv2v_reg <= w_data_i[93];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_92_sv2v_reg <= w_data_i[92];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_91_sv2v_reg <= w_data_i[91];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_90_sv2v_reg <= w_data_i[90];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_89_sv2v_reg <= w_data_i[89];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_88_sv2v_reg <= w_data_i[88];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_87_sv2v_reg <= w_data_i[87];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_86_sv2v_reg <= w_data_i[86];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_85_sv2v_reg <= w_data_i[85];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_84_sv2v_reg <= w_data_i[84];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_83_sv2v_reg <= w_data_i[83];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_82_sv2v_reg <= w_data_i[82];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_81_sv2v_reg <= w_data_i[81];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_80_sv2v_reg <= w_data_i[80];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_79_sv2v_reg <= w_data_i[79];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_78_sv2v_reg <= w_data_i[78];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_77_sv2v_reg <= w_data_i[77];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_76_sv2v_reg <= w_data_i[76];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_75_sv2v_reg <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_74_sv2v_reg <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_73_sv2v_reg <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_72_sv2v_reg <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_71_sv2v_reg <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_70_sv2v_reg <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_69_sv2v_reg <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_68_sv2v_reg <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_67_sv2v_reg <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_66_sv2v_reg <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_65_sv2v_reg <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_64_sv2v_reg <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_63_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_62_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_61_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_60_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_59_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_58_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_57_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_56_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_55_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_54_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_53_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_52_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_51_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_50_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_49_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_48_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_47_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_46_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_45_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_44_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_43_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_42_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_41_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_40_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_39_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_38_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_37_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_36_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_35_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_34_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_33_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_32_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_31_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_30_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_29_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_28_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_27_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_26_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_25_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_24_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_23_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_22_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_21_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_20_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_19_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_18_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_17_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_16_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_15_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_14_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_13_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_12_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_11_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_10_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_9_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_8_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_7_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_6_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_5_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_4_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_3_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_2_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_1_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end

  assign N50 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N50 & w_addr_i[2];
  assign N51 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N51 & w_addr_i[2];
  assign N52 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N52 & w_addr_i[2];
  assign N53 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N53 & w_addr_i[2];
  assign N29 = N50 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N51 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N52 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N53 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N33, N32, N32, N31, N31, N30, N30, N29, N29, N28, N28, N27, N27, N26, N26 } : 
                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

endmodule